
module b20 ( si_31_, si_30_, si_29_, si_28_, si_27_, si_26_, si_25_, si_24_, 
        si_23_, si_22_, si_21_, si_20_, si_19_, si_18_, si_17_, si_16_, si_15_, 
        si_14_, si_13_, si_12_, si_11_, si_10_, si_9_, si_8_, si_7_, si_6_, 
        si_5_, si_4_, si_3_, si_2_, si_1_, si_0_, so_19_, so_18_, so_17_, 
        so_16_, so_15_, so_14_, so_13_, so_12_, so_11_, so_10_, so_9_, so_8_, 
        so_7_, so_6_, so_5_, so_4_, so_3_, so_2_, so_1_, so_0_, clock, 
        test_si6, test_si5, test_si4, test_si3, test_si2, Scan_In, Scan_Enable, 
        reset, test_so2, Scan_Out, wr, rd, test_si10, test_si9, test_si8, 
        test_si7, test_so10, test_so9, test_so8, test_so7, test_so6, test_so5, 
        test_so4, test_so3 );
  input si_31_, si_30_, si_29_, si_28_, si_27_, si_26_, si_25_, si_24_, si_23_,
         si_22_, si_21_, si_20_, si_19_, si_18_, si_17_, si_16_, si_15_,
         si_14_, si_13_, si_12_, si_11_, si_10_, si_9_, si_8_, si_7_, si_6_,
         si_5_, si_4_, si_3_, si_2_, si_1_, si_0_, clock, test_si6, test_si5,
         test_si4, test_si3, test_si2, Scan_In, Scan_Enable, reset, test_si10,
         test_si9, test_si8, test_si7;
  output so_19_, so_18_, so_17_, so_16_, so_15_, so_14_, so_13_, so_12_,
         so_11_, so_10_, so_9_, so_8_, so_7_, so_6_, so_5_, so_4_, so_3_,
         so_2_, so_1_, so_0_, test_so2, Scan_Out, wr, rd, test_so10, test_so9,
         test_so8, test_so7, test_so6, test_so5, test_so4, test_so3;
  wire   SYNOPSYS_UNCONNECTED_0, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12;
  tri   si_31_;
  tri   si_30_;
  tri   si_29_;
  tri   si_28_;
  tri   si_27_;
  tri   si_26_;
  tri   si_25_;
  tri   si_24_;
  tri   si_23_;
  tri   si_22_;
  tri   si_21_;
  tri   si_20_;
  tri   si_19_;
  tri   si_18_;
  tri   si_17_;
  tri   si_16_;
  tri   si_15_;
  tri   si_14_;
  tri   si_13_;
  tri   si_12_;
  tri   si_11_;
  tri   si_10_;
  tri   si_9_;
  tri   si_8_;
  tri   si_7_;
  tri   si_6_;
  tri   si_5_;
  tri   si_4_;
  tri   si_3_;
  tri   si_2_;
  tri   si_1_;
  tri   si_0_;
  tri   so_19_;
  tri   so_18_;
  tri   so_17_;
  tri   so_16_;
  tri   so_15_;
  tri   so_14_;
  tri   so_13_;
  tri   so_12_;
  tri   so_11_;
  tri   so_10_;
  tri   so_9_;
  tri   so_8_;
  tri   so_7_;
  tri   so_6_;
  tri   so_5_;
  tri   so_4_;
  tri   so_3_;
  tri   so_2_;
  tri   so_1_;
  tri   so_0_;
  tri   clock;
  tri   test_si6;
  tri   test_si5;
  tri   test_si4;
  tri   test_si3;
  tri   test_si2;
  tri   Scan_In;
  tri   Scan_Enable;
  tri   reset;
  tri   test_so2;
  tri   Scan_Out;
  tri   wr;
  tri   rd;
  tri   test_si10;
  tri   test_si9;
  tri   test_si8;
  tri   test_si7;
  tri   test_so10;
  tri   test_so9;
  tri   test_so8;
  tri   test_so7;
  tri   test_so6;
  tri   test_so5;
  tri   test_so4;
  tri   test_so3;
  tri   P2_N5203;
  tri   P2_N5352;
  tri   P2_N5351;
  tri   P2_N5350;
  tri   P2_N5349;
  tri   P2_N5348;
  tri   P2_N5347;
  tri   P2_N5346;
  tri   P2_N5345;
  tri   P2_N5344;
  tri   P2_N5343;
  tri   P2_N5342;
  tri   P2_N5341;
  tri   P2_N5340;
  tri   P2_N5339;
  tri   P2_N5338;
  tri   P2_N5337;
  tri   P2_N5336;
  tri   P2_N5335;
  tri   P2_N5334;
  tri   P2_N5333;
  tri   P2_N5332;
  tri   P2_N5331;
  tri   P2_N5330;
  tri   P2_N5329;
  tri   P2_N5328;
  tri   P2_N5327;
  tri   P2_N5326;
  tri   P2_N5325;
  tri   P2_N5324;
  tri   P2_N5323;
  tri   P2_N5322;
  tri   P2_N5321;
  tri   P2_N5037;
  tri   P2_N5036;
  tri   P2_N5035;
  tri   P2_N5034;
  tri   P2_N5033;
  tri   P2_N5032;
  tri   P2_N5031;
  tri   P2_N5030;
  tri   P2_N5029;
  tri   P2_N5028;
  tri   P2_N5027;
  tri   P2_N5026;
  tri   P2_N5025;
  tri   P2_N5024;
  tri   P2_N5023;
  tri   P2_N5022;
  tri   P2_N5021;
  tri   P2_N5020;
  tri   P2_N5019;
  tri   P2_N5018;
  tri   P2_N5017;
  tri   P2_N5016;
  tri   n7275;
  tri   P2_N5014;
  tri   P2_N5013;
  tri   P2_N5012;
  tri   P2_N5011;
  tri   P2_N5010;
  tri   P2_N5009;
  tri   P2_N5008;
  tri   P2_N5007;
  tri   P2_N5006;
  tri   P2_N5284;
  tri   P2_N5353;
  tri   n7263;
  tri   n7259;
  tri   n7252;
  tri   n7248;
  tri   n7247;
  tri   n7243;
  tri   n7239;
  tri   n7234;
  tri   P2_N5097;
  tri   P2_N5098;
  tri   P2_N5081;
  tri   n7216;
  tri   n7210;
  tri   P2_N5084;
  tri   P2_N5085;
  tri   n7202;
  tri   P2_N5087;
  tri   P2_N5088;
  tri   n7187;
  tri   n7181;
  tri   n7177;
  tri   n7173;
  tri   n7165;
  tri   P2_N5077;
  tri   n7157;
  tri   n7153;
  tri   P2_N5080;
  tri   n2919;
  tri   n7242;
  tri   P2_N5079;
  tri   n7222;
  tri   n7224;
  tri   n7229;
  tri   n7237;
  tri   n7238;
  tri   P2_N5094;
  tri   n7253;
  tri   n7260;
  tri   n7264;
  tri   n7188;
  tri   n7195;
  tri   n7197;
  tri   n7201;
  tri   n7205;
  tri   n7208;
  tri   n7211;
  tri   n7214;
  tri   n7219;
  tri   n7149;
  tri   n7158;
  tri   n7164;
  tri   n7166;
  tri   n7174;
  tri   n7178;
  tri   n7182;
  tri   n7186;
  tri   n7035;
  tri   P2_N2633;
  tri   P2_N2632;
  tri   P2_N2631;
  tri   P2_N2630;
  tri   P2_N2629;
  tri   P2_N2628;
  tri   P2_N2627;
  tri   P2_N2626;
  tri   P2_N2625;
  tri   P2_N2624;
  tri   P2_N2623;
  tri   P2_N2622;
  tri   P2_N2621;
  tri   P2_N2620;
  tri   P2_N2619;
  tri   P2_N2618;
  tri   P2_N2617;
  tri   P2_N2616;
  tri   P2_N2615;
  tri   P2_N2614;
  tri   P2_N2613;
  tri   P2_N2612;
  tri   P2_N2611;
  tri   P2_N2610;
  tri   P2_N2609;
  tri   P2_N2608;
  tri   P2_N2607;
  tri   P2_N2606;
  tri   P2_N2605;
  tri   P2_N2875;
  tri   P2_N2874;
  tri   P2_N2873;
  tri   P2_N2872;
  tri   P2_N2871;
  tri   P2_N2870;
  tri   P2_N2869;
  tri   P2_N2868;
  tri   P2_N2867;
  tri   P2_N2866;
  tri   P2_N2865;
  tri   P2_N2864;
  tri   P2_N2863;
  tri   P2_N2862;
  tri   P2_N2861;
  tri   P2_N2860;
  tri   P2_N2859;
  tri   P2_N2858;
  tri   P2_N2857;
  tri   P2_N2856;
  tri   P2_N2855;
  tri   P2_N2854;
  tri   P2_N2853;
  tri   P2_N2852;
  tri   P2_N2851;
  tri   P2_N2850;
  tri   P2_N2849;
  tri   P2_N2848;
  tri   P2_N2847;
  tri   P2_N5072;
  tri   n7231;
  tri   P2_N5095;
  tri   P2_N5092;
  tri   P2_N5091;
  tri   P2_N5090;
  tri   n7194;
  tri   n7198;
  tri   P2_N5086;
  tri   P2_N5083;
  tri   P2_N5082;
  tri   n7151;
  tri   P2_N5078;
  tri   P2_N5075;
  tri   P2_N5074;
  tri   P2_N5073;
  tri   n7184;
  tri   P2_N3006;
  tri   P2_N3005;
  tri   P2_N3004;
  tri   P2_N3003;
  tri   P2_N3002;
  tri   P2_N3001;
  tri   P2_N3000;
  tri   P2_N2999;
  tri   P2_N2998;
  tri   P2_N2997;
  tri   P2_N2996;
  tri   P2_N2995;
  tri   P2_N2994;
  tri   P2_N2993;
  tri   P2_N2992;
  tri   P2_N2991;
  tri   P2_N2990;
  tri   P2_N2989;
  tri   P2_N2988;
  tri   P2_N2987;
  tri   P2_N2986;
  tri   P2_N2985;
  tri   P2_N2984;
  tri   P2_N2983;
  tri   P2_N2982;
  tri   P2_N2981;
  tri   P2_N2980;
  tri   P2_N2979;
  tri   P2_N2978;
  tri   P2_N3248;
  tri   P2_N3247;
  tri   P2_N3246;
  tri   P2_N3245;
  tri   P2_N3244;
  tri   P2_N3243;
  tri   P2_N3242;
  tri   P2_N3241;
  tri   P2_N3240;
  tri   P2_N3239;
  tri   P2_N3238;
  tri   P2_N3237;
  tri   P2_N3236;
  tri   P2_N3235;
  tri   P2_N3234;
  tri   P2_N3233;
  tri   P2_N3232;
  tri   P2_N3231;
  tri   P2_N3230;
  tri   P2_N3229;
  tri   P2_N3228;
  tri   P2_N3227;
  tri   P2_N3226;
  tri   P2_N3225;
  tri   P2_N3224;
  tri   P2_N3223;
  tri   P2_N3222;
  tri   P2_N3221;
  tri   P2_N3220;
  tri   P2_N5093;
  tri   P2_N5089;
  tri   P2_N3379;
  tri   P2_N3378;
  tri   P2_N3377;
  tri   P2_N3376;
  tri   P2_N3375;
  tri   P2_N3374;
  tri   P2_N3373;
  tri   P2_N3372;
  tri   P2_N3371;
  tri   P2_N3370;
  tri   P2_N3369;
  tri   P2_N3368;
  tri   P2_N3367;
  tri   P2_N3366;
  tri   P2_N3365;
  tri   P2_N3364;
  tri   P2_N3363;
  tri   P2_N3362;
  tri   P2_N3361;
  tri   P2_N3360;
  tri   P2_N3359;
  tri   P2_N3358;
  tri   P2_N3357;
  tri   P2_N3356;
  tri   P2_N3355;
  tri   P2_N3354;
  tri   P2_N3353;
  tri   P2_N3352;
  tri   P2_N3351;
  tri   P2_N3621;
  tri   P2_N3620;
  tri   P2_N3619;
  tri   P2_N3618;
  tri   P2_N3617;
  tri   P2_N3616;
  tri   P2_N3615;
  tri   P2_N3614;
  tri   P2_N3613;
  tri   P2_N3612;
  tri   P2_N3611;
  tri   P2_N3610;
  tri   P2_N3609;
  tri   P2_N3608;
  tri   P2_N3607;
  tri   P2_N3606;
  tri   P2_N3605;
  tri   P2_N3604;
  tri   P2_N3603;
  tri   P2_N3602;
  tri   P2_N3601;
  tri   P2_N3600;
  tri   P2_N3599;
  tri   P2_N3598;
  tri   P2_N3597;
  tri   P2_N3596;
  tri   P2_N3595;
  tri   P2_N3594;
  tri   P2_N3593;
  tri   n7206;
  tri   n7209;
  tri   n7154;
  tri   P2_N5076;
  tri   P2_N3752;
  tri   P2_N3751;
  tri   P2_N3750;
  tri   P2_N3749;
  tri   P2_N3748;
  tri   P2_N3747;
  tri   P2_N3746;
  tri   P2_N3745;
  tri   P2_N3744;
  tri   P2_N3743;
  tri   P2_N3742;
  tri   P2_N3741;
  tri   P2_N3740;
  tri   P2_N3739;
  tri   P2_N3738;
  tri   P2_N3737;
  tri   P2_N3736;
  tri   P2_N3735;
  tri   P2_N3734;
  tri   P2_N3733;
  tri   P2_N3732;
  tri   P2_N3731;
  tri   P2_N3730;
  tri   P2_N3729;
  tri   P2_N3728;
  tri   P2_N3727;
  tri   P2_N3726;
  tri   P2_N3725;
  tri   P2_N3724;
  tri   P2_N3994;
  tri   P2_N3993;
  tri   P2_N3992;
  tri   P2_N3991;
  tri   P2_N3990;
  tri   P2_N3989;
  tri   P2_N3988;
  tri   P2_N3987;
  tri   P2_N3986;
  tri   P2_N3985;
  tri   P2_N3984;
  tri   P2_N3983;
  tri   P2_N3982;
  tri   P2_N3981;
  tri   P2_N3980;
  tri   P2_N3979;
  tri   P2_N3978;
  tri   P2_N3977;
  tri   P2_N3976;
  tri   P2_N3975;
  tri   P2_N3974;
  tri   P2_N3973;
  tri   P2_N3972;
  tri   P2_N3971;
  tri   P2_N3970;
  tri   P2_N3969;
  tri   P2_N3968;
  tri   P2_N3967;
  tri   P2_N3966;
  tri   n7220;
  tri   P2_N4125;
  tri   P2_N4124;
  tri   P2_N4123;
  tri   P2_N4122;
  tri   P2_N4121;
  tri   P2_N4120;
  tri   P2_N4119;
  tri   P2_N4118;
  tri   P2_N4117;
  tri   P2_N4116;
  tri   P2_N4115;
  tri   P2_N4114;
  tri   P2_N4113;
  tri   P2_N4112;
  tri   P2_N4111;
  tri   P2_N4110;
  tri   P2_N4109;
  tri   P2_N4108;
  tri   P2_N4107;
  tri   P2_N4106;
  tri   P2_N4105;
  tri   P2_N4104;
  tri   P2_N4103;
  tri   P2_N4102;
  tri   P2_N4101;
  tri   P2_N4100;
  tri   P2_N4099;
  tri   P2_N4098;
  tri   P2_N4097;
  tri   P2_N4277;
  tri   P2_N4276;
  tri   P2_N4275;
  tri   P2_N4274;
  tri   P2_N4273;
  tri   P2_N4272;
  tri   P2_N4271;
  tri   P2_N4270;
  tri   P2_N4269;
  tri   P2_N4268;
  tri   P2_N4267;
  tri   P2_N4266;
  tri   P2_N4265;
  tri   P2_N4264;
  tri   P2_N4263;
  tri   P2_N4262;
  tri   P2_N4261;
  tri   P2_N4260;
  tri   P2_N4259;
  tri   P2_N4258;
  tri   P2_N4257;
  tri   P2_N4256;
  tri   P2_N4255;
  tri   P2_N4254;
  tri   P2_N4253;
  tri   P2_N4252;
  tri   P2_N4251;
  tri   P2_N4250;
  tri   P2_N4249;
  tri   P2_N362;
  tri   n18939;
  tri   n10111;
  tri   n6680;
  tri   n6679;
  tri   n6678;
  tri   n6677;
  tri   n6676;
  tri   n6675;
  tri   n6674;
  tri   n6673;
  tri   n6672;
  tri   n6671;
  tri   n10249;
  tri   n6670;
  tri   n6669;
  tri   n6668;
  tri   n6667;
  tri   n6666;
  tri   n6665;
  tri   n6664;
  tri   n9837;
  tri   P2_N344;
  tri   n6774;
  tri   n6772;
  tri   n6768;
  tri   n6764;
  tri   n6769;
  tri   n6765;
  tri   n6761;
  tri   n6756;
  tri   n6760;
  tri   n6757;
  tri   n6752;
  tri   n6748;
  tri   n6753;
  tri   n6749;
  tri   n6745;
  tri   n6743;
  tri   n6735;
  tri   n6733;
  tri   n6731;
  tri   P2_N4862;
  tri   P2_N4861;
  tri   P2_N4860;
  tri   P2_N4859;
  tri   P2_N4858;
  tri   P2_N4857;
  tri   P2_N4856;
  tri   P2_N4855;
  tri   P2_N4854;
  tri   P2_N4853;
  tri   P2_N4852;
  tri   P2_N4851;
  tri   P2_N4850;
  tri   P2_N4849;
  tri   P2_N4848;
  tri   P2_N4847;
  tri   P2_N4846;
  tri   P2_N4845;
  tri   P2_N4844;
  tri   P2_N4843;
  tri   n18997;
  tri   n10116;
  tri   n6663;
  tri   n6662;
  tri   n6661;
  tri   n6660;
  tri   n6659;
  tri   n6658;
  tri   n6657;
  tri   n6656;
  tri   n6655;
  tri   n6654;
  tri   n6653;
  tri   n6652;
  tri   n6651;
  tri   n6650;
  tri   n6649;
  tri   n6648;
  tri   n6721;
  tri   n6720;
  tri   n9842;
  tri   P2_N4882;
  tri   P2_N4881;
  tri   P2_N4880;
  tri   P2_N4879;
  tri   P2_N4878;
  tri   P2_N4877;
  tri   P2_N4876;
  tri   P2_N4875;
  tri   P2_N4874;
  tri   P2_N4873;
  tri   P2_N4872;
  tri   P2_N4871;
  tri   P2_N4870;
  tri   P2_N4869;
  tri   P2_N4868;
  tri   P2_N4867;
  tri   P2_N4866;
  tri   P2_N4865;
  tri   P2_N4864;
  tri   P2_N4863;
  tri   P2_N5135;
  tri   P1_N5150;
  tri   P1_N5164;
  tri   P1_N5165;
  tri   n7117;
  tri   P1_N5176;
  tri   P1_N5175;
  tri   n7129;
  tri   P1_N5173;
  tri   P1_N5172;
  tri   n7089;
  tri   n7093;
  tri   n7096;
  tri   P1_N5168;
  tri   n7103;
  tri   P1_N5166;
  tri   n7110;
  tri   n7113;
  tri   n7116;
  tri   n7055;
  tri   n7059;
  tri   n7062;
  tri   n7066;
  tri   n7070;
  tri   P1_N5157;
  tri   P1_N5156;
  tri   n7080;
  tri   n7081;
  tri   n7036;
  tri   n7041;
  tri   n7046;
  tri   n7048;
  tri   n7034;
  tri   P1_N4251;
  tri   P1_N4250;
  tri   P1_N4249;
  tri   P1_N4248;
  tri   P1_N4247;
  tri   P1_N4246;
  tri   P1_N4245;
  tri   P1_N4244;
  tri   P1_N4243;
  tri   P1_N4242;
  tri   P1_N4241;
  tri   P1_N4240;
  tri   P1_N4239;
  tri   P1_N4238;
  tri   P1_N4237;
  tri   P1_N4236;
  tri   P1_N4235;
  tri   P1_N4234;
  tri   P1_N4233;
  tri   P1_N4232;
  tri   P1_N4231;
  tri   P1_N4230;
  tri   P1_N4229;
  tri   P1_N4228;
  tri   P1_N4227;
  tri   P1_N4226;
  tri   P1_N4225;
  tri   P1_N4224;
  tri   P1_N4223;
  tri   P1_N4493;
  tri   P1_N4492;
  tri   P1_N4491;
  tri   P1_N4490;
  tri   P1_N4489;
  tri   P1_N4488;
  tri   P1_N4487;
  tri   P1_N4486;
  tri   P1_N4485;
  tri   P1_N4484;
  tri   P1_N4483;
  tri   P1_N4482;
  tri   P1_N4481;
  tri   P1_N4480;
  tri   P1_N4479;
  tri   P1_N4478;
  tri   P1_N4477;
  tri   P1_N4476;
  tri   P1_N4475;
  tri   P1_N4474;
  tri   P1_N4473;
  tri   P1_N4472;
  tri   P1_N4471;
  tri   P1_N4470;
  tri   P1_N4469;
  tri   P1_N4468;
  tri   P1_N4467;
  tri   P1_N4466;
  tri   P1_N4465;
  tri   P1_N5213;
  tri   P1_N5430;
  tri   P1_N5429;
  tri   P1_N5428;
  tri   P1_N5427;
  tri   P1_N5426;
  tri   P1_N5425;
  tri   P1_N5424;
  tri   P1_N5423;
  tri   P1_N5422;
  tri   P1_N5421;
  tri   P1_N5420;
  tri   P1_N5419;
  tri   P1_N5418;
  tri   P1_N5417;
  tri   P1_N5416;
  tri   P1_N5415;
  tri   P1_N5414;
  tri   P1_N5413;
  tri   P1_N5412;
  tri   P1_N5411;
  tri   P1_N5410;
  tri   P1_N5409;
  tri   P1_N5408;
  tri   P1_N5407;
  tri   P1_N5406;
  tri   P1_N5405;
  tri   P1_N5404;
  tri   P1_N5403;
  tri   P1_N5402;
  tri   P1_N5401;
  tri   P1_N5400;
  tri   P1_N5399;
  tri   P1_N5115;
  tri   P1_N5114;
  tri   P1_N5113;
  tri   P1_N5112;
  tri   P1_N5111;
  tri   P1_N5110;
  tri   P1_N5109;
  tri   P1_N5108;
  tri   P1_N5107;
  tri   P1_N5106;
  tri   P1_N5105;
  tri   P1_N5104;
  tri   P1_N5103;
  tri   P1_N5102;
  tri   P1_N5101;
  tri   P1_N5100;
  tri   P1_N5099;
  tri   P1_N5098;
  tri   P1_N5097;
  tri   P1_N5096;
  tri   P1_N5095;
  tri   P1_N5094;
  tri   n7273;
  tri   P1_N5092;
  tri   P1_N5091;
  tri   P1_N5090;
  tri   P1_N5089;
  tri   P1_N5088;
  tri   P1_N5087;
  tri   P1_N5086;
  tri   P1_N5085;
  tri   P1_N5084;
  tri   P1_N5281;
  tri   P1_N5362;
  tri   P1_N5431;
  tri   P2_N1514;
  tri   P2_N1513;
  tri   P2_N1512;
  tri   P2_N1511;
  tri   P2_N1510;
  tri   P2_N1509;
  tri   P2_N1508;
  tri   P2_N1507;
  tri   P2_N1506;
  tri   P2_N1505;
  tri   P2_N1504;
  tri   P2_N1503;
  tri   P2_N1502;
  tri   P2_N1501;
  tri   P2_N1500;
  tri   P2_N1499;
  tri   P2_N1498;
  tri   P2_N1497;
  tri   P2_N1496;
  tri   P2_N1495;
  tri   P2_N1494;
  tri   P2_N1493;
  tri   P2_N1492;
  tri   P2_N1491;
  tri   P2_N1490;
  tri   P2_N1489;
  tri   P2_N1488;
  tri   P2_N1487;
  tri   P2_N1486;
  tri   P2_N1756;
  tri   P2_N1755;
  tri   P2_N1754;
  tri   P2_N1753;
  tri   P2_N1752;
  tri   P2_N1751;
  tri   P2_N1750;
  tri   P2_N1749;
  tri   P2_N1748;
  tri   P2_N1747;
  tri   P2_N1746;
  tri   P2_N1745;
  tri   P2_N1744;
  tri   P2_N1743;
  tri   P2_N1742;
  tri   P2_N1741;
  tri   P2_N1740;
  tri   P2_N1739;
  tri   P2_N1738;
  tri   P2_N1737;
  tri   P2_N1736;
  tri   P2_N1735;
  tri   P2_N1734;
  tri   P2_N1733;
  tri   P2_N1732;
  tri   P2_N1731;
  tri   P2_N1730;
  tri   P2_N1729;
  tri   P2_N1728;
  tri   n7227;
  tri   P2_N1887;
  tri   P2_N1886;
  tri   P2_N1885;
  tri   P2_N1884;
  tri   P2_N1883;
  tri   P2_N1882;
  tri   P2_N1881;
  tri   P2_N1880;
  tri   P2_N1879;
  tri   P2_N1878;
  tri   P2_N1877;
  tri   P2_N1876;
  tri   P2_N1875;
  tri   P2_N1874;
  tri   P2_N1873;
  tri   P2_N1872;
  tri   P2_N1871;
  tri   P2_N1870;
  tri   P2_N1869;
  tri   P2_N1868;
  tri   P2_N1867;
  tri   P2_N1866;
  tri   P2_N1865;
  tri   P2_N1864;
  tri   P2_N1863;
  tri   P2_N1862;
  tri   P2_N1861;
  tri   P2_N1860;
  tri   P2_N1859;
  tri   P2_N2129;
  tri   P2_N2128;
  tri   P2_N2127;
  tri   P2_N2126;
  tri   P2_N2125;
  tri   P2_N2124;
  tri   P2_N2123;
  tri   P2_N2122;
  tri   P2_N2121;
  tri   P2_N2120;
  tri   P2_N2119;
  tri   P2_N2118;
  tri   P2_N2117;
  tri   P2_N2116;
  tri   P2_N2115;
  tri   P2_N2114;
  tri   P2_N2113;
  tri   P2_N2112;
  tri   P2_N2111;
  tri   P2_N2110;
  tri   P2_N2109;
  tri   P2_N2108;
  tri   P2_N2107;
  tri   P2_N2106;
  tri   P2_N2105;
  tri   P2_N2104;
  tri   P2_N2103;
  tri   P2_N2102;
  tri   P2_N2101;
  tri   P2_N5096;
  tri   n7162;
  tri   P2_N2260;
  tri   P2_N2259;
  tri   P2_N2258;
  tri   P2_N2257;
  tri   P2_N2256;
  tri   P2_N2255;
  tri   P2_N2254;
  tri   P2_N2253;
  tri   P2_N2252;
  tri   P2_N2251;
  tri   P2_N2250;
  tri   P2_N2249;
  tri   P2_N2248;
  tri   P2_N2247;
  tri   P2_N2246;
  tri   P2_N2245;
  tri   P2_N2244;
  tri   P2_N2243;
  tri   P2_N2242;
  tri   P2_N2241;
  tri   P2_N2240;
  tri   P2_N2239;
  tri   P2_N2238;
  tri   P2_N2237;
  tri   P2_N2236;
  tri   P2_N2235;
  tri   P2_N2234;
  tri   P2_N2233;
  tri   P2_N2232;
  tri   P2_N2502;
  tri   P2_N2501;
  tri   P2_N2500;
  tri   P2_N2499;
  tri   P2_N2498;
  tri   P2_N2497;
  tri   P2_N2496;
  tri   P2_N2495;
  tri   P2_N2494;
  tri   P2_N2493;
  tri   P2_N2492;
  tri   P2_N2491;
  tri   P2_N2490;
  tri   P2_N2489;
  tri   P2_N2488;
  tri   P2_N2487;
  tri   P2_N2486;
  tri   P2_N2485;
  tri   P2_N2484;
  tri   P2_N2483;
  tri   P2_N2482;
  tri   P2_N2481;
  tri   P2_N2480;
  tri   P2_N2479;
  tri   P2_N2478;
  tri   P2_N2477;
  tri   P2_N2476;
  tri   P2_N2475;
  tri   P2_N2474;
  tri   P1_N630;
  tri   P1_N658;
  tri   P1_N657;
  tri   P1_N656;
  tri   P1_N655;
  tri   P1_N654;
  tri   P1_N653;
  tri   P1_N652;
  tri   P1_N651;
  tri   P1_N650;
  tri   P1_N649;
  tri   P1_N648;
  tri   P1_N647;
  tri   P1_N646;
  tri   P1_N645;
  tri   P1_N644;
  tri   P1_N643;
  tri   P1_N642;
  tri   P1_N641;
  tri   P1_N640;
  tri   P1_N639;
  tri   P1_N638;
  tri   P1_N637;
  tri   P1_N636;
  tri   P1_N635;
  tri   P1_N634;
  tri   P1_N633;
  tri   P1_N632;
  tri   P1_N631;
  tri   n7274;
  tri   P1_N908;
  tri   P1_N907;
  tri   P1_N906;
  tri   P1_N905;
  tri   P1_N904;
  tri   P1_N903;
  tri   P1_N902;
  tri   P1_N901;
  tri   P1_N900;
  tri   P1_N899;
  tri   P1_N898;
  tri   P1_N897;
  tri   P1_N896;
  tri   P1_N895;
  tri   P1_N894;
  tri   P1_N893;
  tri   P1_N892;
  tri   P1_N891;
  tri   P1_N890;
  tri   P1_N889;
  tri   P1_N888;
  tri   P1_N887;
  tri   P1_N886;
  tri   P1_N885;
  tri   P1_N884;
  tri   P1_N883;
  tri   P1_N882;
  tri   P1_N881;
  tri   P1_N5170;
  tri   n7138;
  tri   n7124;
  tri   n7115;
  tri   n7106;
  tri   P1_N5167;
  tri   n7099;
  tri   P1_N5169;
  tri   P1_N5171;
  tri   P1_N5155;
  tri   n7075;
  tri   n4803;
  tri   P1_N5158;
  tri   n7119;
  tri   n7125;
  tri   n7130;
  tri   n7136;
  tri   n7144;
  tri   n7090;
  tri   n7092;
  tri   n7095;
  tri   n7098;
  tri   n7102;
  tri   n7105;
  tri   n7109;
  tri   n7112;
  tri   n7056;
  tri   n7063;
  tri   n7067;
  tri   n7071;
  tri   n7072;
  tri   n7076;
  tri   n7079;
  tri   n7082;
  tri   n7037;
  tri   n7043;
  tri   n7045;
  tri   n7051;
  tri   P1_N1640;
  tri   P1_N1639;
  tri   P1_N1638;
  tri   P1_N1637;
  tri   P1_N1636;
  tri   P1_N1635;
  tri   P1_N1634;
  tri   P1_N1633;
  tri   P1_N1632;
  tri   P1_N1631;
  tri   P1_N1630;
  tri   P1_N1629;
  tri   P1_N1628;
  tri   P1_N1627;
  tri   P1_N1626;
  tri   P1_N1625;
  tri   P1_N1624;
  tri   P1_N1623;
  tri   P1_N1622;
  tri   P1_N1621;
  tri   P1_N1620;
  tri   P1_N1619;
  tri   P1_N1618;
  tri   P1_N1617;
  tri   P1_N1616;
  tri   P1_N1615;
  tri   P1_N1614;
  tri   P1_N1613;
  tri   P1_N1612;
  tri   P1_N1882;
  tri   P1_N1881;
  tri   P1_N1880;
  tri   P1_N1879;
  tri   P1_N1878;
  tri   P1_N1877;
  tri   P1_N1876;
  tri   P1_N1875;
  tri   P1_N1874;
  tri   P1_N1873;
  tri   P1_N1872;
  tri   P1_N1871;
  tri   P1_N1870;
  tri   P1_N1869;
  tri   P1_N1868;
  tri   P1_N1867;
  tri   P1_N1866;
  tri   P1_N1865;
  tri   P1_N1864;
  tri   P1_N1863;
  tri   P1_N1862;
  tri   P1_N1861;
  tri   P1_N1860;
  tri   P1_N1859;
  tri   P1_N1858;
  tri   P1_N1857;
  tri   P1_N1856;
  tri   P1_N1855;
  tri   P1_N1854;
  tri   n7141;
  tri   P1_N5163;
  tri   n7058;
  tri   n7073;
  tri   P1_N2013;
  tri   P1_N2012;
  tri   P1_N2011;
  tri   P1_N2010;
  tri   P1_N2009;
  tri   P1_N2008;
  tri   P1_N2007;
  tri   P1_N2006;
  tri   P1_N2005;
  tri   P1_N2004;
  tri   P1_N2003;
  tri   P1_N2002;
  tri   P1_N2001;
  tri   P1_N2000;
  tri   P1_N1999;
  tri   P1_N1998;
  tri   P1_N1997;
  tri   P1_N1996;
  tri   P1_N1995;
  tri   P1_N1994;
  tri   P1_N1993;
  tri   P1_N1992;
  tri   P1_N1991;
  tri   P1_N1990;
  tri   P1_N1989;
  tri   P1_N1988;
  tri   P1_N1987;
  tri   P1_N1986;
  tri   P1_N1985;
  tri   P1_N2255;
  tri   P1_N2254;
  tri   P1_N2253;
  tri   P1_N2252;
  tri   P1_N2251;
  tri   P1_N2250;
  tri   P1_N2249;
  tri   P1_N2248;
  tri   P1_N2247;
  tri   P1_N2246;
  tri   P1_N2245;
  tri   P1_N2244;
  tri   P1_N2243;
  tri   P1_N2242;
  tri   P1_N2241;
  tri   P1_N2240;
  tri   P1_N2239;
  tri   P1_N2238;
  tri   P1_N2237;
  tri   P1_N2236;
  tri   P1_N2235;
  tri   P1_N2234;
  tri   P1_N2233;
  tri   P1_N2232;
  tri   P1_N2231;
  tri   P1_N2230;
  tri   P1_N2229;
  tri   P1_N2228;
  tri   P1_N2227;
  tri   P1_N5162;
  tri   P1_N5152;
  tri   P1_N2386;
  tri   P1_N2385;
  tri   P1_N2384;
  tri   P1_N2383;
  tri   P1_N2382;
  tri   P1_N2381;
  tri   P1_N2380;
  tri   P1_N2379;
  tri   P1_N2378;
  tri   P1_N2377;
  tri   P1_N2376;
  tri   P1_N2375;
  tri   P1_N2374;
  tri   P1_N2373;
  tri   P1_N2372;
  tri   P1_N2371;
  tri   P1_N2370;
  tri   P1_N2369;
  tri   P1_N2368;
  tri   P1_N2367;
  tri   P1_N2366;
  tri   P1_N2365;
  tri   P1_N2364;
  tri   P1_N2363;
  tri   P1_N2362;
  tri   P1_N2361;
  tri   P1_N2360;
  tri   P1_N2359;
  tri   P1_N2358;
  tri   P1_N2628;
  tri   P1_N2627;
  tri   P1_N2626;
  tri   P1_N2625;
  tri   P1_N2624;
  tri   P1_N2623;
  tri   P1_N2622;
  tri   P1_N2621;
  tri   P1_N2620;
  tri   P1_N2619;
  tri   P1_N2618;
  tri   P1_N2617;
  tri   P1_N2616;
  tri   P1_N2615;
  tri   P1_N2614;
  tri   P1_N2613;
  tri   P1_N2612;
  tri   P1_N2611;
  tri   P1_N2610;
  tri   P1_N2609;
  tri   P1_N2608;
  tri   P1_N2607;
  tri   P1_N2606;
  tri   P1_N2605;
  tri   P1_N2604;
  tri   P1_N2603;
  tri   P1_N2602;
  tri   P1_N2601;
  tri   P1_N2600;
  tri   P1_N5151;
  tri   P1_N5160;
  tri   P1_N2759;
  tri   P1_N2758;
  tri   P1_N2757;
  tri   P1_N2756;
  tri   P1_N2755;
  tri   P1_N2754;
  tri   P1_N2753;
  tri   P1_N2752;
  tri   P1_N2751;
  tri   P1_N2750;
  tri   P1_N2749;
  tri   P1_N2748;
  tri   P1_N2747;
  tri   P1_N2746;
  tri   P1_N2745;
  tri   P1_N2744;
  tri   P1_N2743;
  tri   P1_N2742;
  tri   P1_N2741;
  tri   P1_N2740;
  tri   P1_N2739;
  tri   P1_N2738;
  tri   P1_N2737;
  tri   P1_N2736;
  tri   P1_N2735;
  tri   P1_N2734;
  tri   P1_N2733;
  tri   P1_N2732;
  tri   P1_N2731;
  tri   P1_N3001;
  tri   P1_N3000;
  tri   P1_N2999;
  tri   P1_N2998;
  tri   P1_N2997;
  tri   P1_N2996;
  tri   P1_N2995;
  tri   P1_N2994;
  tri   P1_N2993;
  tri   P1_N2992;
  tri   P1_N2991;
  tri   P1_N2990;
  tri   P1_N2989;
  tri   P1_N2988;
  tri   P1_N2987;
  tri   P1_N2986;
  tri   P1_N2985;
  tri   P1_N2984;
  tri   P1_N2983;
  tri   P1_N2982;
  tri   P1_N2981;
  tri   P1_N2980;
  tri   P1_N2979;
  tri   P1_N2978;
  tri   P1_N2977;
  tri   P1_N2976;
  tri   P1_N2975;
  tri   P1_N2974;
  tri   P1_N2973;
  tri   n7122;
  tri   P1_N5159;
  tri   P1_N5161;
  tri   P1_N3132;
  tri   P1_N3131;
  tri   P1_N3130;
  tri   P1_N3129;
  tri   P1_N3128;
  tri   P1_N3127;
  tri   P1_N3126;
  tri   P1_N3125;
  tri   P1_N3124;
  tri   P1_N3123;
  tri   P1_N3122;
  tri   P1_N3121;
  tri   P1_N3120;
  tri   P1_N3119;
  tri   P1_N3118;
  tri   P1_N3117;
  tri   P1_N3116;
  tri   P1_N3115;
  tri   P1_N3114;
  tri   P1_N3113;
  tri   P1_N3112;
  tri   P1_N3111;
  tri   P1_N3110;
  tri   P1_N3109;
  tri   P1_N3108;
  tri   P1_N3107;
  tri   P1_N3106;
  tri   P1_N3105;
  tri   P1_N3104;
  tri   P1_N3374;
  tri   P1_N3373;
  tri   P1_N3372;
  tri   P1_N3371;
  tri   P1_N3370;
  tri   P1_N3369;
  tri   P1_N3368;
  tri   P1_N3367;
  tri   P1_N3366;
  tri   P1_N3365;
  tri   P1_N3364;
  tri   P1_N3363;
  tri   P1_N3362;
  tri   P1_N3361;
  tri   P1_N3360;
  tri   P1_N3359;
  tri   P1_N3358;
  tri   P1_N3357;
  tri   P1_N3356;
  tri   P1_N3355;
  tri   P1_N3354;
  tri   P1_N3353;
  tri   P1_N3352;
  tri   P1_N3351;
  tri   P1_N3350;
  tri   P1_N3349;
  tri   P1_N3348;
  tri   P1_N3347;
  tri   P1_N3346;
  tri   P1_N3505;
  tri   P1_N3504;
  tri   P1_N3503;
  tri   P1_N3502;
  tri   P1_N3501;
  tri   P1_N3500;
  tri   P1_N3499;
  tri   P1_N3498;
  tri   P1_N3497;
  tri   P1_N3496;
  tri   P1_N3495;
  tri   P1_N3494;
  tri   P1_N3493;
  tri   P1_N3492;
  tri   P1_N3491;
  tri   P1_N3490;
  tri   P1_N3489;
  tri   P1_N3488;
  tri   P1_N3487;
  tri   P1_N3486;
  tri   P1_N3485;
  tri   P1_N3484;
  tri   P1_N3483;
  tri   P1_N3482;
  tri   P1_N3481;
  tri   P1_N3480;
  tri   P1_N3479;
  tri   P1_N3478;
  tri   P1_N3477;
  tri   P1_N3747;
  tri   P1_N3746;
  tri   P1_N3745;
  tri   P1_N3744;
  tri   P1_N3743;
  tri   P1_N3742;
  tri   P1_N3741;
  tri   P1_N3740;
  tri   P1_N3739;
  tri   P1_N3738;
  tri   P1_N3737;
  tri   P1_N3736;
  tri   P1_N3735;
  tri   P1_N3734;
  tri   P1_N3733;
  tri   P1_N3732;
  tri   P1_N3731;
  tri   P1_N3730;
  tri   P1_N3729;
  tri   P1_N3728;
  tri   P1_N3727;
  tri   P1_N3726;
  tri   P1_N3725;
  tri   P1_N3724;
  tri   P1_N3723;
  tri   P1_N3722;
  tri   P1_N3721;
  tri   P1_N3720;
  tri   P1_N3719;
  tri   P1_N3878;
  tri   P1_N3877;
  tri   P1_N3876;
  tri   P1_N3875;
  tri   P1_N3874;
  tri   P1_N3873;
  tri   P1_N3872;
  tri   P1_N3871;
  tri   P1_N3870;
  tri   P1_N3869;
  tri   P1_N3868;
  tri   P1_N3867;
  tri   P1_N3866;
  tri   P1_N3865;
  tri   P1_N3864;
  tri   P1_N3863;
  tri   P1_N3862;
  tri   P1_N3861;
  tri   P1_N3860;
  tri   P1_N3859;
  tri   P1_N3858;
  tri   P1_N3857;
  tri   P1_N3856;
  tri   P1_N3855;
  tri   P1_N3854;
  tri   P1_N3853;
  tri   P1_N3852;
  tri   P1_N3851;
  tri   P1_N3850;
  tri   P1_N4120;
  tri   P1_N4119;
  tri   P1_N4118;
  tri   P1_N4117;
  tri   P1_N4116;
  tri   P1_N4115;
  tri   P1_N4114;
  tri   P1_N4113;
  tri   P1_N4112;
  tri   P1_N4111;
  tri   P1_N4110;
  tri   P1_N4109;
  tri   P1_N4108;
  tri   P1_N4107;
  tri   P1_N4106;
  tri   P1_N4105;
  tri   P1_N4104;
  tri   P1_N4103;
  tri   P1_N4102;
  tri   P1_N4101;
  tri   P1_N4100;
  tri   P1_N4099;
  tri   P1_N4098;
  tri   P1_N4097;
  tri   P1_N4096;
  tri   P1_N4095;
  tri   P1_N4094;
  tri   P1_N4093;
  tri   P1_N4092;
  tri   P2_N5099;
  tri   n7266;
  tri   P2_N2634;
  tri   P2_N2786;
  tri   P2_N2785;
  tri   P2_N2784;
  tri   P2_N2783;
  tri   P2_N2782;
  tri   P2_N2781;
  tri   P2_N2780;
  tri   P2_N2779;
  tri   P2_N2778;
  tri   P2_N2777;
  tri   P2_N2776;
  tri   P2_N2775;
  tri   P2_N2774;
  tri   P2_N2773;
  tri   P2_N2772;
  tri   P2_N2771;
  tri   P2_N2770;
  tri   P2_N2769;
  tri   P2_N2768;
  tri   P2_N2767;
  tri   P2_N2766;
  tri   P2_N2765;
  tri   P2_N2764;
  tri   P2_N2763;
  tri   P2_N2762;
  tri   P2_N2761;
  tri   P2_N2760;
  tri   P2_N2759;
  tri   P2_N2758;
  tri   P2_N2757;
  tri   P2_N3007;
  tri   P2_N3159;
  tri   P2_N3158;
  tri   P2_N3157;
  tri   P2_N3156;
  tri   P2_N3155;
  tri   P2_N3154;
  tri   P2_N3153;
  tri   P2_N3152;
  tri   P2_N3151;
  tri   P2_N3150;
  tri   P2_N3149;
  tri   P2_N3148;
  tri   P2_N3147;
  tri   P2_N3146;
  tri   P2_N3145;
  tri   P2_N3144;
  tri   P2_N3143;
  tri   P2_N3142;
  tri   P2_N3141;
  tri   P2_N3140;
  tri   P2_N3139;
  tri   P2_N3138;
  tri   P2_N3137;
  tri   P2_N3136;
  tri   P2_N3135;
  tri   P2_N3134;
  tri   P2_N3133;
  tri   P2_N3132;
  tri   P2_N3131;
  tri   P2_N3130;
  tri   P2_N3380;
  tri   P2_N3532;
  tri   P2_N3531;
  tri   P2_N3530;
  tri   P2_N3529;
  tri   P2_N3528;
  tri   P2_N3527;
  tri   P2_N3526;
  tri   P2_N3525;
  tri   P2_N3524;
  tri   P2_N3523;
  tri   P2_N3522;
  tri   P2_N3521;
  tri   P2_N3520;
  tri   P2_N3519;
  tri   P2_N3518;
  tri   P2_N3517;
  tri   P2_N3516;
  tri   P2_N3515;
  tri   P2_N3514;
  tri   P2_N3513;
  tri   P2_N3512;
  tri   P2_N3511;
  tri   P2_N3510;
  tri   P2_N3509;
  tri   P2_N3508;
  tri   P2_N3507;
  tri   P2_N3506;
  tri   P2_N3505;
  tri   P2_N3504;
  tri   P2_N3503;
  tri   P2_N3753;
  tri   P2_N3905;
  tri   P2_N3904;
  tri   P2_N3903;
  tri   P2_N3902;
  tri   P2_N3901;
  tri   P2_N3900;
  tri   P2_N3899;
  tri   P2_N3898;
  tri   P2_N3897;
  tri   P2_N3896;
  tri   P2_N3895;
  tri   P2_N3894;
  tri   P2_N3893;
  tri   P2_N3892;
  tri   P2_N3891;
  tri   P2_N3890;
  tri   P2_N3889;
  tri   P2_N3888;
  tri   P2_N3887;
  tri   P2_N3886;
  tri   P2_N3885;
  tri   P2_N3884;
  tri   P2_N3883;
  tri   P2_N3882;
  tri   P2_N3881;
  tri   P2_N3880;
  tri   P2_N3879;
  tri   P2_N3878;
  tri   P2_N3877;
  tri   P2_N3876;
  tri   P2_N4126;
  tri   P2_N4307;
  tri   P2_N4306;
  tri   P2_N4305;
  tri   P2_N4304;
  tri   P2_N4303;
  tri   P2_N4302;
  tri   P2_N4301;
  tri   P2_N4300;
  tri   P2_N4299;
  tri   P2_N4298;
  tri   P2_N4297;
  tri   P2_N4296;
  tri   P2_N4295;
  tri   P2_N4294;
  tri   P2_N4293;
  tri   P2_N4292;
  tri   P2_N4291;
  tri   P2_N4290;
  tri   P2_N4289;
  tri   P2_N4288;
  tri   P2_N4287;
  tri   P2_N4286;
  tri   P2_N4285;
  tri   P2_N4284;
  tri   P2_N4283;
  tri   P2_N4282;
  tri   P2_N4281;
  tri   P2_N4280;
  tri   P2_N4279;
  tri   P2_N4278;
  tri   P2_N5100;
  tri   P2_N4430;
  tri   n2562;
  tri   P2_N497;
  tri   P2_N4462;
  tri   P2_N4461;
  tri   P2_N4460;
  tri   P2_N4459;
  tri   P2_N4458;
  tri   P2_N4457;
  tri   P2_N4456;
  tri   P2_N4455;
  tri   P2_N4454;
  tri   P2_N4453;
  tri   P2_N4452;
  tri   P2_N4451;
  tri   P2_N4450;
  tri   P2_N4449;
  tri   P2_N4448;
  tri   P2_N4447;
  tri   P2_N4446;
  tri   P2_N4445;
  tri   P2_N4444;
  tri   P2_N4443;
  tri   P2_N4442;
  tri   P2_N4441;
  tri   P2_N4440;
  tri   P2_N4439;
  tri   P2_N4438;
  tri   P2_N4437;
  tri   P2_N4436;
  tri   P2_N4435;
  tri   P2_N4434;
  tri   P2_N4433;
  tri   P2_N4432;
  tri   P2_N4431;
  tri   P2_N5059;
  tri   P2_N5065;
  tri   P2_N5062;
  tri   n7265;
  tri   P2_N5015;
  tri   n18245;
  tri   n9565;
  tri   n9569;
  tri   n9573;
  tri   n9577;
  tri   n9581;
  tri   n9585;
  tri   n9589;
  tri   n9593;
  tri   n9597;
  tri   n9601;
  tri   n9605;
  tri   n9609;
  tri   n9613;
  tri   n9617;
  tri   n9621;
  tri   n9625;
  tri   n9629;
  tri   n9318;
  tri   n9329;
  tri   n18209;
  tri   n9417;
  tri   n9421;
  tri   n9425;
  tri   n9429;
  tri   n9433;
  tri   n9437;
  tri   n9441;
  tri   n9445;
  tri   n9449;
  tri   n9453;
  tri   n9457;
  tri   n9461;
  tri   n9465;
  tri   n9469;
  tri   n9473;
  tri   n9477;
  tri   n9481;
  tri   n9485;
  tri   n9489;
  tri   n18347;
  tri   n6688;
  tri   n10137;
  tri   n10133;
  tri   n10141;
  tri   n10369;
  tri   n10183;
  tri   n10377;
  tri   n10191;
  tri   n6719;
  tri   n6608;
  tri   n6609;
  tri   n6610;
  tri   n6611;
  tri   n6612;
  tri   n6613;
  tri   n6614;
  tri   n6615;
  tri   n6616;
  tri   n6617;
  tri   n6607;
  tri   n6606;
  tri   n6605;
  tri   n6604;
  tri   n6603;
  tri   n6602;
  tri   n6601;
  tri   n6600;
  tri   n6599;
  tri   n6598;
  tri   n6597;
  tri   n6596;
  tri   n6595;
  tri   P2_N133;
  tri   P2_N132;
  tri   P2_N131;
  tri   P2_N130;
  tri   P2_N129;
  tri   P2_N128;
  tri   P2_N127;
  tri   P2_N126;
  tri   P2_N125;
  tri   P2_N124;
  tri   P2_N123;
  tri   P2_N122;
  tri   P2_N121;
  tri   P2_N120;
  tri   P2_N119;
  tri   P2_N118;
  tri   P2_N117;
  tri   P2_N116;
  tri   P2_N115;
  tri   P2_N114;
  tri   P2_N113;
  tri   P2_N112;
  tri   P2_N111;
  tri   P2_N110;
  tri   P2_N109;
  tri   P2_N108;
  tri   P2_N107;
  tri   P2_N106;
  tri   P2_N105;
  tri   P2_N104;
  tri   P2_N103;
  tri   n6771;
  tri   P2_N345;
  tri   P2_N346;
  tri   P2_N347;
  tri   P2_N348;
  tri   P2_N349;
  tri   P2_N350;
  tri   P2_N351;
  tri   P2_N352;
  tri   P2_N353;
  tri   P2_N354;
  tri   P2_N355;
  tri   P2_N356;
  tri   P2_N357;
  tri   P2_N358;
  tri   P2_N359;
  tri   P2_N360;
  tri   P2_N361;
  tri   P2_N363;
  tri   n10112;
  tri   n18907;
  tri   n18909;
  tri   n18911;
  tri   n18913;
  tri   n18915;
  tri   n18917;
  tri   n18919;
  tri   n18921;
  tri   n18923;
  tri   n18925;
  tri   n10250;
  tri   n18927;
  tri   n18929;
  tri   n18931;
  tri   n18933;
  tri   n18935;
  tri   n18937;
  tri   n9838;
  tri   n116;
  tri   n117;
  tri   n118;
  tri   n119;
  tri   n120;
  tri   n121;
  tri   n122;
  tri   n123;
  tri   n124;
  tri   n125;
  tri   n126;
  tri   n127;
  tri   n128;
  tri   n129;
  tri   n130;
  tri   n131;
  tri   n132;
  tri   n133;
  tri   n134;
  tri   n135;
  tri   n10117;
  tri   n18963;
  tri   n18965;
  tri   n18967;
  tri   n18969;
  tri   n18971;
  tri   n18973;
  tri   n18975;
  tri   n18977;
  tri   n18979;
  tri   n18981;
  tri   n18983;
  tri   n18985;
  tri   n18987;
  tri   n18989;
  tri   n18991;
  tri   n18993;
  tri   n18995;
  tri   n9843;
  tri   n95;
  tri   n96;
  tri   n97;
  tri   n98;
  tri   n99;
  tri   n100;
  tri   n101;
  tri   n102;
  tri   n103;
  tri   n104;
  tri   n105;
  tri   n106;
  tri   n107;
  tri   n108;
  tri   n109;
  tri   n110;
  tri   n111;
  tri   n112;
  tri   n113;
  tri   n114;
  tri   n9349;
  tri   n9353;
  tri   n9357;
  tri   n9361;
  tri   n9365;
  tri   n9369;
  tri   n9373;
  tri   n9377;
  tri   n9381;
  tri   n9501;
  tri   n9505;
  tri   n9509;
  tri   n9513;
  tri   n9517;
  tri   n9521;
  tri   n9525;
  tri   n9529;
  tri   n9533;
  tri   n9537;
  tri   n9541;
  tri   n9545;
  tri   n9549;
  tri   n9553;
  tri   n9557;
  tri   n9397;
  tri   n6684;
  tri   P2_N394;
  tri   P2_N393;
  tri   P2_N392;
  tri   P2_N391;
  tri   P2_N390;
  tri   P2_N389;
  tri   P2_N388;
  tri   P2_N387;
  tri   P2_N386;
  tri   P2_N385;
  tri   P2_N384;
  tri   P2_N383;
  tri   P2_N382;
  tri   P2_N381;
  tri   P2_N380;
  tri   P2_N379;
  tri   P2_N378;
  tri   P2_N377;
  tri   P2_N376;
  tri   P2_N375;
  tri   P2_N374;
  tri   P2_N373;
  tri   P2_N372;
  tri   P2_N371;
  tri   P2_N370;
  tri   P2_N369;
  tri   P2_N368;
  tri   n9345;
  tri   n10103;
  tri   n10095;
  tri   n9935;
  tri   n9939;
  tri   n9943;
  tri   n9947;
  tri   n9951;
  tri   n9955;
  tri   n9959;
  tri   n9963;
  tri   n9967;
  tri   n9971;
  tri   n9975;
  tri   n9979;
  tri   n9983;
  tri   n9987;
  tri   n9991;
  tri   n9995;
  tri   n9999;
  tri   n10003;
  tri   n10007;
  tri   n9871;
  tri   n9875;
  tri   n9879;
  tri   n9883;
  tri   n9887;
  tri   n9891;
  tri   n9895;
  tri   n9899;
  tri   n9333;
  tri   n9385;
  tri   N70;
  tri   N69;
  tri   N68;
  tri   N67;
  tri   N66;
  tri   N65;
  tri   N64;
  tri   N63;
  tri   N62;
  tri   N61;
  tri   N60;
  tri   N59;
  tri   N58;
  tri   N57;
  tri   N56;
  tri   N55;
  tri   N54;
  tri   N53;
  tri   N52;
  tri   N51;
  tri   N50;
  tri   N49;
  tri   N48;
  tri   N47;
  tri   N46;
  tri   N45;
  tri   N44;
  tri   N43;
  tri   N42;
  tri   N41;
  tri   N40;
  tri   N39;
  tri   P2_N1515;
  tri   P2_N1667;
  tri   P2_N1666;
  tri   P2_N1665;
  tri   P2_N1664;
  tri   P2_N1663;
  tri   P2_N1662;
  tri   P2_N1661;
  tri   P2_N1660;
  tri   P2_N1659;
  tri   P2_N1658;
  tri   P2_N1657;
  tri   P2_N1656;
  tri   P2_N1655;
  tri   P2_N1654;
  tri   P2_N1653;
  tri   P2_N1652;
  tri   P2_N1651;
  tri   P2_N1650;
  tri   P2_N1649;
  tri   P2_N1648;
  tri   P2_N1647;
  tri   P2_N1646;
  tri   P2_N1645;
  tri   P2_N1644;
  tri   P2_N1643;
  tri   P2_N1642;
  tri   P2_N1641;
  tri   P2_N1640;
  tri   P2_N1639;
  tri   P2_N1638;
  tri   P2_N1888;
  tri   P2_N2040;
  tri   P2_N2039;
  tri   P2_N2038;
  tri   P2_N2037;
  tri   P2_N2036;
  tri   P2_N2035;
  tri   P2_N2034;
  tri   P2_N2033;
  tri   P2_N2032;
  tri   P2_N2031;
  tri   P2_N2030;
  tri   P2_N2029;
  tri   P2_N2028;
  tri   P2_N2027;
  tri   P2_N2026;
  tri   P2_N2025;
  tri   P2_N2024;
  tri   P2_N2023;
  tri   P2_N2022;
  tri   P2_N2021;
  tri   P2_N2020;
  tri   P2_N2019;
  tri   P2_N2018;
  tri   P2_N2017;
  tri   P2_N2016;
  tri   P2_N2015;
  tri   P2_N2014;
  tri   P2_N2013;
  tri   P2_N2012;
  tri   P2_N2011;
  tri   P2_N2261;
  tri   P2_N2413;
  tri   P2_N2412;
  tri   P2_N2411;
  tri   P2_N2410;
  tri   P2_N2409;
  tri   P2_N2408;
  tri   P2_N2407;
  tri   P2_N2406;
  tri   P2_N2405;
  tri   P2_N2404;
  tri   P2_N2403;
  tri   P2_N2402;
  tri   P2_N2401;
  tri   P2_N2400;
  tri   P2_N2399;
  tri   P2_N2398;
  tri   P2_N2397;
  tri   P2_N2396;
  tri   P2_N2395;
  tri   P2_N2394;
  tri   P2_N2393;
  tri   P2_N2392;
  tri   P2_N2391;
  tri   P2_N2390;
  tri   P2_N2389;
  tri   P2_N2388;
  tri   P2_N2387;
  tri   P2_N2386;
  tri   P2_N2385;
  tri   P2_N2384;
  tri   n7146;
  tri   P1_N5177;
  tri   P1_N5174;
  tri   P1_N5154;
  tri   P1_N5153;
  tri   P1_N2387;
  tri   P1_N2539;
  tri   P1_N2538;
  tri   P1_N2537;
  tri   P1_N2536;
  tri   P1_N2535;
  tri   P1_N2534;
  tri   P1_N2533;
  tri   P1_N2532;
  tri   P1_N2531;
  tri   P1_N2530;
  tri   P1_N2529;
  tri   P1_N2528;
  tri   P1_N2527;
  tri   P1_N2526;
  tri   P1_N2525;
  tri   P1_N2524;
  tri   P1_N2523;
  tri   P1_N2522;
  tri   P1_N2521;
  tri   P1_N2520;
  tri   P1_N2519;
  tri   P1_N2518;
  tri   P1_N2517;
  tri   P1_N2516;
  tri   P1_N2515;
  tri   P1_N2514;
  tri   P1_N2513;
  tri   P1_N2512;
  tri   P1_N2511;
  tri   P1_N2510;
  tri   P1_N2760;
  tri   P1_N2912;
  tri   P1_N2911;
  tri   P1_N2910;
  tri   P1_N2909;
  tri   P1_N2908;
  tri   P1_N2907;
  tri   P1_N2906;
  tri   P1_N2905;
  tri   P1_N2904;
  tri   P1_N2903;
  tri   P1_N2902;
  tri   P1_N2901;
  tri   P1_N2900;
  tri   P1_N2899;
  tri   P1_N2898;
  tri   P1_N2897;
  tri   P1_N2896;
  tri   P1_N2895;
  tri   P1_N2894;
  tri   P1_N2893;
  tri   P1_N2892;
  tri   P1_N2891;
  tri   P1_N2890;
  tri   P1_N2889;
  tri   P1_N2888;
  tri   P1_N2887;
  tri   P1_N2886;
  tri   P1_N2885;
  tri   P1_N2884;
  tri   P1_N2883;
  tri   P1_N3133;
  tri   P1_N3285;
  tri   P1_N3284;
  tri   P1_N3283;
  tri   P1_N3282;
  tri   P1_N3281;
  tri   P1_N3280;
  tri   P1_N3279;
  tri   P1_N3278;
  tri   P1_N3277;
  tri   P1_N3276;
  tri   P1_N3275;
  tri   P1_N3274;
  tri   P1_N3273;
  tri   P1_N3272;
  tri   P1_N3271;
  tri   P1_N3270;
  tri   P1_N3269;
  tri   P1_N3268;
  tri   P1_N3267;
  tri   P1_N3266;
  tri   P1_N3265;
  tri   P1_N3264;
  tri   P1_N3263;
  tri   P1_N3262;
  tri   P1_N3261;
  tri   P1_N3260;
  tri   P1_N3259;
  tri   P1_N3258;
  tri   P1_N3257;
  tri   P1_N3256;
  tri   P1_N3506;
  tri   P1_N3658;
  tri   P1_N3657;
  tri   P1_N3656;
  tri   P1_N3655;
  tri   P1_N3654;
  tri   P1_N3653;
  tri   P1_N3652;
  tri   P1_N3651;
  tri   P1_N3650;
  tri   P1_N3649;
  tri   P1_N3648;
  tri   P1_N3647;
  tri   P1_N3646;
  tri   P1_N3645;
  tri   P1_N3644;
  tri   P1_N3643;
  tri   P1_N3642;
  tri   P1_N3641;
  tri   P1_N3640;
  tri   P1_N3639;
  tri   P1_N3638;
  tri   P1_N3637;
  tri   P1_N3636;
  tri   P1_N3635;
  tri   P1_N3634;
  tri   P1_N3633;
  tri   P1_N3632;
  tri   P1_N3631;
  tri   P1_N3630;
  tri   P1_N3629;
  tri   P1_N3879;
  tri   P1_N4031;
  tri   P1_N4030;
  tri   P1_N4029;
  tri   P1_N4028;
  tri   P1_N4027;
  tri   P1_N4026;
  tri   P1_N4025;
  tri   P1_N4024;
  tri   P1_N4023;
  tri   P1_N4022;
  tri   P1_N4021;
  tri   P1_N4020;
  tri   P1_N4019;
  tri   P1_N4018;
  tri   P1_N4017;
  tri   P1_N4016;
  tri   P1_N4015;
  tri   P1_N4014;
  tri   P1_N4013;
  tri   P1_N4012;
  tri   P1_N4011;
  tri   P1_N4010;
  tri   P1_N4009;
  tri   P1_N4008;
  tri   P1_N4007;
  tri   P1_N4006;
  tri   P1_N4005;
  tri   P1_N4004;
  tri   P1_N4003;
  tri   P1_N4002;
  tri   P1_N4252;
  tri   P1_N4404;
  tri   P1_N4403;
  tri   P1_N4402;
  tri   P1_N4401;
  tri   P1_N4400;
  tri   P1_N4399;
  tri   P1_N4398;
  tri   P1_N4397;
  tri   P1_N4396;
  tri   P1_N4395;
  tri   P1_N4394;
  tri   P1_N4393;
  tri   P1_N4392;
  tri   P1_N4391;
  tri   P1_N4390;
  tri   P1_N4389;
  tri   P1_N4388;
  tri   P1_N4387;
  tri   P1_N4386;
  tri   P1_N4385;
  tri   P1_N4384;
  tri   P1_N4383;
  tri   P1_N4382;
  tri   P1_N4381;
  tri   P1_N4380;
  tri   P1_N4379;
  tri   P1_N4378;
  tri   P1_N4377;
  tri   P1_N4376;
  tri   P1_N4375;
  tri   P1_N5178;
  tri   P1_N4556;
  tri   n4469;
  tri   P1_N497;
  tri   P1_N4588;
  tri   P1_N4587;
  tri   P1_N4586;
  tri   P1_N4585;
  tri   P1_N4584;
  tri   P1_N4583;
  tri   P1_N4582;
  tri   P1_N4581;
  tri   P1_N4580;
  tri   P1_N4579;
  tri   P1_N4578;
  tri   P1_N4577;
  tri   P1_N4576;
  tri   P1_N4575;
  tri   P1_N4574;
  tri   P1_N4573;
  tri   P1_N4572;
  tri   P1_N4571;
  tri   P1_N4570;
  tri   P1_N4569;
  tri   P1_N4568;
  tri   P1_N4567;
  tri   P1_N4566;
  tri   P1_N4565;
  tri   P1_N4564;
  tri   P1_N4563;
  tri   P1_N4562;
  tri   P1_N4561;
  tri   P1_N4560;
  tri   P1_N4559;
  tri   P1_N4558;
  tri   P1_N4557;
  tri   P1_N5137;
  tri   P1_N5143;
  tri   P1_N5140;
  tri   n7145;
  tri   P1_N5093;
  tri   n18695;
  tri   n6708;
  tri   n10129;
  tri   n10125;
  tri   n10145;
  tri   n10373;
  tri   n10187;
  tri   n10381;
  tri   n10195;
  tri   n6637;
  tri   n6638;
  tri   n6639;
  tri   n6640;
  tri   n6641;
  tri   n6642;
  tri   n6643;
  tri   n6644;
  tri   n6645;
  tri   n6646;
  tri   n6647;
  tri   n6636;
  tri   n6635;
  tri   n6634;
  tri   n6633;
  tri   n6632;
  tri   n6631;
  tri   n6630;
  tri   n6629;
  tri   n6628;
  tri   n6627;
  tri   n6626;
  tri   n6625;
  tri   n6624;
  tri   P1_N133;
  tri   P1_N132;
  tri   P1_N131;
  tri   P1_N130;
  tri   P1_N129;
  tri   P1_N128;
  tri   P1_N127;
  tri   P1_N126;
  tri   P1_N125;
  tri   P1_N124;
  tri   P1_N123;
  tri   P1_N122;
  tri   P1_N121;
  tri   P1_N120;
  tri   P1_N119;
  tri   P1_N118;
  tri   P1_N117;
  tri   P1_N116;
  tri   P1_N115;
  tri   P1_N114;
  tri   P1_N113;
  tri   P1_N112;
  tri   P1_N111;
  tri   P1_N110;
  tri   P1_N109;
  tri   P1_N108;
  tri   P1_N107;
  tri   P1_N106;
  tri   P1_N105;
  tri   P1_N104;
  tri   P1_N103;
  tri   P1_N345;
  tri   P1_N346;
  tri   P1_N349;
  tri   P1_N347;
  tri   P1_N350;
  tri   P1_N348;
  tri   P1_N353;
  tri   P1_N351;
  tri   P1_N354;
  tri   P1_N352;
  tri   P1_N357;
  tri   P1_N355;
  tri   P1_N358;
  tri   P1_N356;
  tri   P1_N359;
  tri   P1_N363;
  tri   P1_N361;
  tri   P1_N360;
  tri   P1_N344;
  tri   n6773;
  tri   n6770;
  tri   n6766;
  tri   n6762;
  tri   n6767;
  tri   n6763;
  tri   n6758;
  tri   n6754;
  tri   n6759;
  tri   n6755;
  tri   n6750;
  tri   n6746;
  tri   n6751;
  tri   n6747;
  tri   n6744;
  tri   n6742;
  tri   n6734;
  tri   n6732;
  tri   n6730;
  tri   n9493;
  tri   n9693;
  tri   n9697;
  tri   n9701;
  tri   n9705;
  tri   n9709;
  tri   n9713;
  tri   n9717;
  tri   n9721;
  tri   n9725;
  tri   n9729;
  tri   n9733;
  tri   n9737;
  tri   n9741;
  tri   n9745;
  tri   n9749;
  tri   n9753;
  tri   n9757;
  tri   n9761;
  tri   n981;
  tri   n192;
  tri   n193;
  tri   n194;
  tri   n195;
  tri   n196;
  tri   n197;
  tri   n198;
  tri   n199;
  tri   n200;
  tri   n201;
  tri   n202;
  tri   n203;
  tri   n204;
  tri   n205;
  tri   n206;
  tri   n207;
  tri   n208;
  tri   n209;
  tri   n210;
  tri   n211;
  tri   n9497;
  tri   n9765;
  tri   n9769;
  tri   n9773;
  tri   n9777;
  tri   n9781;
  tri   n9785;
  tri   n9789;
  tri   n9793;
  tri   n9797;
  tri   n9801;
  tri   n9805;
  tri   n9809;
  tri   n9813;
  tri   n9817;
  tri   n9821;
  tri   n9825;
  tri   n9829;
  tri   n9833;
  tri   n920;
  tri   n171;
  tri   n172;
  tri   n173;
  tri   n174;
  tri   n175;
  tri   n176;
  tri   n177;
  tri   n178;
  tri   n179;
  tri   n180;
  tri   n181;
  tri   n182;
  tri   n183;
  tri   n184;
  tri   n185;
  tri   n186;
  tri   n187;
  tri   n188;
  tri   n189;
  tri   n190;
  tri   n9341;
  tri   n10107;
  tri   n10099;
  tri   n10019;
  tri   n10023;
  tri   n10027;
  tri   n10031;
  tri   n10035;
  tri   n10039;
  tri   n10043;
  tri   n10047;
  tri   n10051;
  tri   n10055;
  tri   n10059;
  tri   n10063;
  tri   n10067;
  tri   n10071;
  tri   n10075;
  tri   n10079;
  tri   n10083;
  tri   n10087;
  tri   n10091;
  tri   n9903;
  tri   n9907;
  tri   n9911;
  tri   n9915;
  tri   n9919;
  tri   n9923;
  tri   n9927;
  tri   n9931;
  tri   n9337;
  tri   n9389;
  tri   N38;
  tri   N37;
  tri   N36;
  tri   N35;
  tri   N34;
  tri   N33;
  tri   N32;
  tri   N31;
  tri   N30;
  tri   N29;
  tri   N28;
  tri   N27;
  tri   N26;
  tri   N25;
  tri   N24;
  tri   N23;
  tri   N22;
  tri   N21;
  tri   N20;
  tri   N19;
  tri   N18;
  tri   N17;
  tri   N16;
  tri   N15;
  tri   N14;
  tri   N13;
  tri   N12;
  tri   N11;
  tri   N10;
  tri   N9;
  tri   N8;
  tri   N7;
  tri   P1_N661;
  tri   P1_N660;
  tri   P1_N659;
  tri   P1_N815;
  tri   P1_N814;
  tri   P1_N813;
  tri   P1_N812;
  tri   P1_N811;
  tri   P1_N810;
  tri   P1_N809;
  tri   P1_N808;
  tri   P1_N807;
  tri   P1_N806;
  tri   P1_N805;
  tri   P1_N804;
  tri   P1_N803;
  tri   P1_N802;
  tri   P1_N801;
  tri   P1_N800;
  tri   P1_N799;
  tri   P1_N798;
  tri   P1_N797;
  tri   P1_N796;
  tri   P1_N795;
  tri   P1_N794;
  tri   P1_N793;
  tri   P1_N792;
  tri   P1_N791;
  tri   P1_N790;
  tri   P1_N789;
  tri   P1_N788;
  tri   P1_N787;
  tri   P1_N786;
  tri   P1_N785;
  tri   n18451;
  tri   n9633;
  tri   n9401;
  tri   n9637;
  tri   n9405;
  tri   n9641;
  tri   n9409;
  tri   n9645;
  tri   n9413;
  tri   n9649;
  tri   n9661;
  tri   n9851;
  tri   n9665;
  tri   n9855;
  tri   n9669;
  tri   n9859;
  tri   n9673;
  tri   n9863;
  tri   n9677;
  tri   n9867;
  tri   n9681;
  tri   n10011;
  tri   n9685;
  tri   n10015;
  tri   n9689;
  tri   n9657;
  tri   n6594;
  tri   P1_N393;
  tri   P1_N392;
  tri   P1_N391;
  tri   P1_N390;
  tri   P1_N389;
  tri   P1_N388;
  tri   P1_N387;
  tri   P1_N386;
  tri   P1_N385;
  tri   P1_N384;
  tri   P1_N383;
  tri   P1_N382;
  tri   P1_N381;
  tri   P1_N380;
  tri   P1_N379;
  tri   P1_N378;
  tri   P1_N377;
  tri   P1_N376;
  tri   P1_N375;
  tri   P1_N374;
  tri   P1_N373;
  tri   P1_N372;
  tri   P1_N371;
  tri   P1_N370;
  tri   P1_N369;
  tri   P1_N368;
  tri   P1_N1641;
  tri   P1_N1793;
  tri   P1_N1792;
  tri   P1_N1791;
  tri   P1_N1790;
  tri   P1_N1789;
  tri   P1_N1788;
  tri   P1_N1787;
  tri   P1_N1786;
  tri   P1_N1785;
  tri   P1_N1784;
  tri   P1_N1783;
  tri   P1_N1782;
  tri   P1_N1781;
  tri   P1_N1780;
  tri   P1_N1779;
  tri   P1_N1778;
  tri   P1_N1777;
  tri   P1_N1776;
  tri   P1_N1775;
  tri   P1_N1774;
  tri   P1_N1773;
  tri   P1_N1772;
  tri   P1_N1771;
  tri   P1_N1770;
  tri   P1_N1769;
  tri   P1_N1768;
  tri   P1_N1767;
  tri   P1_N1766;
  tri   P1_N1765;
  tri   P1_N1764;
  tri   P1_N2014;
  tri   P1_N2166;
  tri   P1_N2165;
  tri   P1_N2164;
  tri   P1_N2163;
  tri   P1_N2162;
  tri   P1_N2161;
  tri   P1_N2160;
  tri   P1_N2159;
  tri   P1_N2158;
  tri   P1_N2157;
  tri   P1_N2156;
  tri   P1_N2155;
  tri   P1_N2154;
  tri   P1_N2153;
  tri   P1_N2152;
  tri   P1_N2151;
  tri   P1_N2150;
  tri   P1_N2149;
  tri   P1_N2148;
  tri   P1_N2147;
  tri   P1_N2146;
  tri   P1_N2145;
  tri   P1_N2144;
  tri   P1_N2143;
  tri   P1_N2142;
  tri   P1_N2141;
  tri   P1_N2140;
  tri   P1_N2139;
  tri   P1_N2138;
  tri   P1_N2137;
  tri   clock_G1B2I1_1;
  tri   clock_G1B1I2_1;
  tri   clock_G1B1I1_1;
  tri   clock_G1B2I38_1;
  tri   clock_G1B2I37_1;
  tri   clock_G1B2I34_1;
  tri   clock_G1B2I33_1;
  tri   clock_G1B2I36_1;
  tri   clock_G1B1I3_1;
  tri   clock_G1B2I32_1;
  tri   clock_G1B2I27_1;
  tri   clock_G1B2I35_1;
  tri   clock_G1B2I15_1;
  tri   clock_G1B2I31_1;
  tri   clock_G1B2I9_1;
  tri   clock_G1B2I30_1;
  tri   clock_G1B2I29_1;
  tri   clock_G1B2I17_1;
  tri   clock_G1B2I21_1;
  tri   clock_G1B2I23_1;
  tri   clock_G1B2I28_1;
  tri   clock_G1B2I14_1;
  tri   clock_G1B2I26_1;
  tri   clock_G1B2I18_1;
  tri   clock_G1B2I12_1;
  tri   clock_G1B2I13_1;
  tri   clock_G1B2I24_1;
  tri   clock_G1B2I25_1;
  tri   clock_G1B2I3_1;
  tri   clock_G1B2I22_1;
  tri   clock_G1B2I20_1;
  tri   clock_G1B2I19_1;
  tri   clock_G1B2I8_1;
  tri   clock_G1B2I16_1;
  tri   clock_G1B2I7_1;
  tri   clock_G1B2I11_1;
  tri   clock_G1B2I2_1;
  tri   clock_G1B2I4_1;
  tri   clock_G1B2I6_1;
  tri   clock_G1B2I5_1;
  tri   clock_G1B2I10_1;
  tri   P2_N5470;
  tri   n6729;
  tri   n6931;
  tri   n7460;
  tri   n6967;
  tri   P2_N294;
  tri   n6705;
  tri   n7480;
  tri   n7462;
  tri   n7007;
  tri   n7479;
  tri   n6693;
  tri   n4169;
  tri   n7580;
  tri   n7582;
  tri   n18293;
  tri   n6580;
  tri   n2166;
  tri   n7501;
  tri   n6573;
  tri   n18762;
  tri   n6589;
  tri   n18345;
  tri   n18343;
  tri   n18341;
  tri   n6715;
  tri   n6699;
  tri   n6685;
  tri   n6703;
  tri   n6716;
  tri   n6687;
  tri   n6706;
  tri   n6704;
  tri   n6712;
  tri   n6694;
  tri   n19025;
  tri   n6690;
  tri   n6718;
  tri   n6692;
  tri   n19009;
  tri   n6710;
  tri   n6737;
  tri   n6736;
  tri   n6739;
  tri   N5;
  tri   n6621;
  tri   n18465;
  tri   n6681;
  tri   n18819;
  tri   n4480;
  tri   n4615;
  tri   n4616;
  tri   n2569;
  tri   n2660;
  tri   n2661;
  tri   n6622;
  tri   n18459;
  tri   n6682;
  tri   n18817;
  tri   P1_N583;
  tri   n4157;
  tri   n4158;
  tri   n2693;
  tri   n2153;
  tri   n2154;
  tri   n4804;
  tri   n4805;
  tri   n2920;
  tri   n2921;
  tri   n6683;
  tri   n18815;
  tri   n6623;
  tri   n18455;
  tri   P1_N5147;
  tri   n7281;
  tri   n2205;
  tri   n7311;
  tri   P2_N914;
  tri   n7015;
  tri   n7314;
  tri   n4202;
  tri   n2199;
  tri   n7315;
  tri   n2202;
  tri   n7313;
  tri   n7316;
  tri   n4199;
  tri   n2196;
  tri   n7317;
  tri   n7318;
  tri   n4196;
  tri   n7319;
  tri   n2193;
  tri   n7322;
  tri   n4190;
  tri   n7320;
  tri   n4193;
  tri   n2187;
  tri   n7323;
  tri   n2190;
  tri   n7321;
  tri   n7324;
  tri   n4187;
  tri   n2184;
  tri   n7325;
  tri   n2181;
  tri   n7327;
  tri   n7326;
  tri   n4184;
  tri   n7328;
  tri   n4181;
  tri   n6592;
  tri   n18207;
  tri   n6620;
  tri   n18285;
  tri   n18287;
  tri   n6619;
  tri   n6593;
  tri   n18205;
  tri   n7271;
  tri   P1_N536;
  tri   n7272;
  tri   P2_N536;
  tri   n6895;
  tri   n7483;
  tri   n6999;
  tri   P2_N584;
  tri   n7485;
  tri   n6837;
  tri   n6896;
  tri   n6838;
  tri   n6910;
  tri   n6332;
  tri   n6333;
  tri   n7458;
  tri   P1_N584;
  tri   n6996;
  tri   n7484;
  tri   n6847;
  tri   n6869;
  tri   n6809;
  tri   n6893;
  tri   n7482;
  tri   n6897;
  tri   n6899;
  tri   n6848;
  tri   n6915;
  tri   n6870;
  tri   n6808;
  tri   n6807;
  tri   n6854;
  tri   n7459;
  tri   n6883;
  tri   n6898;
  tri   n6900;
  tri   n6916;
  tri   n6917;
  tri   n6819;
  tri   n2992;
  tri   n7354;
  tri   n2934;
  tri   n5709;
  tri   n7356;
  tri   n7355;
  tri   n4022;
  tri   n7376;
  tri   n7375;
  tri   n3796;
  tri   n7378;
  tri   n7377;
  tri   n3710;
  tri   n7380;
  tri   n7379;
  tri   n3624;
  tri   n7382;
  tri   n7381;
  tri   n3512;
  tri   n7384;
  tri   n7383;
  tri   n3403;
  tri   n7386;
  tri   n7385;
  tri   n3299;
  tri   n7388;
  tri   n7387;
  tri   n3213;
  tri   n7390;
  tri   n7389;
  tri   n3105;
  tri   n7392;
  tri   n7391;
  tri   n3019;
  tri   n7394;
  tri   n7393;
  tri   n2069;
  tri   n7395;
  tri   n7396;
  tri   n1466;
  tri   P2_N4244;
  tri   P2_N5509;
  tri   n1485;
  tri   P1_N3434;
  tri   P1_N5581;
  tri   n6891;
  tri   P1_N292;
  tri   P1_N293;
  tri   n6949;
  tri   P2_N292;
  tri   n6851;
  tri   n6835;
  tri   n6834;
  tri   n7486;
  tri   n6815;
  tri   P1_N506;
  tri   n6618;
  tri   P2_N506;
  tri   n6591;
  tri   P1_N2878;
  tri   P1_N3062;
  tri   P1_N2880;
  tri   P1_N3031;
  tri   P1_N3251;
  tri   P1_N3435;
  tri   P1_N3253;
  tri   P1_N3404;
  tri   P1_N3624;
  tri   P1_N3808;
  tri   P1_N3626;
  tri   P1_N3777;
  tri   P1_N3997;
  tri   P1_N4181;
  tri   P1_N3999;
  tri   P1_N4150;
  tri   P1_N4370;
  tri   P1_N4554;
  tri   P1_N4372;
  tri   P1_N4523;
  tri   P1_N6685;
  tri   P1_N6686;
  tri   P1_N6688;
  tri   P1_N779;
  tri   P1_N969;
  tri   P1_N781;
  tri   P1_N938;
  tri   P1_N1250;
  tri   P1_N1315;
  tri   P1_N1252;
  tri   P1_N1284;
  tri   P1_N1759;
  tri   P1_N1943;
  tri   P1_N1761;
  tri   P1_N1912;
  tri   P1_N2132;
  tri   P1_N2316;
  tri   P1_N2134;
  tri   P1_N2285;
  tri   P1_N2505;
  tri   P1_N2689;
  tri   P1_N2507;
  tri   P1_N2658;
  tri   P2_N6610;
  tri   P2_N1633;
  tri   P2_N1817;
  tri   P2_N1635;
  tri   P2_N1786;
  tri   P2_N2006;
  tri   P2_N2190;
  tri   P2_N2008;
  tri   P2_N2159;
  tri   P2_N2379;
  tri   P2_N2563;
  tri   P2_N2381;
  tri   P2_N2532;
  tri   P2_N2752;
  tri   P2_N2936;
  tri   P2_N2754;
  tri   P2_N2905;
  tri   P2_N3125;
  tri   P2_N3309;
  tri   P2_N3127;
  tri   P2_N3278;
  tri   P2_N3498;
  tri   P2_N3682;
  tri   P2_N3500;
  tri   P2_N3651;
  tri   P2_N3871;
  tri   P2_N4055;
  tri   P2_N3873;
  tri   P2_N4024;
  tri   P2_N4428;
  tri   P2_N6607;
  tri   P2_N6608;
  tri   n6940;
  tri   P2_N778;
  tri   P2_N843;
  tri   P2_N780;
  tri   P2_N812;
  tri   P2_N1124;
  tri   P2_N1189;
  tri   P2_N1126;
  tri   P2_N1158;
  tri   n6979;
  tri   P1_N294;
  tri   n6824;
  tri   n6823;
  tri   n6843;
  tri   n6781;
  tri   P2_N291;
  tri   n6829;
  tri   n4510;
  tri   n7400;
  tri   n7399;
  tri   P1_N5282;
  tri   P1_N1505;
  tri   P1_N1570;
  tri   P1_N1507;
  tri   P1_N1539;
  tri   P2_N5204;
  tri   P2_N1379;
  tri   P2_N1444;
  tri   P2_N1381;
  tri   P2_N1413;
  tri   n6980;
  tri   n6972;
  tri   n6802;
  tri   n6860;
  tri   P1_N291;
  tri   n6855;
  tri   n14523;
  tri   n14763;
  tri   n11310;
  tri   n11550;
  tri   P1_N4752;
  tri   P1_N4817;
  tri   P1_N4754;
  tri   P1_N4786;
  tri   P2_N4626;
  tri   P2_N4691;
  tri   n6934;
  tri   n6975;
  tri   n7461;
  tri   n6954;
  tri   n6977;
  tri   n6966;
  tri   n6984;
  tri   n6583;
  tri   n6584;
  tri   n2168;
  tri   P2_N499;
  tri   n4164;
  tri   n4356;
  tri   n6585;
  tri   n4171;
  tri   P1_N499;
  tri   n6582;
  tri   n6586;
  tri   n7455;
  tri   n7449;
  tri   n7456;
  tri   n7448;
  tri   n598;
  tri   n2459;
  tri   n599;
  tri   n2452;
  tri   n480;
  tri   n4366;
  tri   n481;
  tri   n6579;
  tri   n6570;
  tri   n7285;
  tri   P2_N5419;
  tri   P1_N5554;
  tri   n7031;
  tri   n7284;
  tri   P1_N5497;
  tri   n6572;
  tri   n7457;
  tri   n6568;
  tri   n7540;
  tri   n6577;
  tri   n6578;
  tri   n7454;
  tri   n7478;
  tri   n7539;
  tri   n6576;
  tri   n7536;
  tri   n7535;
  tri   n7549;
  tri   n7553;
  tri   n7554;
  tri   n7555;
  tri   n6569;
  tri   n6574;
  tri   n7584;
  tri   n7581;
  tri   n7585;
  tri   n7586;
  tri   n7583;
  tri   n7505;
  tri   n7504;
  tri   n7506;
  tri   n6713;
  tri   n6787;
  tri   n7487;
  tri   n6943;
  tri   n6932;
  tri   P2_N293;
  tri   n6937;
  tri   n6946;
  tri   n7606;
  tri   n7605;
  tri   n7604;
  tri   n7603;
  tri   n7602;
  tri   n7601;
  tri   n7600;
  tri   n7599;
  tri   n7598;
  tri   n7597;
  tri   n7596;
  tri   n7595;
  tri   n7594;
  tri   n7593;
  tri   n7592;
  tri   n7591;
  tri   n7590;
  tri   n7589;
  tri   n7588;
  tri   n7587;
  tri   n7579;
  tri   n7578;
  tri   n7577;
  tri   n7576;
  tri   n7575;
  tri   n7574;
  tri   n7573;
  tri   n6571;
  tri   n7572;
  tri   n7453;
  tri   n7571;
  tri   n7570;
  tri   n7569;
  tri   n7568;
  tri   n7567;
  tri   n7566;
  tri   n7565;
  tri   n7564;
  tri   n7563;
  tri   n7562;
  tri   n7561;
  tri   n7560;
  tri   n7559;
  tri   n7558;
  tri   n7557;
  tri   n7548;
  tri   n7547;
  tri   n7546;
  tri   n7545;
  tri   n7544;
  tri   n7543;
  tri   n7542;
  tri   n7541;
  tri   n7538;
  tri   n6560;
  tri   n7537;
  tri   n7534;
  tri   n7533;
  tri   n7532;
  tri   n7531;
  tri   n7530;
  tri   n7529;
  tri   n7528;
  tri   n7527;
  tri   n7526;
  tri   n7525;
  tri   n6556;
  tri   n7524;
  tri   n7523;
  tri   n7522;
  tri   n7521;
  tri   n7520;
  tri   n7519;
  tri   n7518;
  tri   n7517;
  tri   n7516;
  tri   n7515;
  tri   n7514;
  tri   n7513;
  tri   n6567;
  tri   n7512;
  tri   n7511;
  tri   n7510;
  tri   n7509;
  tri   n7508;
  tri   n7507;
  tri   n6561;
  tri   n7502;
  tri   n7500;
  tri   n7499;
  tri   n7498;
  tri   n7497;
  tri   n7496;
  tri   n7495;
  tri   n7494;
  tri   n7493;
  tri   n7492;
  tri   n7491;
  tri   n7490;
  tri   n7489;
  tri   n6382;
  tri   n6383;
  tri   n7488;
  tri   n6384;
  tri   n6385;
  tri   n6334;
  tri   n6335;
  tri   n7481;
  tri   n6566;
  tri   n7477;
  tri   n7476;
  tri   n7475;
  tri   n6575;
  tri   n7474;
  tri   n7473;
  tri   n7472;
  tri   n6563;
  tri   n7471;
  tri   n7470;
  tri   n7469;
  tri   n7468;
  tri   n7467;
  tri   n7466;
  tri   n7465;
  tri   n7464;
  tri   n1502;
  tri   n7463;
  tri   n1481;
  tri   n6338;
  tri   n6339;
  tri   n6388;
  tri   n6389;
  tri   n7550;
  tri   n7452;
  tri   n7451;
  tri   n7450;
  tri   n7556;
  tri   n7503;
  tri   n7552;
  tri   n7551;
  tri   n2586;
  tri   n2587;
  tri   n7447;
  tri   n2579;
  tri   n2580;
  tri   n7446;
  tri   n4499;
  tri   n4498;
  tri   n7445;
  tri   n4491;
  tri   n4490;
  tri   n7444;
  tri   P1_N5433;
  tri   n4367;
  tri   n7443;
  tri   P2_N5355;
  tri   n2460;
  tri   n7442;
  tri   P1_N663;
  tri   n7441;
  tri   P1_N664;
  tri   n7440;
  tri   P1_N666;
  tri   n7439;
  tri   P1_N668;
  tri   n7438;
  tri   P1_N669;
  tri   n7437;
  tri   P1_N670;
  tri   n7436;
  tri   P1_N671;
  tri   n7435;
  tri   P1_N672;
  tri   n7434;
  tri   P1_N673;
  tri   n7433;
  tri   P1_N674;
  tri   n7432;
  tri   P1_N675;
  tri   n7431;
  tri   P1_N676;
  tri   n7430;
  tri   P1_N677;
  tri   n7429;
  tri   P1_N678;
  tri   n7428;
  tri   P1_N679;
  tri   n7427;
  tri   P1_N680;
  tri   n7426;
  tri   P1_N681;
  tri   n7425;
  tri   P1_N682;
  tri   n7424;
  tri   n7422;
  tri   n7409;
  tri   n7423;
  tri   n6784;
  tri   n7412;
  tri   n7411;
  tri   n7421;
  tri   n7413;
  tri   n7420;
  tri   n7408;
  tri   n7407;
  tri   n7419;
  tri   n7410;
  tri   n7418;
  tri   n7406;
  tri   n7405;
  tri   n7417;
  tri   n7404;
  tri   n7416;
  tri   P2_N245;
  tri   n6381;
  tri   n7415;
  tri   P1_N245;
  tri   n6331;
  tri   n7414;
  tri   n6793;
  tri   n6963;
  tri   n6857;
  tri   n6956;
  tri   n7403;
  tri   P1_N5755;
  tri   P1_N5756;
  tri   n7398;
  tri   P2_N4561;
  tri   n7402;
  tri   n7401;
  tri   P2_N5677;
  tri   P2_N5678;
  tri   P1_N6683;
  tri   P1_N6684;
  tri   P1_N6681;
  tri   P1_N6682;
  tri   P2_N6605;
  tri   P2_N6606;
  tri   P2_N4178;
  tri   n7397;
  tri   P2_N5899;
  tri   P2_N5900;
  tri   P2_N5901;
  tri   P2_N5902;
  tri   P2_N6477;
  tri   P2_N6478;
  tri   P2_N6475;
  tri   P2_N6476;
  tri   P2_N6413;
  tri   P2_N6414;
  tri   P2_N6411;
  tri   P2_N6412;
  tri   P2_N6349;
  tri   P2_N6350;
  tri   P2_N6347;
  tri   P2_N6348;
  tri   P2_N6285;
  tri   P2_N6286;
  tri   P2_N6283;
  tri   P2_N6284;
  tri   P2_N6221;
  tri   P2_N6222;
  tri   P2_N6219;
  tri   P2_N6220;
  tri   P2_N6157;
  tri   P2_N6158;
  tri   P2_N6155;
  tri   P2_N6156;
  tri   P2_N6093;
  tri   P2_N6094;
  tri   P2_N6091;
  tri   P2_N6092;
  tri   P2_N6029;
  tri   P2_N6030;
  tri   P2_N6027;
  tri   P2_N6028;
  tri   P2_N5965;
  tri   P2_N5966;
  tri   P2_N5963;
  tri   P2_N5964;
  tri   P1_N5979;
  tri   P1_N5980;
  tri   P1_N5977;
  tri   P1_N5978;
  tri   n7374;
  tri   P1_N6619;
  tri   P1_N6620;
  tri   n7373;
  tri   P1_N6617;
  tri   P1_N6618;
  tri   n7372;
  tri   P1_N6555;
  tri   P1_N6556;
  tri   n7371;
  tri   P1_N6553;
  tri   P1_N6554;
  tri   n7370;
  tri   P1_N6491;
  tri   P1_N6492;
  tri   n7369;
  tri   P1_N6489;
  tri   P1_N6490;
  tri   n7368;
  tri   P1_N6427;
  tri   P1_N6428;
  tri   n7367;
  tri   P1_N6425;
  tri   P1_N6426;
  tri   n7366;
  tri   P1_N6363;
  tri   P1_N6364;
  tri   n7365;
  tri   P1_N6361;
  tri   P1_N6362;
  tri   n7364;
  tri   P1_N6299;
  tri   P1_N6300;
  tri   n7363;
  tri   P1_N6297;
  tri   P1_N6298;
  tri   n7362;
  tri   P1_N6235;
  tri   P1_N6236;
  tri   n7361;
  tri   P1_N6233;
  tri   P1_N6234;
  tri   n7360;
  tri   P1_N6171;
  tri   P1_N6172;
  tri   n7359;
  tri   P1_N6169;
  tri   P1_N6170;
  tri   n7358;
  tri   P1_N6107;
  tri   P1_N6108;
  tri   n7357;
  tri   P1_N6105;
  tri   P1_N6106;
  tri   P1_N6043;
  tri   P1_N6044;
  tri   P1_N6041;
  tri   P1_N6042;
  tri   P2_N6541;
  tri   P2_N6542;
  tri   n7353;
  tri   P2_N5631;
  tri   P2_N5632;
  tri   n7352;
  tri   P1_N5709;
  tri   P1_N5710;
  tri   n7351;
  tri   P1_N5653;
  tri   P1_N5654;
  tri   n7350;
  tri   P2_N5575;
  tri   P2_N5576;
  tri   n9310;
  tri   n7349;
  tri   n9314;
  tri   n7348;
  tri   n7347;
  tri   n7346;
  tri   n7336;
  tri   n7345;
  tri   n7335;
  tri   n7344;
  tri   n7339;
  tri   n7343;
  tri   n7338;
  tri   n7342;
  tri   n7341;
  tri   n7340;
  tri   n6415;
  tri   n6414;
  tri   n6418;
  tri   n6417;
  tri   n7331;
  tri   n7337;
  tri   n6365;
  tri   n6364;
  tri   n6368;
  tri   n6367;
  tri   n7333;
  tri   n7334;
  tri   n6401;
  tri   n6400;
  tri   n6404;
  tri   n6403;
  tri   n7332;
  tri   n6351;
  tri   n6350;
  tri   n6354;
  tri   n6353;
  tri   n7330;
  tri   n7052;
  tri   P2_N5069;
  tri   n7147;
  tri   P1_N662;
  tri   n7019;
  tri   n7012;
  tri   n7013;
  tri   n6810;
  tri   n17734;
  tri   n2657;
  tri   n14521;
  tri   n6779;
  tri   n6782;
  tri   n6813;
  tri   n6842;
  tri   n6827;
  tri   n6907;
  tri   n6923;
  tri   n6922;
  tri   n6921;
  tri   n6874;
  tri   n6878;
  tri   n6941;
  tri   n6969;
  tri   n7309;
  tri   P2_N5485;
  tri   n6564;
  tri   n6562;
  tri   n6559;
  tri   n6557;
  tri   n6565;
  tri   n6558;
  tri   n2178;
  tri   n7329;
  tri   n7312;
  tri   n4205;
  tri   n4208;
  tri   n7310;
  tri   P2_N5486;
  tri   n7303;
  tri   P1_N5563;
  tri   n7299;
  tri   P1_N5564;
  tri   n7295;
  tri   n7291;
  tri   P2_N5484;
  tri   P1_N5562;
  tri   n7287;
  tri   n7279;
  tri   P2_N5476;
  tri   n7270;
  tri   n7029;
  tri   n7028;
  tri   n7027;
  tri   n7026;
  tri   n7024;
  tri   n7022;
  tri   n7023;
  tri   n7021;
  tri   n7016;
  tri   n7011;
  tri   n7010;
  tri   n7009;
  tri   n7006;
  tri   n6993;
  tri   n6992;
  tri   n11309;
  tri   n14522;
  tri   n6986;
  tri   n6981;
  tri   n6982;
  tri   n6976;
  tri   n6974;
  tri   n6970;
  tri   n6961;
  tri   n6962;
  tri   n6959;
  tri   n6957;
  tri   n6958;
  tri   n6955;
  tri   n6952;
  tri   n6948;
  tri   n6942;
  tri   n6928;
  tri   n6927;
  tri   n6926;
  tri   n6901;
  tri   n6920;
  tri   n6919;
  tri   n6906;
  tri   n6904;
  tri   n6894;
  tri   n6892;
  tri   n6890;
  tri   n6887;
  tri   n6888;
  tri   n6886;
  tri   n6884;
  tri   n6881;
  tri   n6882;
  tri   n6871;
  tri   n6872;
  tri   n6867;
  tri   n6865;
  tri   n6866;
  tri   n6864;
  tri   n6861;
  tri   n6862;
  tri   n6856;
  tri   n6852;
  tri   n6836;
  tri   n6831;
  tri   n6832;
  tri   n6830;
  tri   n6828;
  tri   n6825;
  tri   n6822;
  tri   n6820;
  tri   n6818;
  tri   n6816;
  tri   n6812;
  tri   n6803;
  tri   n6804;
  tri   n6794;
  tri   n6792;
  tri   n6790;
  tri   n6789;
  tri   n6775;
  tri   n6786;
  tri   n6780;
  tri   n6776;
  tri   P1_N362;
  tri   n6725;
  tri   P1_N5548;
  tri   n19001;
  tri   n6714;
  tri   n6702;
  tri   n6700;
  tri   n6698;
  tri   n6696;
  tri   n6686;
  tri   n18813;
  tri   n18643;
  tri   n18645;
  tri   n18647;
  tri   n18649;
  tri   n18651;
  tri   n18653;
  tri   n18655;
  tri   n18657;
  tri   n18659;
  tri   n18661;
  tri   n18663;
  tri   n18671;
  tri   n18673;
  tri   n18675;
  tri   n18677;
  tri   n18679;
  tri   n18681;
  tri   n18683;
  tri   n18685;
  tri   n18687;
  tri   n18689;
  tri   n18691;
  tri   n18693;
  tri   n18297;
  tri   n18299;
  tri   n18301;
  tri   n18303;
  tri   n18305;
  tri   n18307;
  tri   n18309;
  tri   n18311;
  tri   n18313;
  tri   n18315;
  tri   n18323;
  tri   n18325;
  tri   n18327;
  tri   n18329;
  tri   n18331;
  tri   n18333;
  tri   n18335;
  tri   n18337;
  tri   n18339;
  tri   n6590;
  tri   n6588;
  tri   n5945;
  tri   n5946;
  tri   n4150;
  tri   n5948;
  tri   n5949;
  tri   n4153;
  tri   n5951;
  tri   n5952;
  tri   n4156;
  tri   n5942;
  tri   n5943;
  tri   n4147;
  tri   n5939;
  tri   n5940;
  tri   n4144;
  tri   n5936;
  tri   n5937;
  tri   n4141;
  tri   n5933;
  tri   n5934;
  tri   n4138;
  tri   n3886;
  tri   n3887;
  tri   n2044;
  tri   n6348;
  tri   n6347;
  tri   n3881;
  tri   n3882;
  tri   n2041;
  tri   n3963;
  tri   n3964;
  tri   P2_N925;
  tri   n3861;
  tri   n3862;
  tri   n2029;
  tri   n3856;
  tri   n3857;
  tri   n2026;
  tri   n3951;
  tri   n3952;
  tri   P2_N928;
  tri   n3851;
  tri   n3852;
  tri   n2023;
  tri   n3947;
  tri   n3948;
  tri   P2_N929;
  tri   n3846;
  tri   n3847;
  tri   n2020;
  tri   n3841;
  tri   n3842;
  tri   n2017;
  tri   n3836;
  tri   n3837;
  tri   n2014;
  tri   n5894;
  tri   n5895;
  tri   n4099;
  tri   n3826;
  tri   n3827;
  tri   n2008;
  tri   n6398;
  tri   n6397;
  tri   n5924;
  tri   n5925;
  tri   n4129;
  tri   n4112;
  tri   n4115;
  tri   n4118;
  tri   n4121;
  tri   n4124;
  tri   n4127;
  tri   n4136;
  tri   n2024;
  tri   n2027;
  tri   n2030;
  tri   n5921;
  tri   n5922;
  tri   n4126;
  tri   n5918;
  tri   n5919;
  tri   n4123;
  tri   n4375;
  tri   n4376;
  tri   n2468;
  tri   n2469;
  tri   n5915;
  tri   n5916;
  tri   n4120;
  tri   n5912;
  tri   n5913;
  tri   n4117;
  tri   n5623;
  tri   n5511;
  tri   n5425;
  tri   n5316;
  tri   n5212;
  tri   n5104;
  tri   n5018;
  tri   n4932;
  tri   n4818;
  tri   n5909;
  tri   n5910;
  tri   n4114;
  tri   n1474;
  tri   P2_N5497;
  tri   n5906;
  tri   n5907;
  tri   n4111;
  tri   n5903;
  tri   n5904;
  tri   n4108;
  tri   n3831;
  tri   n3832;
  tri   n2011;
  tri   n18952;
  tri   n18953;
  tri   n18954;
  tri   n18955;
  tri   n18956;
  tri   n18957;
  tri   n18958;
  tri   n18959;
  tri   n18960;
  tri   n18961;
  tri   n18998;
  tri   n18999;
  tri   n19002;
  tri   n19003;
  tri   n19004;
  tri   n19005;
  tri   n19006;
  tri   n19007;
  tri   n19010;
  tri   n19011;
  tri   n19012;
  tri   n19013;
  tri   n19014;
  tri   n19015;
  tri   n19016;
  tri   n19017;
  tri   n19018;
  tri   n19019;
  tri   n19020;
  tri   n19021;
  tri   n19022;
  tri   n19023;
  tri   n18766;
  tri   n18767;
  tri   n18768;
  tri   n18769;
  tri   n18770;
  tri   n18771;
  tri   n18772;
  tri   n18773;
  tri   n18774;
  tri   n18775;
  tri   n18776;
  tri   n18777;
  tri   n18778;
  tri   n18779;
  tri   n18780;
  tri   n18781;
  tri   n18782;
  tri   n18783;
  tri   n18784;
  tri   n18785;
  tri   n18786;
  tri   n18787;
  tri   n18788;
  tri   n18789;
  tri   n18790;
  tri   n18791;
  tri   n18792;
  tri   n18793;
  tri   n18794;
  tri   n18795;
  tri   n18796;
  tri   n18797;
  tri   n18798;
  tri   n18799;
  tri   n18800;
  tri   n18801;
  tri   n18802;
  tri   n18803;
  tri   n18804;
  tri   n18805;
  tri   n18806;
  tri   n18807;
  tri   n18808;
  tri   n18809;
  tri   n18810;
  tri   n18811;
  tri   n18820;
  tri   n18821;
  tri   n18822;
  tri   n18823;
  tri   n18824;
  tri   n18825;
  tri   n18826;
  tri   n18827;
  tri   n18828;
  tri   n18829;
  tri   n18830;
  tri   n18831;
  tri   n18832;
  tri   n18833;
  tri   n18834;
  tri   n18835;
  tri   n18836;
  tri   n18837;
  tri   n18838;
  tri   n18839;
  tri   n18840;
  tri   n18841;
  tri   n18842;
  tri   n18843;
  tri   n18844;
  tri   n18845;
  tri   n18846;
  tri   n18847;
  tri   n18848;
  tri   n18849;
  tri   n18850;
  tri   n18851;
  tri   n18852;
  tri   n18853;
  tri   n18854;
  tri   n18855;
  tri   n18856;
  tri   n18857;
  tri   n18858;
  tri   n18859;
  tri   n18860;
  tri   n18861;
  tri   n18862;
  tri   n18863;
  tri   n18864;
  tri   n18865;
  tri   n18866;
  tri   n18867;
  tri   n18868;
  tri   n18869;
  tri   n18870;
  tri   n18871;
  tri   n18872;
  tri   n18873;
  tri   n18874;
  tri   n18875;
  tri   n18876;
  tri   n18877;
  tri   n18878;
  tri   n18879;
  tri   n18880;
  tri   n18881;
  tri   n18882;
  tri   n18883;
  tri   n18884;
  tri   n18885;
  tri   n18886;
  tri   n18887;
  tri   n18888;
  tri   n18889;
  tri   n18890;
  tri   n18891;
  tri   n18892;
  tri   n18893;
  tri   n18894;
  tri   n18895;
  tri   n18896;
  tri   n18897;
  tri   n18898;
  tri   n18899;
  tri   n18900;
  tri   n18901;
  tri   n18902;
  tri   n18903;
  tri   n18904;
  tri   n18905;
  tri   n18940;
  tri   n18941;
  tri   n18942;
  tri   n18943;
  tri   n18944;
  tri   n18945;
  tri   n18946;
  tri   n18947;
  tri   n18948;
  tri   n18949;
  tri   n18950;
  tri   n18951;
  tri   n18580;
  tri   n18581;
  tri   n18582;
  tri   n18583;
  tri   n18584;
  tri   n18585;
  tri   n18586;
  tri   n18587;
  tri   n18588;
  tri   n18589;
  tri   n18590;
  tri   n18591;
  tri   n18592;
  tri   n18593;
  tri   n18594;
  tri   n18595;
  tri   n18596;
  tri   n18597;
  tri   n18598;
  tri   n18599;
  tri   n18600;
  tri   n18601;
  tri   n18602;
  tri   n18603;
  tri   n18604;
  tri   n18605;
  tri   n18606;
  tri   n18607;
  tri   n18608;
  tri   n18609;
  tri   n18610;
  tri   n18611;
  tri   n18612;
  tri   n18613;
  tri   n18614;
  tri   n18615;
  tri   n18616;
  tri   n18617;
  tri   n18618;
  tri   n18619;
  tri   n18620;
  tri   n18621;
  tri   n18622;
  tri   n18623;
  tri   n18624;
  tri   n18625;
  tri   n18626;
  tri   n18627;
  tri   n18628;
  tri   n18629;
  tri   n18630;
  tri   n18631;
  tri   n18632;
  tri   n18633;
  tri   n18634;
  tri   n18635;
  tri   n18636;
  tri   n18637;
  tri   n18638;
  tri   n18639;
  tri   n18640;
  tri   n18641;
  tri   n18664;
  tri   n18665;
  tri   n18666;
  tri   n18667;
  tri   n18668;
  tri   n18669;
  tri   n18696;
  tri   n18697;
  tri   n18698;
  tri   n18699;
  tri   n18700;
  tri   n18701;
  tri   n18702;
  tri   n18703;
  tri   n18704;
  tri   n18705;
  tri   n18706;
  tri   n18707;
  tri   n18708;
  tri   n18709;
  tri   n18710;
  tri   n18711;
  tri   n18712;
  tri   n18713;
  tri   n18714;
  tri   n18715;
  tri   n18716;
  tri   n18717;
  tri   n18718;
  tri   n18719;
  tri   n18720;
  tri   n18721;
  tri   n18722;
  tri   n18723;
  tri   n18724;
  tri   n18725;
  tri   n18726;
  tri   n18727;
  tri   n18728;
  tri   n18729;
  tri   n18730;
  tri   n18731;
  tri   n18732;
  tri   n18733;
  tri   n18734;
  tri   n18735;
  tri   n18736;
  tri   n18737;
  tri   n18738;
  tri   n18739;
  tri   n18740;
  tri   n18741;
  tri   n18742;
  tri   n18743;
  tri   n18744;
  tri   n18745;
  tri   n18746;
  tri   n18747;
  tri   n18748;
  tri   n18749;
  tri   n18750;
  tri   n18751;
  tri   n18752;
  tri   n18753;
  tri   n18754;
  tri   n18755;
  tri   n18756;
  tri   n18757;
  tri   n18758;
  tri   n18759;
  tri   n18760;
  tri   n18761;
  tri   n18763;
  tri   n18764;
  tri   n18765;
  tri   n18394;
  tri   n18395;
  tri   n18396;
  tri   n18397;
  tri   n18398;
  tri   n18399;
  tri   n18400;
  tri   n18401;
  tri   n18402;
  tri   n18403;
  tri   n18404;
  tri   n18405;
  tri   n18406;
  tri   n18407;
  tri   n18408;
  tri   n18409;
  tri   n18410;
  tri   n18411;
  tri   n18412;
  tri   n18413;
  tri   n18414;
  tri   n18415;
  tri   n18416;
  tri   n18417;
  tri   n18418;
  tri   n18419;
  tri   n18420;
  tri   n18421;
  tri   n18422;
  tri   n18423;
  tri   n18424;
  tri   n18425;
  tri   n18426;
  tri   n18427;
  tri   n18428;
  tri   n18429;
  tri   n18430;
  tri   n18431;
  tri   n18432;
  tri   n18433;
  tri   n18434;
  tri   n18435;
  tri   n18436;
  tri   n18437;
  tri   n18438;
  tri   n18439;
  tri   n18440;
  tri   n18441;
  tri   n18442;
  tri   n18443;
  tri   n18444;
  tri   n18445;
  tri   n18446;
  tri   n18447;
  tri   n18448;
  tri   n18449;
  tri   n18452;
  tri   n18453;
  tri   n18456;
  tri   n18457;
  tri   n18460;
  tri   n18461;
  tri   n18462;
  tri   n18463;
  tri   n18466;
  tri   n18467;
  tri   n18468;
  tri   n18469;
  tri   n18470;
  tri   n18471;
  tri   n18472;
  tri   n18473;
  tri   n18474;
  tri   n18475;
  tri   n18476;
  tri   n18477;
  tri   n18478;
  tri   n18479;
  tri   n18480;
  tri   n18481;
  tri   n18482;
  tri   n18483;
  tri   n18484;
  tri   n18485;
  tri   n18486;
  tri   n18487;
  tri   n18488;
  tri   n18489;
  tri   n18490;
  tri   n18491;
  tri   n18492;
  tri   n18493;
  tri   n18494;
  tri   n18495;
  tri   n18496;
  tri   n18497;
  tri   n18498;
  tri   n18499;
  tri   n18500;
  tri   n18501;
  tri   n18502;
  tri   n18503;
  tri   n18504;
  tri   n18505;
  tri   n18506;
  tri   n18507;
  tri   n18508;
  tri   n18509;
  tri   n18510;
  tri   n18511;
  tri   n18512;
  tri   n18513;
  tri   n18514;
  tri   n18515;
  tri   n18516;
  tri   n18517;
  tri   n18518;
  tri   n18519;
  tri   n18520;
  tri   n18521;
  tri   n18522;
  tri   n18523;
  tri   n18524;
  tri   n18525;
  tri   n18526;
  tri   n18527;
  tri   n18528;
  tri   n18529;
  tri   n18530;
  tri   n18531;
  tri   n18532;
  tri   n18533;
  tri   n18534;
  tri   n18535;
  tri   n18536;
  tri   n18537;
  tri   n18538;
  tri   n18539;
  tri   n18540;
  tri   n18541;
  tri   n18542;
  tri   n18543;
  tri   n18544;
  tri   n18545;
  tri   n18546;
  tri   n18547;
  tri   n18548;
  tri   n18549;
  tri   n18550;
  tri   n18551;
  tri   n18552;
  tri   n18553;
  tri   n18554;
  tri   n18555;
  tri   n18556;
  tri   n18557;
  tri   n18558;
  tri   n18559;
  tri   n18560;
  tri   n18561;
  tri   n18562;
  tri   n18563;
  tri   n18564;
  tri   n18565;
  tri   n18566;
  tri   n18567;
  tri   n18568;
  tri   n18569;
  tri   n18570;
  tri   n18571;
  tri   n18572;
  tri   n18573;
  tri   n18574;
  tri   n18575;
  tri   n18576;
  tri   n18577;
  tri   n18578;
  tri   n18579;
  tri   n18211;
  tri   n18212;
  tri   n18213;
  tri   n18214;
  tri   n18215;
  tri   n18216;
  tri   n18217;
  tri   n18218;
  tri   n18219;
  tri   n18220;
  tri   n18221;
  tri   n18222;
  tri   n18223;
  tri   n18224;
  tri   n18225;
  tri   n18226;
  tri   n18227;
  tri   n18228;
  tri   n18229;
  tri   n18230;
  tri   n18231;
  tri   n18232;
  tri   n18233;
  tri   n18234;
  tri   n18235;
  tri   n18236;
  tri   n18237;
  tri   n18238;
  tri   n18239;
  tri   n18240;
  tri   n18241;
  tri   n18242;
  tri   n18243;
  tri   n18244;
  tri   n18246;
  tri   n18247;
  tri   n18248;
  tri   n18249;
  tri   n18250;
  tri   n18251;
  tri   n18252;
  tri   n18253;
  tri   n18254;
  tri   n18255;
  tri   n18256;
  tri   n18257;
  tri   n18258;
  tri   n18259;
  tri   n18260;
  tri   n18261;
  tri   n18262;
  tri   n18263;
  tri   n18264;
  tri   n18265;
  tri   n18266;
  tri   n18267;
  tri   n18268;
  tri   n18269;
  tri   n18270;
  tri   n18271;
  tri   n18272;
  tri   n18273;
  tri   n18274;
  tri   n18275;
  tri   n18276;
  tri   n18277;
  tri   n18278;
  tri   n18279;
  tri   n18280;
  tri   n18281;
  tri   n18282;
  tri   n18283;
  tri   N74;
  tri   n18289;
  tri   n18290;
  tri   n18291;
  tri   n18292;
  tri   n18294;
  tri   n18295;
  tri   N71;
  tri   n18316;
  tri   n18317;
  tri   n18318;
  tri   n18319;
  tri   n18320;
  tri   n18321;
  tri   n18348;
  tri   n18349;
  tri   n18350;
  tri   n18351;
  tri   n18352;
  tri   n18353;
  tri   n18354;
  tri   n18355;
  tri   n18356;
  tri   n18357;
  tri   n18358;
  tri   n18359;
  tri   n18360;
  tri   n18361;
  tri   n18362;
  tri   n18363;
  tri   n18364;
  tri   n18365;
  tri   n18366;
  tri   n18367;
  tri   n18368;
  tri   n18369;
  tri   n18370;
  tri   n18371;
  tri   n18372;
  tri   n18373;
  tri   n18374;
  tri   n18375;
  tri   n18376;
  tri   n18377;
  tri   n18378;
  tri   n18379;
  tri   n18380;
  tri   n18381;
  tri   n18382;
  tri   n18383;
  tri   n18384;
  tri   n18385;
  tri   n18386;
  tri   n18387;
  tri   n18388;
  tri   n18389;
  tri   n18390;
  tri   n18391;
  tri   n18392;
  tri   n18393;
  tri   n17624;
  tri   n17623;
  tri   n17628;
  tri   n17626;
  tri   n17625;
  tri   n17630;
  tri   n17629;
  tri   n17627;
  tri   n17634;
  tri   n17633;
  tri   n17631;
  tri   n17643;
  tri   n17636;
  tri   n17635;
  tri   n17640;
  tri   n17638;
  tri   n17637;
  tri   n17642;
  tri   n17641;
  tri   n17639;
  tri   n17644;
  tri   n17646;
  tri   n17645;
  tri   n17650;
  tri   n17648;
  tri   n17647;
  tri   n17652;
  tri   n17651;
  tri   n17649;
  tri   n17662;
  tri   n17654;
  tri   n17653;
  tri   n17658;
  tri   n17656;
  tri   n17655;
  tri   n17660;
  tri   n17659;
  tri   n17657;
  tri   n17664;
  tri   n17663;
  tri   n17661;
  tri   n17673;
  tri   n17666;
  tri   n17665;
  tri   n17670;
  tri   n17668;
  tri   n17667;
  tri   n17672;
  tri   n17671;
  tri   n17669;
  tri   n17674;
  tri   n17676;
  tri   n17675;
  tri   n17680;
  tri   n17678;
  tri   n17677;
  tri   n17682;
  tri   n17681;
  tri   n17679;
  tri   n17692;
  tri   n17684;
  tri   n17683;
  tri   n17688;
  tri   n17686;
  tri   n17685;
  tri   n17690;
  tri   n17689;
  tri   n17687;
  tri   n17694;
  tri   n17693;
  tri   n17691;
  tri   n17703;
  tri   n17696;
  tri   n17695;
  tri   n17700;
  tri   n17698;
  tri   n17697;
  tri   n17702;
  tri   n17701;
  tri   n17699;
  tri   n17704;
  tri   n17706;
  tri   n17705;
  tri   n17710;
  tri   n17708;
  tri   n17707;
  tri   n17712;
  tri   n17711;
  tri   n17709;
  tri   n17722;
  tri   n17714;
  tri   n17713;
  tri   n17718;
  tri   n17716;
  tri   n17715;
  tri   n17720;
  tri   n17719;
  tri   n17717;
  tri   n17724;
  tri   n17723;
  tri   n17721;
  tri   n17733;
  tri   n17727;
  tri   n17726;
  tri   n17730;
  tri   n17729;
  tri   n17725;
  tri   n17732;
  tri   n17728;
  tri   n17731;
  tri   n17736;
  tri   n17735;
  tri   P1_N5180;
  tri   n17738;
  tri   n17737;
  tri   P2_N5102;
  tri   n18194;
  tri   n1503;
  tri   n18195;
  tri   n1504;
  tri   n18198;
  tri   n18199;
  tri   n18200;
  tri   n18201;
  tri   n18202;
  tri   n18203;
  tri   n18210;
  tri   n17346;
  tri   n17345;
  tri   n17350;
  tri   n17348;
  tri   n17347;
  tri   n17352;
  tri   n17351;
  tri   n17349;
  tri   n17362;
  tri   n17354;
  tri   n17353;
  tri   n17358;
  tri   n17356;
  tri   n17355;
  tri   n17360;
  tri   n17359;
  tri   n17357;
  tri   n17364;
  tri   n17363;
  tri   n17361;
  tri   n17373;
  tri   n17366;
  tri   n17365;
  tri   n17370;
  tri   n17368;
  tri   n17367;
  tri   n17372;
  tri   n17371;
  tri   n17369;
  tri   n17374;
  tri   n17376;
  tri   n17375;
  tri   n17380;
  tri   n17378;
  tri   n17377;
  tri   n17382;
  tri   n17381;
  tri   n17379;
  tri   n17392;
  tri   n17384;
  tri   n17383;
  tri   n17388;
  tri   n17386;
  tri   n17385;
  tri   n17390;
  tri   n17389;
  tri   n17387;
  tri   n17394;
  tri   n17393;
  tri   n17391;
  tri   n17403;
  tri   n17396;
  tri   n17395;
  tri   n17400;
  tri   n17398;
  tri   n17397;
  tri   n17402;
  tri   n17401;
  tri   n17399;
  tri   n17404;
  tri   n17406;
  tri   n17405;
  tri   n17410;
  tri   n17408;
  tri   n17407;
  tri   n17412;
  tri   n17411;
  tri   n17409;
  tri   n17422;
  tri   n17414;
  tri   n17413;
  tri   n17418;
  tri   n17416;
  tri   n17415;
  tri   n17420;
  tri   n17419;
  tri   n17417;
  tri   n17424;
  tri   n17423;
  tri   n17421;
  tri   n17433;
  tri   n17426;
  tri   n17425;
  tri   n17430;
  tri   n17428;
  tri   n17427;
  tri   n17432;
  tri   n17431;
  tri   n17429;
  tri   n17434;
  tri   n17436;
  tri   n17435;
  tri   n17440;
  tri   n17438;
  tri   n17437;
  tri   n17442;
  tri   n17441;
  tri   n17439;
  tri   n17452;
  tri   n17444;
  tri   n17443;
  tri   n17448;
  tri   n17446;
  tri   n17445;
  tri   n17450;
  tri   n17449;
  tri   n17447;
  tri   n17454;
  tri   n17453;
  tri   n17451;
  tri   n17463;
  tri   n17456;
  tri   n17455;
  tri   n17460;
  tri   n17458;
  tri   n17457;
  tri   n17462;
  tri   n17461;
  tri   n17459;
  tri   n17464;
  tri   n17466;
  tri   n17465;
  tri   n17470;
  tri   n17468;
  tri   n17467;
  tri   n17472;
  tri   n17471;
  tri   n17469;
  tri   n17482;
  tri   n17474;
  tri   n17473;
  tri   n17478;
  tri   n17476;
  tri   n17475;
  tri   n17480;
  tri   n17479;
  tri   n17477;
  tri   n17484;
  tri   n17483;
  tri   n17481;
  tri   n17493;
  tri   n17486;
  tri   n17485;
  tri   n17490;
  tri   n17488;
  tri   n17487;
  tri   n17492;
  tri   n17491;
  tri   n17489;
  tri   n17494;
  tri   n17496;
  tri   n17495;
  tri   n17500;
  tri   n17498;
  tri   n17497;
  tri   n17502;
  tri   n17501;
  tri   n17499;
  tri   n17512;
  tri   n17504;
  tri   n17503;
  tri   n17508;
  tri   n17506;
  tri   n17505;
  tri   n17510;
  tri   n17509;
  tri   n17507;
  tri   n17514;
  tri   n17513;
  tri   n17511;
  tri   n17523;
  tri   n17516;
  tri   n17515;
  tri   n17520;
  tri   n17518;
  tri   n17517;
  tri   n17522;
  tri   n17521;
  tri   n17519;
  tri   n17524;
  tri   n17526;
  tri   n17525;
  tri   n17530;
  tri   n17528;
  tri   n17527;
  tri   n17532;
  tri   n17531;
  tri   n17529;
  tri   n17542;
  tri   n17534;
  tri   n17533;
  tri   n17538;
  tri   n17536;
  tri   n17535;
  tri   n17540;
  tri   n17539;
  tri   n17537;
  tri   n17544;
  tri   n17543;
  tri   n17541;
  tri   n17553;
  tri   n17546;
  tri   n17545;
  tri   n17550;
  tri   n17548;
  tri   n17547;
  tri   n17552;
  tri   n17551;
  tri   n17549;
  tri   n17554;
  tri   n17556;
  tri   n17555;
  tri   n17560;
  tri   n17558;
  tri   n17557;
  tri   n17562;
  tri   n17561;
  tri   n17559;
  tri   n17572;
  tri   n17564;
  tri   n17563;
  tri   n17568;
  tri   n17566;
  tri   n17565;
  tri   n17570;
  tri   n17569;
  tri   n17567;
  tri   n17574;
  tri   n17573;
  tri   n17571;
  tri   n17583;
  tri   n17576;
  tri   n17575;
  tri   n17580;
  tri   n17578;
  tri   n17577;
  tri   n17582;
  tri   n17581;
  tri   n17579;
  tri   n17584;
  tri   n17586;
  tri   n17585;
  tri   n17590;
  tri   n17588;
  tri   n17587;
  tri   n17592;
  tri   n17591;
  tri   n17589;
  tri   n17602;
  tri   n17594;
  tri   n17593;
  tri   n17598;
  tri   n17596;
  tri   n17595;
  tri   n17600;
  tri   n17599;
  tri   n17597;
  tri   n17604;
  tri   n17603;
  tri   n17601;
  tri   n17613;
  tri   n17606;
  tri   n17605;
  tri   n17610;
  tri   n17608;
  tri   n17607;
  tri   n17612;
  tri   n17611;
  tri   n17609;
  tri   n17614;
  tri   n17616;
  tri   n17615;
  tri   n17620;
  tri   n17618;
  tri   n17617;
  tri   n17622;
  tri   n17621;
  tri   n17619;
  tri   n17632;
  tri   n17065;
  tri   n17064;
  tri   n17069;
  tri   n17068;
  tri   n17066;
  tri   n17071;
  tri   n17072;
  tri   n17070;
  tri   n17074;
  tri   n17076;
  tri   n17075;
  tri   n17078;
  tri   n17079;
  tri   n17077;
  tri   n17089;
  tri   n17081;
  tri   n17080;
  tri   n17085;
  tri   n17083;
  tri   n17082;
  tri   n17087;
  tri   n17086;
  tri   n17084;
  tri   n17091;
  tri   n17090;
  tri   n17088;
  tri   n17103;
  tri   n17093;
  tri   n17092;
  tri   n17097;
  tri   n17095;
  tri   n17094;
  tri   n17099;
  tri   n17098;
  tri   n17096;
  tri   n17101;
  tri   n17102;
  tri   n17100;
  tri   n17104;
  tri   n17106;
  tri   n17105;
  tri   n17110;
  tri   n17108;
  tri   n17107;
  tri   n17112;
  tri   n17111;
  tri   n17109;
  tri   n17122;
  tri   n17114;
  tri   n17113;
  tri   n17118;
  tri   n17116;
  tri   n17115;
  tri   n17120;
  tri   n17119;
  tri   n17117;
  tri   n17124;
  tri   n17123;
  tri   n17121;
  tri   n17133;
  tri   n17126;
  tri   n17125;
  tri   n17130;
  tri   n17128;
  tri   n17127;
  tri   n17132;
  tri   n17131;
  tri   n17129;
  tri   n17134;
  tri   n17136;
  tri   n17135;
  tri   n17140;
  tri   n17138;
  tri   n17137;
  tri   n17142;
  tri   n17141;
  tri   n17139;
  tri   n17152;
  tri   n17144;
  tri   n17143;
  tri   n17148;
  tri   n17146;
  tri   n17145;
  tri   n17150;
  tri   n17149;
  tri   n17147;
  tri   n17154;
  tri   n17153;
  tri   n17151;
  tri   n17163;
  tri   n17156;
  tri   n17155;
  tri   n17160;
  tri   n17158;
  tri   n17157;
  tri   n17162;
  tri   n17161;
  tri   n17159;
  tri   n17164;
  tri   n17166;
  tri   n17165;
  tri   n17170;
  tri   n17168;
  tri   n17167;
  tri   n17172;
  tri   n17171;
  tri   n17169;
  tri   n17182;
  tri   n17174;
  tri   n17173;
  tri   n17178;
  tri   n17176;
  tri   n17175;
  tri   n17180;
  tri   n17179;
  tri   n17177;
  tri   n17184;
  tri   n17183;
  tri   n17181;
  tri   n17193;
  tri   n17186;
  tri   n17185;
  tri   n17190;
  tri   n17188;
  tri   n17187;
  tri   n17192;
  tri   n17191;
  tri   n17189;
  tri   n17194;
  tri   n17196;
  tri   n17195;
  tri   n17200;
  tri   n17198;
  tri   n17197;
  tri   n17202;
  tri   n17201;
  tri   n17199;
  tri   n17212;
  tri   n17204;
  tri   n17203;
  tri   n17208;
  tri   n17206;
  tri   n17205;
  tri   n17210;
  tri   n17209;
  tri   n17207;
  tri   n17214;
  tri   n17213;
  tri   n17211;
  tri   n17223;
  tri   n17216;
  tri   n17215;
  tri   n17220;
  tri   n17218;
  tri   n17217;
  tri   n17222;
  tri   n17221;
  tri   n17219;
  tri   n17224;
  tri   n17226;
  tri   n17225;
  tri   n17230;
  tri   n17228;
  tri   n17227;
  tri   n17232;
  tri   n17231;
  tri   n17229;
  tri   n17242;
  tri   n17234;
  tri   n17233;
  tri   n17238;
  tri   n17236;
  tri   n17235;
  tri   n17240;
  tri   n17239;
  tri   n17237;
  tri   n17244;
  tri   n17243;
  tri   n17241;
  tri   n17253;
  tri   n17246;
  tri   n17245;
  tri   n17250;
  tri   n17248;
  tri   n17247;
  tri   n17252;
  tri   n17251;
  tri   n17249;
  tri   n17254;
  tri   n17256;
  tri   n17255;
  tri   n17260;
  tri   n17258;
  tri   n17257;
  tri   n17262;
  tri   n17261;
  tri   n17259;
  tri   n17272;
  tri   n17264;
  tri   n17263;
  tri   n17268;
  tri   n17266;
  tri   n17265;
  tri   n17270;
  tri   n17269;
  tri   n17267;
  tri   n17274;
  tri   n17273;
  tri   n17271;
  tri   n17283;
  tri   n17276;
  tri   n17275;
  tri   n17280;
  tri   n17278;
  tri   n17277;
  tri   n17282;
  tri   n17281;
  tri   n17279;
  tri   n17284;
  tri   n17286;
  tri   n17285;
  tri   n17290;
  tri   n17288;
  tri   n17287;
  tri   n17292;
  tri   n17291;
  tri   n17289;
  tri   n17302;
  tri   n17294;
  tri   n17293;
  tri   n17298;
  tri   n17296;
  tri   n17295;
  tri   n17300;
  tri   n17299;
  tri   n17297;
  tri   n17304;
  tri   n17303;
  tri   n17301;
  tri   n17313;
  tri   n17306;
  tri   n17305;
  tri   n17310;
  tri   n17308;
  tri   n17307;
  tri   n17312;
  tri   n17311;
  tri   n17309;
  tri   n17314;
  tri   n17316;
  tri   n17315;
  tri   n17320;
  tri   n17318;
  tri   n17317;
  tri   n17322;
  tri   n17321;
  tri   n17319;
  tri   n17332;
  tri   n17324;
  tri   n17323;
  tri   n17328;
  tri   n17326;
  tri   n17325;
  tri   n17330;
  tri   n17329;
  tri   n17327;
  tri   n17334;
  tri   n17333;
  tri   n17331;
  tri   n17343;
  tri   n17336;
  tri   n17335;
  tri   n17340;
  tri   n17338;
  tri   n17337;
  tri   n17342;
  tri   n17341;
  tri   n17339;
  tri   n17344;
  tri   n16786;
  tri   n16784;
  tri   n16799;
  tri   n16789;
  tri   n16788;
  tri   n16793;
  tri   n16791;
  tri   n16790;
  tri   n16795;
  tri   n16794;
  tri   n16792;
  tri   n16798;
  tri   n16797;
  tri   n16796;
  tri   n16800;
  tri   n16802;
  tri   n16801;
  tri   n16806;
  tri   n16804;
  tri   n16803;
  tri   n16808;
  tri   n16807;
  tri   n16805;
  tri   n16818;
  tri   n16810;
  tri   n16809;
  tri   n16814;
  tri   n16812;
  tri   n16811;
  tri   n16816;
  tri   n16815;
  tri   n16813;
  tri   n16820;
  tri   n16819;
  tri   n16817;
  tri   n16832;
  tri   n16822;
  tri   n16821;
  tri   n16826;
  tri   n16824;
  tri   n16823;
  tri   n16828;
  tri   n16827;
  tri   n16825;
  tri   n16831;
  tri   n16830;
  tri   n16829;
  tri   n16833;
  tri   n16835;
  tri   n16834;
  tri   n16838;
  tri   n16837;
  tri   n16836;
  tri   n16839;
  tri   n16841;
  tri   n16840;
  tri   n16844;
  tri   n16843;
  tri   n16842;
  tri   n16845;
  tri   n16847;
  tri   n16846;
  tri   n16850;
  tri   n16849;
  tri   n16848;
  tri   n16851;
  tri   n16853;
  tri   n16852;
  tri   n16856;
  tri   n16855;
  tri   n16854;
  tri   n16857;
  tri   n16859;
  tri   n16858;
  tri   n16862;
  tri   n16861;
  tri   n16860;
  tri   n16863;
  tri   n16865;
  tri   n16864;
  tri   n16868;
  tri   n16867;
  tri   n16866;
  tri   n16869;
  tri   n16871;
  tri   n16870;
  tri   n16874;
  tri   n16873;
  tri   n16872;
  tri   n16875;
  tri   n16877;
  tri   n16876;
  tri   n16880;
  tri   n16879;
  tri   n16878;
  tri   n16881;
  tri   n16883;
  tri   n16882;
  tri   n16886;
  tri   n16885;
  tri   n16884;
  tri   n16887;
  tri   n16889;
  tri   n16888;
  tri   n16892;
  tri   n16891;
  tri   n16890;
  tri   n16893;
  tri   n16895;
  tri   n16894;
  tri   n16898;
  tri   n16897;
  tri   n16896;
  tri   n16899;
  tri   n16901;
  tri   n16900;
  tri   n16904;
  tri   n16903;
  tri   n16902;
  tri   n16905;
  tri   n16907;
  tri   n16906;
  tri   n16910;
  tri   n16909;
  tri   n16908;
  tri   n16911;
  tri   n16913;
  tri   n16912;
  tri   n16916;
  tri   n16915;
  tri   n16914;
  tri   n16917;
  tri   n16919;
  tri   n16918;
  tri   n16922;
  tri   n16921;
  tri   n16920;
  tri   n16923;
  tri   n16925;
  tri   n16924;
  tri   n16928;
  tri   n16927;
  tri   n16926;
  tri   n16929;
  tri   n16931;
  tri   n16930;
  tri   n16934;
  tri   n16933;
  tri   n16932;
  tri   n16935;
  tri   n16937;
  tri   n16936;
  tri   n16940;
  tri   n16939;
  tri   n16938;
  tri   n16941;
  tri   n16943;
  tri   n16942;
  tri   n16946;
  tri   n16945;
  tri   n16944;
  tri   n16947;
  tri   n16949;
  tri   n16948;
  tri   n16952;
  tri   n16951;
  tri   n16950;
  tri   n16953;
  tri   n16955;
  tri   n16954;
  tri   n16958;
  tri   n16957;
  tri   n16956;
  tri   n16959;
  tri   n16961;
  tri   n16960;
  tri   n16964;
  tri   n16963;
  tri   n16962;
  tri   n16965;
  tri   n16967;
  tri   n16966;
  tri   n16970;
  tri   n16969;
  tri   n16968;
  tri   n16971;
  tri   n16973;
  tri   n16972;
  tri   n16976;
  tri   n16975;
  tri   n16974;
  tri   n16977;
  tri   n16979;
  tri   n16978;
  tri   n16982;
  tri   n16981;
  tri   n16980;
  tri   n16983;
  tri   n16985;
  tri   n16984;
  tri   n16988;
  tri   n16987;
  tri   n16986;
  tri   n16989;
  tri   n16991;
  tri   n16990;
  tri   n16994;
  tri   n16993;
  tri   n16992;
  tri   n16995;
  tri   n16997;
  tri   n16996;
  tri   n17000;
  tri   n16999;
  tri   n16998;
  tri   n17001;
  tri   n17003;
  tri   n17002;
  tri   n17006;
  tri   n17005;
  tri   n17004;
  tri   n17007;
  tri   n17009;
  tri   n17008;
  tri   n17012;
  tri   n17011;
  tri   n17010;
  tri   n17013;
  tri   n17015;
  tri   n17014;
  tri   n17017;
  tri   n17018;
  tri   n17016;
  tri   n17029;
  tri   n17021;
  tri   n17020;
  tri   n17025;
  tri   n17023;
  tri   n17022;
  tri   n17027;
  tri   n17026;
  tri   n17024;
  tri   n17031;
  tri   n17030;
  tri   n17028;
  tri   n17043;
  tri   n17033;
  tri   n17032;
  tri   n17037;
  tri   n17035;
  tri   n17034;
  tri   n17039;
  tri   n17038;
  tri   n17036;
  tri   n17041;
  tri   n17042;
  tri   n17040;
  tri   n17044;
  tri   n17046;
  tri   n17045;
  tri   n17048;
  tri   n17049;
  tri   n17047;
  tri   n17059;
  tri   n17051;
  tri   n17050;
  tri   n17055;
  tri   n17053;
  tri   n17052;
  tri   n17057;
  tri   n17056;
  tri   n17054;
  tri   n17061;
  tri   n17060;
  tri   n17058;
  tri   n17073;
  tri   n17063;
  tri   n17062;
  tri   n17067;
  tri   n16507;
  tri   n16506;
  tri   n16511;
  tri   n16510;
  tri   n16508;
  tri   n16521;
  tri   n16513;
  tri   n16512;
  tri   n16517;
  tri   n16515;
  tri   n16514;
  tri   n16519;
  tri   n16518;
  tri   n16516;
  tri   n16523;
  tri   n16522;
  tri   n16520;
  tri   n16535;
  tri   n16525;
  tri   n16524;
  tri   n16529;
  tri   n16527;
  tri   n16526;
  tri   n16531;
  tri   n16530;
  tri   n16528;
  tri   n16534;
  tri   n16533;
  tri   n16532;
  tri   n16536;
  tri   n16538;
  tri   n16537;
  tri   n16542;
  tri   n16540;
  tri   n16539;
  tri   n16544;
  tri   n16543;
  tri   n16541;
  tri   n16554;
  tri   n16546;
  tri   n16545;
  tri   n16550;
  tri   n16548;
  tri   n16547;
  tri   n16552;
  tri   n16551;
  tri   n16549;
  tri   n16556;
  tri   n16555;
  tri   n16553;
  tri   n16568;
  tri   n16558;
  tri   n16557;
  tri   n16562;
  tri   n16560;
  tri   n16559;
  tri   n16564;
  tri   n16563;
  tri   n16561;
  tri   n16567;
  tri   n16566;
  tri   n16565;
  tri   n16569;
  tri   n16571;
  tri   n16570;
  tri   n16575;
  tri   n16573;
  tri   n16572;
  tri   n16577;
  tri   n16576;
  tri   n16574;
  tri   n16587;
  tri   n16579;
  tri   n16578;
  tri   n16583;
  tri   n16581;
  tri   n16580;
  tri   n16585;
  tri   n16584;
  tri   n16582;
  tri   n16589;
  tri   n16588;
  tri   n16586;
  tri   n16601;
  tri   n16591;
  tri   n16590;
  tri   n16595;
  tri   n16593;
  tri   n16592;
  tri   n16597;
  tri   n16596;
  tri   n16594;
  tri   n16600;
  tri   n16599;
  tri   n16598;
  tri   n16602;
  tri   n16604;
  tri   n16603;
  tri   n16608;
  tri   n16606;
  tri   n16605;
  tri   n16610;
  tri   n16609;
  tri   n16607;
  tri   n16620;
  tri   n16612;
  tri   n16611;
  tri   n16616;
  tri   n16614;
  tri   n16613;
  tri   n16618;
  tri   n16617;
  tri   n16615;
  tri   n16622;
  tri   n16621;
  tri   n16619;
  tri   n16634;
  tri   n16624;
  tri   n16623;
  tri   n16628;
  tri   n16626;
  tri   n16625;
  tri   n16630;
  tri   n16629;
  tri   n16627;
  tri   n16633;
  tri   n16632;
  tri   n16631;
  tri   n16635;
  tri   n16637;
  tri   n16636;
  tri   n16641;
  tri   n16639;
  tri   n16638;
  tri   n16643;
  tri   n16642;
  tri   n16640;
  tri   n16653;
  tri   n16645;
  tri   n16644;
  tri   n16649;
  tri   n16647;
  tri   n16646;
  tri   n16651;
  tri   n16650;
  tri   n16648;
  tri   n16655;
  tri   n16654;
  tri   n16652;
  tri   n16667;
  tri   n16657;
  tri   n16656;
  tri   n16661;
  tri   n16659;
  tri   n16658;
  tri   n16663;
  tri   n16662;
  tri   n16660;
  tri   n16666;
  tri   n16665;
  tri   n16664;
  tri   n16668;
  tri   n16670;
  tri   n16669;
  tri   n16674;
  tri   n16672;
  tri   n16671;
  tri   n16676;
  tri   n16675;
  tri   n16673;
  tri   n16686;
  tri   n16678;
  tri   n16677;
  tri   n16682;
  tri   n16680;
  tri   n16679;
  tri   n16684;
  tri   n16683;
  tri   n16681;
  tri   n16688;
  tri   n16687;
  tri   n16685;
  tri   n16700;
  tri   n16690;
  tri   n16689;
  tri   n16694;
  tri   n16692;
  tri   n16691;
  tri   n16696;
  tri   n16695;
  tri   n16693;
  tri   n16699;
  tri   n16698;
  tri   n16697;
  tri   n16701;
  tri   n16703;
  tri   n16702;
  tri   n16707;
  tri   n16705;
  tri   n16704;
  tri   n16709;
  tri   n16708;
  tri   n16706;
  tri   n16719;
  tri   n16711;
  tri   n16710;
  tri   n16715;
  tri   n16713;
  tri   n16712;
  tri   n16717;
  tri   n16716;
  tri   n16714;
  tri   n16721;
  tri   n16720;
  tri   n16718;
  tri   n16733;
  tri   n16723;
  tri   n16722;
  tri   n16727;
  tri   n16725;
  tri   n16724;
  tri   n16729;
  tri   n16728;
  tri   n16726;
  tri   n16732;
  tri   n16731;
  tri   n16730;
  tri   n16734;
  tri   n16736;
  tri   n16735;
  tri   n16740;
  tri   n16738;
  tri   n16737;
  tri   n16742;
  tri   n16741;
  tri   n16739;
  tri   n16752;
  tri   n16744;
  tri   n16743;
  tri   n16748;
  tri   n16746;
  tri   n16745;
  tri   n16750;
  tri   n16749;
  tri   n16747;
  tri   n16754;
  tri   n16753;
  tri   n16751;
  tri   n16766;
  tri   n16756;
  tri   n16755;
  tri   n16760;
  tri   n16758;
  tri   n16757;
  tri   n16762;
  tri   n16761;
  tri   n16759;
  tri   n16765;
  tri   n16764;
  tri   n16763;
  tri   n16767;
  tri   n16769;
  tri   n16768;
  tri   n16773;
  tri   n16771;
  tri   n16770;
  tri   n16775;
  tri   n16774;
  tri   n16772;
  tri   n16785;
  tri   n16777;
  tri   n16776;
  tri   n16781;
  tri   n16779;
  tri   n16778;
  tri   n16783;
  tri   n16782;
  tri   n16780;
  tri   n16787;
  tri   n16228;
  tri   n16227;
  tri   n16232;
  tri   n16230;
  tri   n16229;
  tri   n16234;
  tri   n16233;
  tri   n16231;
  tri   n16237;
  tri   n16236;
  tri   n16235;
  tri   n16239;
  tri   n16241;
  tri   n16240;
  tri   n16245;
  tri   n16243;
  tri   n16242;
  tri   n16247;
  tri   n16246;
  tri   n16244;
  tri   n16257;
  tri   n16249;
  tri   n16248;
  tri   n16253;
  tri   n16251;
  tri   n16250;
  tri   n16255;
  tri   n16254;
  tri   n16252;
  tri   n16259;
  tri   n16258;
  tri   n16256;
  tri   n16271;
  tri   n16261;
  tri   n16260;
  tri   n16265;
  tri   n16263;
  tri   n16262;
  tri   n16267;
  tri   n16266;
  tri   n16264;
  tri   n16270;
  tri   n16269;
  tri   n16268;
  tri   n16272;
  tri   n16274;
  tri   n16273;
  tri   n16278;
  tri   n16276;
  tri   n16275;
  tri   n16280;
  tri   n16279;
  tri   n16277;
  tri   n16290;
  tri   n16282;
  tri   n16281;
  tri   n16286;
  tri   n16284;
  tri   n16283;
  tri   n16288;
  tri   n16287;
  tri   n16285;
  tri   n16292;
  tri   n16291;
  tri   n16289;
  tri   n16304;
  tri   n16294;
  tri   n16293;
  tri   n16298;
  tri   n16296;
  tri   n16295;
  tri   n16300;
  tri   n16299;
  tri   n16297;
  tri   n16303;
  tri   n16302;
  tri   n16301;
  tri   n16305;
  tri   n16307;
  tri   n16306;
  tri   n16311;
  tri   n16309;
  tri   n16308;
  tri   n16313;
  tri   n16312;
  tri   n16310;
  tri   n16323;
  tri   n16315;
  tri   n16314;
  tri   n16319;
  tri   n16317;
  tri   n16316;
  tri   n16321;
  tri   n16320;
  tri   n16318;
  tri   n16325;
  tri   n16324;
  tri   n16322;
  tri   n16337;
  tri   n16327;
  tri   n16326;
  tri   n16331;
  tri   n16329;
  tri   n16328;
  tri   n16333;
  tri   n16332;
  tri   n16330;
  tri   n16336;
  tri   n16335;
  tri   n16334;
  tri   n16338;
  tri   n16340;
  tri   n16339;
  tri   n16344;
  tri   n16342;
  tri   n16341;
  tri   n16346;
  tri   n16345;
  tri   n16343;
  tri   n16356;
  tri   n16348;
  tri   n16347;
  tri   n16352;
  tri   n16350;
  tri   n16349;
  tri   n16354;
  tri   n16353;
  tri   n16351;
  tri   n16358;
  tri   n16357;
  tri   n16355;
  tri   n16370;
  tri   n16360;
  tri   n16359;
  tri   n16364;
  tri   n16362;
  tri   n16361;
  tri   n16366;
  tri   n16365;
  tri   n16363;
  tri   n16369;
  tri   n16368;
  tri   n16367;
  tri   n16371;
  tri   n16373;
  tri   n16372;
  tri   n16377;
  tri   n16375;
  tri   n16374;
  tri   n16379;
  tri   n16378;
  tri   n16376;
  tri   n16389;
  tri   n16381;
  tri   n16380;
  tri   n16385;
  tri   n16383;
  tri   n16382;
  tri   n16387;
  tri   n16386;
  tri   n16384;
  tri   n16391;
  tri   n16390;
  tri   n16388;
  tri   n16403;
  tri   n16393;
  tri   n16392;
  tri   n16397;
  tri   n16395;
  tri   n16394;
  tri   n16399;
  tri   n16398;
  tri   n16396;
  tri   n16402;
  tri   n16401;
  tri   n16400;
  tri   n16404;
  tri   n16406;
  tri   n16405;
  tri   n16410;
  tri   n16408;
  tri   n16407;
  tri   n16412;
  tri   n16411;
  tri   n16409;
  tri   n16422;
  tri   n16414;
  tri   n16413;
  tri   n16418;
  tri   n16416;
  tri   n16415;
  tri   n16420;
  tri   n16419;
  tri   n16417;
  tri   n16424;
  tri   n16423;
  tri   n16421;
  tri   n16436;
  tri   n16426;
  tri   n16425;
  tri   n16430;
  tri   n16428;
  tri   n16427;
  tri   n16432;
  tri   n16431;
  tri   n16429;
  tri   n16435;
  tri   n16434;
  tri   n16433;
  tri   n16437;
  tri   n16439;
  tri   n16438;
  tri   n16443;
  tri   n16441;
  tri   n16440;
  tri   n16445;
  tri   n16444;
  tri   n16442;
  tri   n16455;
  tri   n16447;
  tri   n16446;
  tri   n16451;
  tri   n16449;
  tri   n16448;
  tri   n16453;
  tri   n16452;
  tri   n16450;
  tri   n16457;
  tri   n16456;
  tri   n16454;
  tri   n16469;
  tri   n16459;
  tri   n16458;
  tri   n16463;
  tri   n16461;
  tri   n16460;
  tri   n16465;
  tri   n16464;
  tri   n16462;
  tri   n16468;
  tri   n16467;
  tri   n16466;
  tri   n16470;
  tri   n16472;
  tri   n16471;
  tri   n16476;
  tri   n16474;
  tri   n16473;
  tri   n16478;
  tri   n16477;
  tri   n16475;
  tri   n16488;
  tri   n16480;
  tri   n16479;
  tri   n16484;
  tri   n16482;
  tri   n16481;
  tri   n16486;
  tri   n16485;
  tri   n16483;
  tri   n16490;
  tri   n16489;
  tri   n16487;
  tri   n16502;
  tri   n16492;
  tri   n16491;
  tri   n16496;
  tri   n16494;
  tri   n16493;
  tri   n16498;
  tri   n16497;
  tri   n16495;
  tri   n16501;
  tri   n16500;
  tri   n16499;
  tri   n16503;
  tri   n16505;
  tri   n16504;
  tri   n16509;
  tri   n15949;
  tri   n15947;
  tri   n15960;
  tri   n15952;
  tri   n15951;
  tri   n15956;
  tri   n15954;
  tri   n15953;
  tri   n15958;
  tri   n15957;
  tri   n15955;
  tri   n15962;
  tri   n15961;
  tri   n15959;
  tri   n15974;
  tri   n15964;
  tri   n15963;
  tri   n15968;
  tri   n15966;
  tri   n15965;
  tri   n15970;
  tri   n15969;
  tri   n15967;
  tri   n15973;
  tri   n15972;
  tri   n15971;
  tri   n15975;
  tri   n15977;
  tri   n15976;
  tri   n15981;
  tri   n15979;
  tri   n15978;
  tri   n15983;
  tri   n15982;
  tri   n15980;
  tri   n15993;
  tri   n15985;
  tri   n15984;
  tri   n15989;
  tri   n15987;
  tri   n15986;
  tri   n15991;
  tri   n15990;
  tri   n15988;
  tri   n15995;
  tri   n15994;
  tri   n15992;
  tri   n16007;
  tri   n15997;
  tri   n15996;
  tri   n16001;
  tri   n15999;
  tri   n15998;
  tri   n16003;
  tri   n16002;
  tri   n16000;
  tri   n16006;
  tri   n16005;
  tri   n16004;
  tri   n16008;
  tri   n16010;
  tri   n16009;
  tri   n16014;
  tri   n16012;
  tri   n16011;
  tri   n16016;
  tri   n16015;
  tri   n16013;
  tri   n16026;
  tri   n16018;
  tri   n16017;
  tri   n16022;
  tri   n16020;
  tri   n16019;
  tri   n16024;
  tri   n16023;
  tri   n16021;
  tri   n16028;
  tri   n16027;
  tri   n16025;
  tri   n16040;
  tri   n16030;
  tri   n16029;
  tri   n16034;
  tri   n16032;
  tri   n16031;
  tri   n16036;
  tri   n16035;
  tri   n16033;
  tri   n16039;
  tri   n16038;
  tri   n16037;
  tri   n16041;
  tri   n16043;
  tri   n16042;
  tri   n16047;
  tri   n16045;
  tri   n16044;
  tri   n16049;
  tri   n16048;
  tri   n16046;
  tri   n16059;
  tri   n16051;
  tri   n16050;
  tri   n16055;
  tri   n16053;
  tri   n16052;
  tri   n16057;
  tri   n16056;
  tri   n16054;
  tri   n16061;
  tri   n16060;
  tri   n16058;
  tri   n16073;
  tri   n16063;
  tri   n16062;
  tri   n16067;
  tri   n16065;
  tri   n16064;
  tri   n16069;
  tri   n16068;
  tri   n16066;
  tri   n16072;
  tri   n16071;
  tri   n16070;
  tri   n16074;
  tri   n16076;
  tri   n16075;
  tri   n16080;
  tri   n16078;
  tri   n16077;
  tri   n16082;
  tri   n16081;
  tri   n16079;
  tri   n16092;
  tri   n16084;
  tri   n16083;
  tri   n16088;
  tri   n16086;
  tri   n16085;
  tri   n16090;
  tri   n16089;
  tri   n16087;
  tri   n16094;
  tri   n16093;
  tri   n16091;
  tri   n16106;
  tri   n16096;
  tri   n16095;
  tri   n16100;
  tri   n16098;
  tri   n16097;
  tri   n16102;
  tri   n16101;
  tri   n16099;
  tri   n16105;
  tri   n16104;
  tri   n16103;
  tri   n16107;
  tri   n16109;
  tri   n16108;
  tri   n16113;
  tri   n16111;
  tri   n16110;
  tri   n16115;
  tri   n16114;
  tri   n16112;
  tri   n16125;
  tri   n16117;
  tri   n16116;
  tri   n16121;
  tri   n16119;
  tri   n16118;
  tri   n16123;
  tri   n16122;
  tri   n16120;
  tri   n16127;
  tri   n16126;
  tri   n16124;
  tri   n16139;
  tri   n16129;
  tri   n16128;
  tri   n16133;
  tri   n16131;
  tri   n16130;
  tri   n16135;
  tri   n16134;
  tri   n16132;
  tri   n16138;
  tri   n16137;
  tri   n16136;
  tri   n16140;
  tri   n16142;
  tri   n16141;
  tri   n16146;
  tri   n16144;
  tri   n16143;
  tri   n16148;
  tri   n16147;
  tri   n16145;
  tri   n16158;
  tri   n16150;
  tri   n16149;
  tri   n16154;
  tri   n16152;
  tri   n16151;
  tri   n16156;
  tri   n16155;
  tri   n16153;
  tri   n16160;
  tri   n16159;
  tri   n16157;
  tri   n16172;
  tri   n16162;
  tri   n16161;
  tri   n16166;
  tri   n16164;
  tri   n16163;
  tri   n16168;
  tri   n16167;
  tri   n16165;
  tri   n16171;
  tri   n16170;
  tri   n16169;
  tri   n16173;
  tri   n16175;
  tri   n16174;
  tri   n16179;
  tri   n16177;
  tri   n16176;
  tri   n16181;
  tri   n16180;
  tri   n16178;
  tri   n16191;
  tri   n16183;
  tri   n16182;
  tri   n16187;
  tri   n16185;
  tri   n16184;
  tri   n16189;
  tri   n16188;
  tri   n16186;
  tri   n16193;
  tri   n16192;
  tri   n16190;
  tri   n16205;
  tri   n16195;
  tri   n16194;
  tri   n16199;
  tri   n16197;
  tri   n16196;
  tri   n16201;
  tri   n16200;
  tri   n16198;
  tri   n16204;
  tri   n16203;
  tri   n16202;
  tri   n16206;
  tri   n16208;
  tri   n16207;
  tri   n16212;
  tri   n16210;
  tri   n16209;
  tri   n16214;
  tri   n16213;
  tri   n16211;
  tri   n16224;
  tri   n16216;
  tri   n16215;
  tri   n16220;
  tri   n16218;
  tri   n16217;
  tri   n16222;
  tri   n16221;
  tri   n16219;
  tri   n16226;
  tri   n16225;
  tri   n16223;
  tri   n16238;
  tri   n15670;
  tri   n15668;
  tri   n15681;
  tri   n15673;
  tri   n15672;
  tri   n15677;
  tri   n15675;
  tri   n15674;
  tri   n15679;
  tri   n15678;
  tri   n15676;
  tri   n15683;
  tri   n15682;
  tri   n15680;
  tri   n15698;
  tri   n15685;
  tri   n15684;
  tri   n15689;
  tri   n15687;
  tri   n15686;
  tri   n15691;
  tri   n15690;
  tri   n15688;
  tri   n15695;
  tri   n15693;
  tri   n15692;
  tri   n15697;
  tri   n15696;
  tri   n15694;
  tri   n15699;
  tri   n15701;
  tri   n15700;
  tri   n15705;
  tri   n15703;
  tri   n15702;
  tri   n15707;
  tri   n15706;
  tri   n15704;
  tri   n15717;
  tri   n15709;
  tri   n15708;
  tri   n15713;
  tri   n15711;
  tri   n15710;
  tri   n15715;
  tri   n15714;
  tri   n15712;
  tri   n15719;
  tri   n15718;
  tri   n15716;
  tri   n15734;
  tri   n15721;
  tri   n15720;
  tri   n15725;
  tri   n15723;
  tri   n15722;
  tri   n15727;
  tri   n15726;
  tri   n15724;
  tri   n15731;
  tri   n15729;
  tri   n15728;
  tri   n15733;
  tri   n15732;
  tri   n15730;
  tri   n15735;
  tri   n15737;
  tri   n15736;
  tri   n15741;
  tri   n15739;
  tri   n15738;
  tri   n15743;
  tri   n15742;
  tri   n15740;
  tri   n15753;
  tri   n15745;
  tri   n15744;
  tri   n15749;
  tri   n15747;
  tri   n15746;
  tri   n15751;
  tri   n15750;
  tri   n15748;
  tri   n15755;
  tri   n15754;
  tri   n15752;
  tri   n15770;
  tri   n15757;
  tri   n15756;
  tri   n15761;
  tri   n15759;
  tri   n15758;
  tri   n15763;
  tri   n15762;
  tri   n15760;
  tri   n15767;
  tri   n15765;
  tri   n15764;
  tri   n15769;
  tri   n15768;
  tri   n15766;
  tri   n15771;
  tri   n15773;
  tri   n15772;
  tri   n15777;
  tri   n15775;
  tri   n15774;
  tri   n15779;
  tri   n15778;
  tri   n15776;
  tri   n15789;
  tri   n15781;
  tri   n15780;
  tri   n15785;
  tri   n15783;
  tri   n15782;
  tri   n15787;
  tri   n15786;
  tri   n15784;
  tri   n15791;
  tri   n15790;
  tri   n15788;
  tri   n15806;
  tri   n15793;
  tri   n15792;
  tri   n15797;
  tri   n15795;
  tri   n15794;
  tri   n15799;
  tri   n15798;
  tri   n15796;
  tri   n15803;
  tri   n15801;
  tri   n15800;
  tri   n15805;
  tri   n15804;
  tri   n15802;
  tri   n15807;
  tri   n15809;
  tri   n15808;
  tri   n15813;
  tri   n15811;
  tri   n15810;
  tri   n15815;
  tri   n15814;
  tri   n15812;
  tri   n15825;
  tri   n15817;
  tri   n15816;
  tri   n15821;
  tri   n15819;
  tri   n15818;
  tri   n15823;
  tri   n15822;
  tri   n15820;
  tri   n15827;
  tri   n15826;
  tri   n15824;
  tri   n15842;
  tri   n15829;
  tri   n15828;
  tri   n15833;
  tri   n15831;
  tri   n15830;
  tri   n15835;
  tri   n15834;
  tri   n15832;
  tri   n15839;
  tri   n15837;
  tri   n15836;
  tri   n15841;
  tri   n15840;
  tri   n15838;
  tri   n15843;
  tri   n15845;
  tri   n15844;
  tri   n15849;
  tri   n15847;
  tri   n15846;
  tri   n15851;
  tri   n15850;
  tri   n15848;
  tri   n15861;
  tri   n15853;
  tri   n15852;
  tri   n15857;
  tri   n15855;
  tri   n15854;
  tri   n15859;
  tri   n15858;
  tri   n15856;
  tri   n15863;
  tri   n15862;
  tri   n15860;
  tri   n15875;
  tri   n15865;
  tri   n15864;
  tri   n15869;
  tri   n15867;
  tri   n15866;
  tri   n15871;
  tri   n15870;
  tri   n15868;
  tri   n15874;
  tri   n15873;
  tri   n15872;
  tri   n15876;
  tri   n15878;
  tri   n15877;
  tri   n15882;
  tri   n15880;
  tri   n15879;
  tri   n15884;
  tri   n15883;
  tri   n15881;
  tri   n15894;
  tri   n15886;
  tri   n15885;
  tri   n15890;
  tri   n15888;
  tri   n15887;
  tri   n15892;
  tri   n15891;
  tri   n15889;
  tri   n15896;
  tri   n15895;
  tri   n15893;
  tri   n15908;
  tri   n15898;
  tri   n15897;
  tri   n15902;
  tri   n15900;
  tri   n15899;
  tri   n15904;
  tri   n15903;
  tri   n15901;
  tri   n15907;
  tri   n15906;
  tri   n15905;
  tri   n15909;
  tri   n15911;
  tri   n15910;
  tri   n15915;
  tri   n15913;
  tri   n15912;
  tri   n15917;
  tri   n15916;
  tri   n15914;
  tri   n15927;
  tri   n15919;
  tri   n15918;
  tri   n15923;
  tri   n15921;
  tri   n15920;
  tri   n15925;
  tri   n15924;
  tri   n15922;
  tri   n15929;
  tri   n15928;
  tri   n15926;
  tri   n15941;
  tri   n15931;
  tri   n15930;
  tri   n15935;
  tri   n15933;
  tri   n15932;
  tri   n15937;
  tri   n15936;
  tri   n15934;
  tri   n15940;
  tri   n15939;
  tri   n15938;
  tri   n15942;
  tri   n15944;
  tri   n15943;
  tri   n15948;
  tri   n15946;
  tri   n15945;
  tri   n15950;
  tri   n15390;
  tri   n15388;
  tri   n15395;
  tri   n15394;
  tri   n15392;
  tri   n15410;
  tri   n15397;
  tri   n15396;
  tri   n15401;
  tri   n15399;
  tri   n15398;
  tri   n15403;
  tri   n15402;
  tri   n15400;
  tri   n15407;
  tri   n15405;
  tri   n15404;
  tri   n15409;
  tri   n15408;
  tri   n15406;
  tri   n15411;
  tri   n15413;
  tri   n15412;
  tri   n15417;
  tri   n15415;
  tri   n15414;
  tri   n15419;
  tri   n15418;
  tri   n15416;
  tri   n15429;
  tri   n15421;
  tri   n15420;
  tri   n15425;
  tri   n15423;
  tri   n15422;
  tri   n15427;
  tri   n15426;
  tri   n15424;
  tri   n15431;
  tri   n15430;
  tri   n15428;
  tri   n15446;
  tri   n15433;
  tri   n15432;
  tri   n15437;
  tri   n15435;
  tri   n15434;
  tri   n15439;
  tri   n15438;
  tri   n15436;
  tri   n15443;
  tri   n15441;
  tri   n15440;
  tri   n15445;
  tri   n15444;
  tri   n15442;
  tri   n15447;
  tri   n15449;
  tri   n15448;
  tri   n15453;
  tri   n15451;
  tri   n15450;
  tri   n15455;
  tri   n15454;
  tri   n15452;
  tri   n15465;
  tri   n15457;
  tri   n15456;
  tri   n15461;
  tri   n15459;
  tri   n15458;
  tri   n15463;
  tri   n15462;
  tri   n15460;
  tri   n15467;
  tri   n15466;
  tri   n15464;
  tri   n15482;
  tri   n15469;
  tri   n15468;
  tri   n15473;
  tri   n15471;
  tri   n15470;
  tri   n15475;
  tri   n15474;
  tri   n15472;
  tri   n15479;
  tri   n15477;
  tri   n15476;
  tri   n15481;
  tri   n15480;
  tri   n15478;
  tri   n15483;
  tri   n15485;
  tri   n15484;
  tri   n15489;
  tri   n15487;
  tri   n15486;
  tri   n15491;
  tri   n15490;
  tri   n15488;
  tri   n15501;
  tri   n15493;
  tri   n15492;
  tri   n15497;
  tri   n15495;
  tri   n15494;
  tri   n15499;
  tri   n15498;
  tri   n15496;
  tri   n15503;
  tri   n15502;
  tri   n15500;
  tri   n15518;
  tri   n15505;
  tri   n15504;
  tri   n15509;
  tri   n15507;
  tri   n15506;
  tri   n15511;
  tri   n15510;
  tri   n15508;
  tri   n15515;
  tri   n15513;
  tri   n15512;
  tri   n15517;
  tri   n15516;
  tri   n15514;
  tri   n15519;
  tri   n15521;
  tri   n15520;
  tri   n15525;
  tri   n15523;
  tri   n15522;
  tri   n15527;
  tri   n15526;
  tri   n15524;
  tri   n15537;
  tri   n15529;
  tri   n15528;
  tri   n15533;
  tri   n15531;
  tri   n15530;
  tri   n15535;
  tri   n15534;
  tri   n15532;
  tri   n15539;
  tri   n15538;
  tri   n15536;
  tri   n15554;
  tri   n15541;
  tri   n15540;
  tri   n15545;
  tri   n15543;
  tri   n15542;
  tri   n15547;
  tri   n15546;
  tri   n15544;
  tri   n15551;
  tri   n15549;
  tri   n15548;
  tri   n15553;
  tri   n15552;
  tri   n15550;
  tri   n15555;
  tri   n15557;
  tri   n15556;
  tri   n15561;
  tri   n15559;
  tri   n15558;
  tri   n15563;
  tri   n15562;
  tri   n15560;
  tri   n15573;
  tri   n15565;
  tri   n15564;
  tri   n15569;
  tri   n15567;
  tri   n15566;
  tri   n15571;
  tri   n15570;
  tri   n15568;
  tri   n15575;
  tri   n15574;
  tri   n15572;
  tri   n15590;
  tri   n15577;
  tri   n15576;
  tri   n15581;
  tri   n15579;
  tri   n15578;
  tri   n15583;
  tri   n15582;
  tri   n15580;
  tri   n15587;
  tri   n15585;
  tri   n15584;
  tri   n15589;
  tri   n15588;
  tri   n15586;
  tri   n15591;
  tri   n15593;
  tri   n15592;
  tri   n15597;
  tri   n15595;
  tri   n15594;
  tri   n15599;
  tri   n15598;
  tri   n15596;
  tri   n15609;
  tri   n15601;
  tri   n15600;
  tri   n15605;
  tri   n15603;
  tri   n15602;
  tri   n15607;
  tri   n15606;
  tri   n15604;
  tri   n15611;
  tri   n15610;
  tri   n15608;
  tri   n15626;
  tri   n15613;
  tri   n15612;
  tri   n15617;
  tri   n15615;
  tri   n15614;
  tri   n15619;
  tri   n15618;
  tri   n15616;
  tri   n15623;
  tri   n15621;
  tri   n15620;
  tri   n15625;
  tri   n15624;
  tri   n15622;
  tri   n15627;
  tri   n15629;
  tri   n15628;
  tri   n15633;
  tri   n15631;
  tri   n15630;
  tri   n15635;
  tri   n15634;
  tri   n15632;
  tri   n15645;
  tri   n15637;
  tri   n15636;
  tri   n15641;
  tri   n15639;
  tri   n15638;
  tri   n15643;
  tri   n15642;
  tri   n15640;
  tri   n15647;
  tri   n15646;
  tri   n15644;
  tri   n15662;
  tri   n15649;
  tri   n15648;
  tri   n15653;
  tri   n15651;
  tri   n15650;
  tri   n15655;
  tri   n15654;
  tri   n15652;
  tri   n15659;
  tri   n15657;
  tri   n15656;
  tri   n15661;
  tri   n15660;
  tri   n15658;
  tri   n15663;
  tri   n15665;
  tri   n15664;
  tri   n15669;
  tri   n15667;
  tri   n15666;
  tri   n15671;
  tri   n15111;
  tri   n15110;
  tri   n15115;
  tri   n15114;
  tri   n15112;
  tri   n15119;
  tri   n15117;
  tri   n15116;
  tri   n15121;
  tri   n15120;
  tri   n15118;
  tri   n15123;
  tri   n15125;
  tri   n15124;
  tri   n15129;
  tri   n15127;
  tri   n15126;
  tri   n15131;
  tri   n15130;
  tri   n15128;
  tri   n15141;
  tri   n15133;
  tri   n15132;
  tri   n15137;
  tri   n15135;
  tri   n15134;
  tri   n15139;
  tri   n15138;
  tri   n15136;
  tri   n15143;
  tri   n15142;
  tri   n15140;
  tri   n15158;
  tri   n15145;
  tri   n15144;
  tri   n15149;
  tri   n15147;
  tri   n15146;
  tri   n15151;
  tri   n15150;
  tri   n15148;
  tri   n15155;
  tri   n15153;
  tri   n15152;
  tri   n15157;
  tri   n15156;
  tri   n15154;
  tri   n15159;
  tri   n15161;
  tri   n15160;
  tri   n15165;
  tri   n15163;
  tri   n15162;
  tri   n15167;
  tri   n15166;
  tri   n15164;
  tri   n15177;
  tri   n15169;
  tri   n15168;
  tri   n15173;
  tri   n15171;
  tri   n15170;
  tri   n15175;
  tri   n15174;
  tri   n15172;
  tri   n15179;
  tri   n15178;
  tri   n15176;
  tri   n15194;
  tri   n15181;
  tri   n15180;
  tri   n15185;
  tri   n15183;
  tri   n15182;
  tri   n15187;
  tri   n15186;
  tri   n15184;
  tri   n15191;
  tri   n15189;
  tri   n15188;
  tri   n15193;
  tri   n15192;
  tri   n15190;
  tri   n15195;
  tri   n15197;
  tri   n15196;
  tri   n15201;
  tri   n15199;
  tri   n15198;
  tri   n15203;
  tri   n15202;
  tri   n15200;
  tri   n15213;
  tri   n15205;
  tri   n15204;
  tri   n15209;
  tri   n15207;
  tri   n15206;
  tri   n15211;
  tri   n15210;
  tri   n15208;
  tri   n15215;
  tri   n15214;
  tri   n15212;
  tri   n15230;
  tri   n15217;
  tri   n15216;
  tri   n15221;
  tri   n15219;
  tri   n15218;
  tri   n15223;
  tri   n15222;
  tri   n15220;
  tri   n15227;
  tri   n15225;
  tri   n15224;
  tri   n15229;
  tri   n15228;
  tri   n15226;
  tri   n15231;
  tri   n15233;
  tri   n15232;
  tri   n15237;
  tri   n15235;
  tri   n15234;
  tri   n15239;
  tri   n15238;
  tri   n15236;
  tri   n15249;
  tri   n15241;
  tri   n15240;
  tri   n15245;
  tri   n15243;
  tri   n15242;
  tri   n15247;
  tri   n15246;
  tri   n15244;
  tri   n15251;
  tri   n15250;
  tri   n15248;
  tri   n15266;
  tri   n15253;
  tri   n15252;
  tri   n15257;
  tri   n15255;
  tri   n15254;
  tri   n15259;
  tri   n15258;
  tri   n15256;
  tri   n15263;
  tri   n15261;
  tri   n15260;
  tri   n15265;
  tri   n15264;
  tri   n15262;
  tri   n15267;
  tri   n15269;
  tri   n15268;
  tri   n15273;
  tri   n15271;
  tri   n15270;
  tri   n15275;
  tri   n15274;
  tri   n15272;
  tri   n15285;
  tri   n15277;
  tri   n15276;
  tri   n15281;
  tri   n15279;
  tri   n15278;
  tri   n15283;
  tri   n15282;
  tri   n15280;
  tri   n15287;
  tri   n15286;
  tri   n15284;
  tri   n15302;
  tri   n15289;
  tri   n15288;
  tri   n15293;
  tri   n15291;
  tri   n15290;
  tri   n15295;
  tri   n15294;
  tri   n15292;
  tri   n15299;
  tri   n15297;
  tri   n15296;
  tri   n15301;
  tri   n15300;
  tri   n15298;
  tri   n15303;
  tri   n15305;
  tri   n15304;
  tri   n15309;
  tri   n15307;
  tri   n15306;
  tri   n15311;
  tri   n15310;
  tri   n15308;
  tri   n15321;
  tri   n15313;
  tri   n15312;
  tri   n15317;
  tri   n15315;
  tri   n15314;
  tri   n15319;
  tri   n15318;
  tri   n15316;
  tri   n15323;
  tri   n15322;
  tri   n15320;
  tri   n15338;
  tri   n15325;
  tri   n15324;
  tri   n15329;
  tri   n15327;
  tri   n15326;
  tri   n15331;
  tri   n15330;
  tri   n15328;
  tri   n15335;
  tri   n15333;
  tri   n15332;
  tri   n15337;
  tri   n15336;
  tri   n15334;
  tri   n15339;
  tri   n15341;
  tri   n15340;
  tri   n15345;
  tri   n15343;
  tri   n15342;
  tri   n15347;
  tri   n15346;
  tri   n15344;
  tri   n15357;
  tri   n15349;
  tri   n15348;
  tri   n15353;
  tri   n15351;
  tri   n15350;
  tri   n15355;
  tri   n15354;
  tri   n15352;
  tri   n15359;
  tri   n15358;
  tri   n15356;
  tri   n15374;
  tri   n15361;
  tri   n15360;
  tri   n15365;
  tri   n15363;
  tri   n15362;
  tri   n15367;
  tri   n15366;
  tri   n15364;
  tri   n15371;
  tri   n15369;
  tri   n15368;
  tri   n15373;
  tri   n15372;
  tri   n15370;
  tri   n15375;
  tri   n15377;
  tri   n15376;
  tri   n15381;
  tri   n15379;
  tri   n15378;
  tri   n15383;
  tri   n15382;
  tri   n15380;
  tri   n15393;
  tri   n15385;
  tri   n15384;
  tri   n15389;
  tri   n15387;
  tri   n15386;
  tri   n15391;
  tri   n14832;
  tri   n14830;
  tri   n14835;
  tri   n14837;
  tri   n14836;
  tri   n14841;
  tri   n14839;
  tri   n14838;
  tri   n14843;
  tri   n14842;
  tri   n14840;
  tri   n14853;
  tri   n14845;
  tri   n14844;
  tri   n14849;
  tri   n14847;
  tri   n14846;
  tri   n14851;
  tri   n14850;
  tri   n14848;
  tri   n14855;
  tri   n14854;
  tri   n14852;
  tri   n14870;
  tri   n14857;
  tri   n14856;
  tri   n14861;
  tri   n14859;
  tri   n14858;
  tri   n14863;
  tri   n14862;
  tri   n14860;
  tri   n14867;
  tri   n14865;
  tri   n14864;
  tri   n14869;
  tri   n14868;
  tri   n14866;
  tri   n14871;
  tri   n14873;
  tri   n14872;
  tri   n14877;
  tri   n14875;
  tri   n14874;
  tri   n14879;
  tri   n14878;
  tri   n14876;
  tri   n14889;
  tri   n14881;
  tri   n14880;
  tri   n14885;
  tri   n14883;
  tri   n14882;
  tri   n14887;
  tri   n14886;
  tri   n14884;
  tri   n14891;
  tri   n14890;
  tri   n14888;
  tri   n14906;
  tri   n14893;
  tri   n14892;
  tri   n14897;
  tri   n14895;
  tri   n14894;
  tri   n14899;
  tri   n14898;
  tri   n14896;
  tri   n14903;
  tri   n14901;
  tri   n14900;
  tri   n14905;
  tri   n14904;
  tri   n14902;
  tri   n14907;
  tri   n14909;
  tri   n14908;
  tri   n14913;
  tri   n14911;
  tri   n14910;
  tri   n14915;
  tri   n14914;
  tri   n14912;
  tri   n14925;
  tri   n14917;
  tri   n14916;
  tri   n14921;
  tri   n14919;
  tri   n14918;
  tri   n14923;
  tri   n14922;
  tri   n14920;
  tri   n14927;
  tri   n14926;
  tri   n14924;
  tri   n14942;
  tri   n14929;
  tri   n14928;
  tri   n14933;
  tri   n14931;
  tri   n14930;
  tri   n14935;
  tri   n14934;
  tri   n14932;
  tri   n14939;
  tri   n14937;
  tri   n14936;
  tri   n14941;
  tri   n14940;
  tri   n14938;
  tri   n14943;
  tri   n14945;
  tri   n14944;
  tri   n14949;
  tri   n14947;
  tri   n14946;
  tri   n14951;
  tri   n14950;
  tri   n14948;
  tri   n14961;
  tri   n14953;
  tri   n14952;
  tri   n14957;
  tri   n14955;
  tri   n14954;
  tri   n14959;
  tri   n14958;
  tri   n14956;
  tri   n14963;
  tri   n14962;
  tri   n14960;
  tri   n14978;
  tri   n14965;
  tri   n14964;
  tri   n14969;
  tri   n14967;
  tri   n14966;
  tri   n14971;
  tri   n14970;
  tri   n14968;
  tri   n14975;
  tri   n14973;
  tri   n14972;
  tri   n14977;
  tri   n14976;
  tri   n14974;
  tri   n14979;
  tri   n14981;
  tri   n14980;
  tri   n14985;
  tri   n14983;
  tri   n14982;
  tri   n14987;
  tri   n14986;
  tri   n14984;
  tri   n14997;
  tri   n14989;
  tri   n14988;
  tri   n14993;
  tri   n14991;
  tri   n14990;
  tri   n14995;
  tri   n14994;
  tri   n14992;
  tri   n14999;
  tri   n14998;
  tri   n14996;
  tri   n15014;
  tri   n15001;
  tri   n15000;
  tri   n15005;
  tri   n15003;
  tri   n15002;
  tri   n15007;
  tri   n15006;
  tri   n15004;
  tri   n15011;
  tri   n15009;
  tri   n15008;
  tri   n15013;
  tri   n15012;
  tri   n15010;
  tri   n15015;
  tri   n15017;
  tri   n15016;
  tri   n15021;
  tri   n15019;
  tri   n15018;
  tri   n15023;
  tri   n15022;
  tri   n15020;
  tri   n15033;
  tri   n15025;
  tri   n15024;
  tri   n15029;
  tri   n15027;
  tri   n15026;
  tri   n15031;
  tri   n15030;
  tri   n15028;
  tri   n15035;
  tri   n15034;
  tri   n15032;
  tri   n15050;
  tri   n15037;
  tri   n15036;
  tri   n15041;
  tri   n15039;
  tri   n15038;
  tri   n15043;
  tri   n15042;
  tri   n15040;
  tri   n15047;
  tri   n15045;
  tri   n15044;
  tri   n15049;
  tri   n15048;
  tri   n15046;
  tri   n15051;
  tri   n15053;
  tri   n15052;
  tri   n15057;
  tri   n15055;
  tri   n15054;
  tri   n15059;
  tri   n15058;
  tri   n15056;
  tri   n15069;
  tri   n15061;
  tri   n15060;
  tri   n15065;
  tri   n15063;
  tri   n15062;
  tri   n15067;
  tri   n15066;
  tri   n15064;
  tri   n15071;
  tri   n15070;
  tri   n15068;
  tri   n15086;
  tri   n15073;
  tri   n15072;
  tri   n15077;
  tri   n15075;
  tri   n15074;
  tri   n15079;
  tri   n15078;
  tri   n15076;
  tri   n15083;
  tri   n15081;
  tri   n15080;
  tri   n15085;
  tri   n15084;
  tri   n15082;
  tri   n15087;
  tri   n15089;
  tri   n15088;
  tri   n15093;
  tri   n15091;
  tri   n15090;
  tri   n15095;
  tri   n15094;
  tri   n15092;
  tri   n15105;
  tri   n15097;
  tri   n15096;
  tri   n15101;
  tri   n15099;
  tri   n15098;
  tri   n15103;
  tri   n15102;
  tri   n15100;
  tri   n15107;
  tri   n15106;
  tri   n15104;
  tri   n15122;
  tri   n15109;
  tri   n15108;
  tri   n15113;
  tri   n14752;
  tri   n14753;
  tri   P2_N933;
  tri   n14754;
  tri   n14755;
  tri   P2_N934;
  tri   n14756;
  tri   n14757;
  tri   n14759;
  tri   n14760;
  tri   n14758;
  tri   n14761;
  tri   n17019;
  tri   n14764;
  tri   n14762;
  tri   n14774;
  tri   n14766;
  tri   n14765;
  tri   n14770;
  tri   n14768;
  tri   n14767;
  tri   n14772;
  tri   n14771;
  tri   n14769;
  tri   n14776;
  tri   n14775;
  tri   n14773;
  tri   n14798;
  tri   n14778;
  tri   n14777;
  tri   n14782;
  tri   n14780;
  tri   n14779;
  tri   n14784;
  tri   n14783;
  tri   n14781;
  tri   n14794;
  tri   n14786;
  tri   n14785;
  tri   n14790;
  tri   n14788;
  tri   n14787;
  tri   n14792;
  tri   n14791;
  tri   n14789;
  tri   n14796;
  tri   n14795;
  tri   n14793;
  tri   n14799;
  tri   n14801;
  tri   n14800;
  tri   n14805;
  tri   n14803;
  tri   n14802;
  tri   n14807;
  tri   n14806;
  tri   n14804;
  tri   n14817;
  tri   n14809;
  tri   n14808;
  tri   n14813;
  tri   n14811;
  tri   n14810;
  tri   n14815;
  tri   n14814;
  tri   n14812;
  tri   n14819;
  tri   n14818;
  tri   n14816;
  tri   n14834;
  tri   n14821;
  tri   n14820;
  tri   n14825;
  tri   n14823;
  tri   n14822;
  tri   n14827;
  tri   n14826;
  tri   n14824;
  tri   n14831;
  tri   n14829;
  tri   n14828;
  tri   n14833;
  tri   n14744;
  tri   n14745;
  tri   n14746;
  tri   n14747;
  tri   P2_N930;
  tri   n14748;
  tri   n14749;
  tri   P2_N931;
  tri   n14750;
  tri   n14751;
  tri   P2_N932;
  tri   P2_N924;
  tri   n14736;
  tri   n14737;
  tri   n14738;
  tri   n14739;
  tri   P2_N926;
  tri   n14740;
  tri   n14741;
  tri   P2_N927;
  tri   n14742;
  tri   n14743;
  tri   P2_N920;
  tri   n14728;
  tri   n14729;
  tri   P2_N921;
  tri   n14730;
  tri   n14731;
  tri   P2_N922;
  tri   n14732;
  tri   n14733;
  tri   P2_N923;
  tri   n14734;
  tri   n14735;
  tri   n14718;
  tri   n14719;
  tri   P2_N916;
  tri   n14720;
  tri   n14721;
  tri   P2_N917;
  tri   n14722;
  tri   n14723;
  tri   P2_N918;
  tri   n14724;
  tri   n14725;
  tri   P2_N919;
  tri   n14726;
  tri   n14727;
  tri   n14703;
  tri   P2_N1260;
  tri   n14704;
  tri   n14705;
  tri   n14706;
  tri   n14708;
  tri   n14709;
  tri   n14711;
  tri   n14710;
  tri   n14712;
  tri   n14713;
  tri   P2_N842;
  tri   P2_N1188;
  tri   n14715;
  tri   P2_N1816;
  tri   P2_N2562;
  tri   P2_N2189;
  tri   P2_N2935;
  tri   P2_N3308;
  tri   P2_N4054;
  tri   P2_N3681;
  tri   P2_N4398;
  tri   n14714;
  tri   n14716;
  tri   n14717;
  tri   P2_N915;
  tri   n14672;
  tri   n14673;
  tri   P2_N1245;
  tri   n14674;
  tri   n14675;
  tri   P2_N1246;
  tri   n14676;
  tri   n14677;
  tri   P2_N1247;
  tri   n14678;
  tri   n14679;
  tri   P2_N1248;
  tri   n14680;
  tri   n14681;
  tri   P2_N1249;
  tri   n14682;
  tri   n14683;
  tri   P2_N1250;
  tri   n14684;
  tri   n14685;
  tri   P2_N1251;
  tri   n14686;
  tri   n14687;
  tri   P2_N1252;
  tri   n14688;
  tri   n14689;
  tri   P2_N1253;
  tri   n14690;
  tri   n14691;
  tri   P2_N1254;
  tri   n14692;
  tri   n14693;
  tri   P2_N1255;
  tri   n14694;
  tri   n14695;
  tri   P2_N1256;
  tri   n14696;
  tri   n14697;
  tri   P2_N1257;
  tri   n14698;
  tri   n14699;
  tri   P2_N1258;
  tri   n14700;
  tri   n14701;
  tri   P2_N1259;
  tri   n14702;
  tri   P2_N4528;
  tri   n14644;
  tri   n14645;
  tri   P2_N1231;
  tri   n14646;
  tri   n14647;
  tri   P2_N1232;
  tri   n14648;
  tri   n14649;
  tri   P2_N1233;
  tri   n14650;
  tri   n14651;
  tri   P2_N1234;
  tri   n14652;
  tri   n14653;
  tri   P2_N1235;
  tri   n14654;
  tri   n14655;
  tri   P2_N1236;
  tri   n14656;
  tri   n14657;
  tri   P2_N1237;
  tri   n14658;
  tri   n14659;
  tri   P2_N1238;
  tri   n14660;
  tri   n14661;
  tri   P2_N1239;
  tri   n14662;
  tri   n14663;
  tri   P2_N1240;
  tri   n14664;
  tri   n14665;
  tri   P2_N1241;
  tri   n14666;
  tri   n14667;
  tri   P2_N1242;
  tri   n14668;
  tri   n14669;
  tri   P2_N1243;
  tri   n14670;
  tri   n14671;
  tri   P2_N1244;
  tri   P2_N4524;
  tri   n14636;
  tri   n14637;
  tri   P2_N656;
  tri   P2_N1002;
  tri   P2_N4525;
  tri   n14638;
  tri   n14639;
  tri   P2_N657;
  tri   P2_N1003;
  tri   P2_N4526;
  tri   n14640;
  tri   n14641;
  tri   P2_N658;
  tri   P2_N1004;
  tri   P2_N4527;
  tri   n14642;
  tri   n14643;
  tri   P2_N659;
  tri   P2_N1005;
  tri   P2_N4520;
  tri   n14628;
  tri   n14629;
  tri   P2_N652;
  tri   P2_N998;
  tri   P2_N4521;
  tri   n14630;
  tri   n14631;
  tri   P2_N653;
  tri   P2_N999;
  tri   P2_N4522;
  tri   n14632;
  tri   n14633;
  tri   P2_N654;
  tri   P2_N1000;
  tri   P2_N4523;
  tri   n14634;
  tri   n14635;
  tri   P2_N655;
  tri   P2_N1001;
  tri   P2_N4516;
  tri   n14620;
  tri   n14621;
  tri   P2_N648;
  tri   P2_N994;
  tri   P2_N4517;
  tri   n14622;
  tri   n14623;
  tri   P2_N649;
  tri   P2_N995;
  tri   P2_N4518;
  tri   n14624;
  tri   n14625;
  tri   P2_N650;
  tri   P2_N996;
  tri   P2_N4519;
  tri   n14626;
  tri   n14627;
  tri   P2_N651;
  tri   P2_N997;
  tri   n14613;
  tri   P2_N644;
  tri   P2_N990;
  tri   P2_N4513;
  tri   n14614;
  tri   n14615;
  tri   P2_N645;
  tri   P2_N991;
  tri   P2_N4514;
  tri   n14616;
  tri   n14617;
  tri   P2_N646;
  tri   P2_N992;
  tri   P2_N4515;
  tri   n14618;
  tri   n14619;
  tri   P2_N647;
  tri   P2_N993;
  tri   P2_N4509;
  tri   n14606;
  tri   n14607;
  tri   P2_N641;
  tri   P2_N987;
  tri   P2_N4510;
  tri   n14608;
  tri   n14609;
  tri   P2_N642;
  tri   P2_N988;
  tri   P2_N4511;
  tri   n14610;
  tri   n14611;
  tri   P2_N643;
  tri   P2_N989;
  tri   P2_N4512;
  tri   n14612;
  tri   P2_N4505;
  tri   n14598;
  tri   n14599;
  tri   P2_N637;
  tri   P2_N983;
  tri   P2_N4506;
  tri   n14600;
  tri   n14601;
  tri   P2_N638;
  tri   P2_N984;
  tri   P2_N4507;
  tri   n14602;
  tri   n14603;
  tri   P2_N639;
  tri   P2_N985;
  tri   P2_N4508;
  tri   n14604;
  tri   n14605;
  tri   P2_N640;
  tri   P2_N986;
  tri   P2_N4501;
  tri   n14590;
  tri   n14591;
  tri   P2_N633;
  tri   P2_N979;
  tri   P2_N4502;
  tri   n14592;
  tri   n14593;
  tri   P2_N634;
  tri   P2_N980;
  tri   P2_N4503;
  tri   n14594;
  tri   n14595;
  tri   P2_N635;
  tri   P2_N981;
  tri   P2_N4504;
  tri   n14596;
  tri   n14597;
  tri   P2_N636;
  tri   P2_N982;
  tri   P2_N4052;
  tri   P2_N3679;
  tri   P2_N4426;
  tri   P2_N4689;
  tri   n14582;
  tri   n14583;
  tri   P2_N841;
  tri   P2_N1187;
  tri   P2_N913;
  tri   P2_N1442;
  tri   P2_N1815;
  tri   P2_N2561;
  tri   P2_N2188;
  tri   P2_N2934;
  tri   P2_N3307;
  tri   P2_N4053;
  tri   P2_N3680;
  tri   P2_N4427;
  tri   P2_N4690;
  tri   n14584;
  tri   n14585;
  tri   P2_N630;
  tri   P2_N976;
  tri   P2_N4499;
  tri   n14586;
  tri   n14587;
  tri   P2_N631;
  tri   P2_N977;
  tri   P2_N4500;
  tri   n14588;
  tri   n14589;
  tri   P2_N632;
  tri   P2_N978;
  tri   P2_N837;
  tri   P2_N1183;
  tri   P2_N909;
  tri   P2_N1438;
  tri   P2_N1811;
  tri   P2_N2557;
  tri   P2_N2184;
  tri   P2_N2930;
  tri   P2_N3303;
  tri   P2_N4049;
  tri   P2_N3676;
  tri   P2_N4423;
  tri   P2_N4686;
  tri   n14576;
  tri   n14577;
  tri   P2_N838;
  tri   P2_N1184;
  tri   P2_N910;
  tri   P2_N1439;
  tri   P2_N1812;
  tri   P2_N2558;
  tri   P2_N2185;
  tri   P2_N2931;
  tri   P2_N3304;
  tri   P2_N4050;
  tri   P2_N3677;
  tri   P2_N4424;
  tri   P2_N4687;
  tri   n14578;
  tri   n14579;
  tri   P2_N839;
  tri   P2_N1185;
  tri   P2_N911;
  tri   P2_N1440;
  tri   P2_N1813;
  tri   P2_N2559;
  tri   P2_N2186;
  tri   P2_N2932;
  tri   P2_N3305;
  tri   P2_N4051;
  tri   P2_N3678;
  tri   P2_N4425;
  tri   P2_N4688;
  tri   n14580;
  tri   n14581;
  tri   P2_N840;
  tri   P2_N1186;
  tri   P2_N912;
  tri   P2_N1441;
  tri   P2_N1814;
  tri   P2_N2560;
  tri   P2_N2187;
  tri   P2_N2933;
  tri   P2_N3306;
  tri   P2_N3299;
  tri   P2_N4045;
  tri   P2_N3672;
  tri   P2_N4419;
  tri   P2_N4682;
  tri   n14568;
  tri   n14569;
  tri   P2_N834;
  tri   P2_N1180;
  tri   P2_N906;
  tri   P2_N1435;
  tri   P2_N1808;
  tri   P2_N2554;
  tri   P2_N2181;
  tri   P2_N2927;
  tri   P2_N3300;
  tri   P2_N4046;
  tri   P2_N3673;
  tri   P2_N4420;
  tri   P2_N4683;
  tri   n14570;
  tri   n14571;
  tri   P2_N835;
  tri   P2_N1181;
  tri   P2_N907;
  tri   P2_N1436;
  tri   P2_N1809;
  tri   P2_N2555;
  tri   P2_N2182;
  tri   P2_N2928;
  tri   P2_N3301;
  tri   P2_N4047;
  tri   P2_N3674;
  tri   P2_N4421;
  tri   P2_N4684;
  tri   n14572;
  tri   n14573;
  tri   P2_N836;
  tri   P2_N1182;
  tri   P2_N908;
  tri   P2_N1437;
  tri   P2_N1810;
  tri   P2_N2556;
  tri   P2_N2183;
  tri   P2_N2929;
  tri   P2_N3302;
  tri   P2_N4048;
  tri   P2_N3675;
  tri   P2_N4422;
  tri   P2_N4685;
  tri   n14574;
  tri   n14575;
  tri   n14560;
  tri   n14561;
  tri   P2_N830;
  tri   P2_N1176;
  tri   P2_N902;
  tri   P2_N1431;
  tri   P2_N1804;
  tri   P2_N2550;
  tri   P2_N2177;
  tri   P2_N2923;
  tri   P2_N3296;
  tri   P2_N4042;
  tri   P2_N3669;
  tri   P2_N4416;
  tri   P2_N4679;
  tri   n14562;
  tri   n14563;
  tri   P2_N831;
  tri   P2_N1177;
  tri   P2_N903;
  tri   P2_N1432;
  tri   P2_N1805;
  tri   P2_N2551;
  tri   P2_N2178;
  tri   P2_N2924;
  tri   P2_N3297;
  tri   P2_N4043;
  tri   P2_N3670;
  tri   P2_N4417;
  tri   P2_N4680;
  tri   n14564;
  tri   n14565;
  tri   P2_N832;
  tri   P2_N1178;
  tri   P2_N904;
  tri   P2_N1433;
  tri   P2_N1806;
  tri   P2_N2552;
  tri   P2_N2179;
  tri   P2_N2925;
  tri   P2_N3298;
  tri   P2_N4044;
  tri   P2_N3671;
  tri   P2_N4418;
  tri   P2_N4681;
  tri   n14566;
  tri   n14567;
  tri   P2_N833;
  tri   P2_N1179;
  tri   P2_N905;
  tri   P2_N1434;
  tri   P2_N1807;
  tri   P2_N2553;
  tri   P2_N2180;
  tri   P2_N2926;
  tri   P2_N2546;
  tri   P2_N2173;
  tri   P2_N2919;
  tri   P2_N3292;
  tri   P2_N4038;
  tri   P2_N3665;
  tri   P2_N4412;
  tri   P2_N4675;
  tri   n14554;
  tri   n14555;
  tri   P2_N827;
  tri   P2_N1173;
  tri   P2_N899;
  tri   P2_N1428;
  tri   P2_N1801;
  tri   P2_N2547;
  tri   P2_N2174;
  tri   P2_N2920;
  tri   P2_N3293;
  tri   P2_N4039;
  tri   P2_N3666;
  tri   P2_N4413;
  tri   P2_N4676;
  tri   n14556;
  tri   n14557;
  tri   P2_N828;
  tri   P2_N1174;
  tri   P2_N900;
  tri   P2_N1429;
  tri   P2_N1802;
  tri   P2_N2548;
  tri   P2_N2175;
  tri   P2_N2921;
  tri   P2_N3294;
  tri   P2_N4040;
  tri   P2_N3667;
  tri   P2_N4414;
  tri   P2_N4677;
  tri   n14558;
  tri   n14559;
  tri   P2_N829;
  tri   P2_N1175;
  tri   P2_N901;
  tri   P2_N1430;
  tri   P2_N1803;
  tri   P2_N2549;
  tri   P2_N2176;
  tri   P2_N2922;
  tri   P2_N3295;
  tri   P2_N4041;
  tri   P2_N3668;
  tri   P2_N4415;
  tri   P2_N4678;
  tri   P2_N4671;
  tri   n14546;
  tri   n14547;
  tri   P2_N823;
  tri   P2_N1169;
  tri   P2_N895;
  tri   P2_N1424;
  tri   P2_N1797;
  tri   P2_N2543;
  tri   P2_N2170;
  tri   P2_N2916;
  tri   P2_N3289;
  tri   P2_N4035;
  tri   P2_N3662;
  tri   P2_N4409;
  tri   P2_N4672;
  tri   n14548;
  tri   n14549;
  tri   P2_N824;
  tri   P2_N1170;
  tri   P2_N896;
  tri   P2_N1425;
  tri   P2_N1798;
  tri   P2_N2544;
  tri   P2_N2171;
  tri   P2_N2917;
  tri   P2_N3290;
  tri   P2_N4036;
  tri   P2_N3663;
  tri   P2_N4410;
  tri   P2_N4673;
  tri   n14550;
  tri   n14551;
  tri   P2_N825;
  tri   P2_N1171;
  tri   P2_N897;
  tri   P2_N1426;
  tri   P2_N1799;
  tri   P2_N2545;
  tri   P2_N2172;
  tri   P2_N2918;
  tri   P2_N3291;
  tri   P2_N4037;
  tri   P2_N3664;
  tri   P2_N4411;
  tri   P2_N4674;
  tri   n14552;
  tri   n14553;
  tri   P2_N826;
  tri   P2_N1172;
  tri   P2_N898;
  tri   P2_N1427;
  tri   P2_N1800;
  tri   P2_N1420;
  tri   P2_N1793;
  tri   P2_N2539;
  tri   P2_N2166;
  tri   P2_N2912;
  tri   P2_N3285;
  tri   P2_N4031;
  tri   P2_N3658;
  tri   P2_N4405;
  tri   P2_N4668;
  tri   n14540;
  tri   n14541;
  tri   P2_N820;
  tri   P2_N1166;
  tri   P2_N892;
  tri   P2_N1421;
  tri   P2_N1794;
  tri   P2_N2540;
  tri   P2_N2167;
  tri   P2_N2913;
  tri   P2_N3286;
  tri   P2_N4032;
  tri   P2_N3659;
  tri   P2_N4406;
  tri   P2_N4669;
  tri   n14542;
  tri   n14543;
  tri   P2_N821;
  tri   P2_N1167;
  tri   P2_N893;
  tri   P2_N1422;
  tri   P2_N1795;
  tri   P2_N2541;
  tri   P2_N2168;
  tri   P2_N2914;
  tri   P2_N3287;
  tri   P2_N4033;
  tri   P2_N3660;
  tri   P2_N4407;
  tri   P2_N4670;
  tri   n14544;
  tri   n14545;
  tri   P2_N822;
  tri   P2_N1168;
  tri   P2_N894;
  tri   P2_N1423;
  tri   P2_N1796;
  tri   P2_N2542;
  tri   P2_N2169;
  tri   P2_N2915;
  tri   P2_N3288;
  tri   P2_N4034;
  tri   P2_N3661;
  tri   P2_N4408;
  tri   P2_N3281;
  tri   P2_N4027;
  tri   P2_N3654;
  tri   P2_N4401;
  tri   P2_N4664;
  tri   n14532;
  tri   n14533;
  tri   P2_N816;
  tri   P2_N1162;
  tri   P2_N888;
  tri   P2_N1417;
  tri   P2_N1790;
  tri   P2_N2536;
  tri   P2_N2163;
  tri   P2_N2909;
  tri   P2_N3282;
  tri   P2_N4028;
  tri   P2_N3655;
  tri   P2_N4402;
  tri   P2_N4665;
  tri   n14534;
  tri   n14535;
  tri   P2_N817;
  tri   P2_N1163;
  tri   P2_N889;
  tri   P2_N1418;
  tri   P2_N1791;
  tri   P2_N2537;
  tri   P2_N2164;
  tri   P2_N2910;
  tri   P2_N3283;
  tri   P2_N4029;
  tri   P2_N3656;
  tri   P2_N4403;
  tri   P2_N4666;
  tri   n14536;
  tri   n14537;
  tri   P2_N818;
  tri   P2_N1164;
  tri   P2_N890;
  tri   P2_N1419;
  tri   P2_N1792;
  tri   P2_N2538;
  tri   P2_N2165;
  tri   P2_N2911;
  tri   P2_N3284;
  tri   P2_N4030;
  tri   P2_N3657;
  tri   P2_N4404;
  tri   P2_N4667;
  tri   n14538;
  tri   n14539;
  tri   P2_N819;
  tri   P2_N1165;
  tri   P2_N891;
  tri   P2_N5206;
  tri   P2_N5210;
  tri   P2_N5208;
  tri   P2_N5212;
  tri   P2_N5214;
  tri   P2_N5285;
  tri   P2_N5216;
  tri   P2_N5354;
  tri   n14526;
  tri   n14527;
  tri   P2_N813;
  tri   P2_N1159;
  tri   P2_N885;
  tri   P2_N1414;
  tri   P2_N1787;
  tri   P2_N2533;
  tri   P2_N2160;
  tri   P2_N2906;
  tri   P2_N3279;
  tri   P2_N4025;
  tri   P2_N3652;
  tri   P2_N4399;
  tri   P2_N4662;
  tri   n14528;
  tri   n14529;
  tri   P2_N814;
  tri   P2_N1160;
  tri   P2_N886;
  tri   P2_N1415;
  tri   P2_N1788;
  tri   P2_N2534;
  tri   P2_N2161;
  tri   P2_N2907;
  tri   P2_N3280;
  tri   P2_N4026;
  tri   P2_N3653;
  tri   P2_N4400;
  tri   P2_N4663;
  tri   n14530;
  tri   n14531;
  tri   P2_N815;
  tri   P2_N1161;
  tri   P2_N887;
  tri   P2_N1416;
  tri   P2_N1789;
  tri   P2_N2535;
  tri   P2_N2162;
  tri   P2_N2908;
  tri   P2_N4838;
  tri   P2_N4778;
  tri   P2_N4779;
  tri   P2_N4780;
  tri   P2_N4781;
  tri   P2_N4782;
  tri   P2_N4783;
  tri   P2_N4784;
  tri   P2_N4785;
  tri   P2_N4786;
  tri   P2_N4787;
  tri   P2_N4788;
  tri   P2_N4789;
  tri   P2_N4790;
  tri   P2_N4791;
  tri   P2_N4792;
  tri   P2_N4793;
  tri   P2_N4794;
  tri   P2_N4795;
  tri   P2_N4796;
  tri   P2_N4797;
  tri   P2_N4798;
  tri   P2_N4799;
  tri   P2_N4800;
  tri   P2_N4801;
  tri   P2_N4802;
  tri   P2_N4803;
  tri   P2_N4804;
  tri   P2_N4805;
  tri   P2_N4806;
  tri   P2_N4807;
  tri   P2_N4745;
  tri   P2_N4746;
  tri   P2_N4747;
  tri   P2_N4748;
  tri   P2_N4749;
  tri   P2_N4750;
  tri   P2_N4751;
  tri   P2_N4752;
  tri   P2_N4753;
  tri   P2_N4754;
  tri   P2_N4755;
  tri   P2_N4756;
  tri   P2_N4757;
  tri   P2_N4758;
  tri   P2_N4759;
  tri   P2_N4760;
  tri   P2_N4761;
  tri   P2_N4762;
  tri   P2_N4763;
  tri   P2_N4764;
  tri   P2_N4765;
  tri   P2_N4766;
  tri   P2_N4767;
  tri   P2_N4768;
  tri   P2_N4769;
  tri   P2_N4770;
  tri   P2_N4771;
  tri   P2_N4772;
  tri   P2_N4773;
  tri   P2_N4774;
  tri   P2_N4777;
  tri   P2_N4744;
  tri   P2_N4661;
  tri   P2_N1443;
  tri   P2_N4713;
  tri   P2_N4693;
  tri   P2_N4694;
  tri   P2_N4695;
  tri   P2_N4696;
  tri   P2_N4697;
  tri   P2_N4698;
  tri   P2_N4699;
  tri   P2_N4700;
  tri   P2_N4701;
  tri   P2_N4702;
  tri   P2_N4703;
  tri   P2_N4704;
  tri   P2_N4705;
  tri   P2_N4706;
  tri   P2_N4707;
  tri   P2_N4708;
  tri   P2_N4709;
  tri   P2_N4710;
  tri   P2_N4711;
  tri   P2_N4712;
  tri   P2_N4692;
  tri   n14524;
  tri   n14525;
  tri   n14348;
  tri   n14346;
  tri   n14359;
  tri   n14351;
  tri   n14350;
  tri   n14355;
  tri   n14353;
  tri   n14352;
  tri   n14357;
  tri   n14356;
  tri   n14354;
  tri   n14361;
  tri   n14360;
  tri   n14358;
  tri   n14370;
  tri   n14363;
  tri   n14362;
  tri   n14367;
  tri   n14365;
  tri   n14364;
  tri   n14369;
  tri   n14368;
  tri   n14366;
  tri   n14371;
  tri   n14373;
  tri   n14372;
  tri   n14377;
  tri   n14375;
  tri   n14374;
  tri   n14379;
  tri   n14378;
  tri   n14376;
  tri   n14389;
  tri   n14381;
  tri   n14380;
  tri   n14385;
  tri   n14383;
  tri   n14382;
  tri   n14387;
  tri   n14386;
  tri   n14384;
  tri   n14391;
  tri   n14390;
  tri   n14388;
  tri   n14400;
  tri   n14393;
  tri   n14392;
  tri   n14397;
  tri   n14395;
  tri   n14394;
  tri   n14399;
  tri   n14398;
  tri   n14396;
  tri   n14401;
  tri   n14403;
  tri   n14402;
  tri   n14407;
  tri   n14405;
  tri   n14404;
  tri   n14409;
  tri   n14408;
  tri   n14406;
  tri   n14419;
  tri   n14411;
  tri   n14410;
  tri   n14415;
  tri   n14413;
  tri   n14412;
  tri   n14417;
  tri   n14416;
  tri   n14414;
  tri   n14421;
  tri   n14420;
  tri   n14418;
  tri   n14430;
  tri   n14423;
  tri   n14422;
  tri   n14427;
  tri   n14425;
  tri   n14424;
  tri   n14429;
  tri   n14428;
  tri   n14426;
  tri   n14431;
  tri   n14433;
  tri   n14432;
  tri   n14437;
  tri   n14435;
  tri   n14434;
  tri   n14439;
  tri   n14438;
  tri   n14436;
  tri   n14449;
  tri   n14441;
  tri   n14440;
  tri   n14445;
  tri   n14443;
  tri   n14442;
  tri   n14447;
  tri   n14446;
  tri   n14444;
  tri   n14451;
  tri   n14450;
  tri   n14448;
  tri   n14460;
  tri   n14453;
  tri   n14452;
  tri   n14457;
  tri   n14455;
  tri   n14454;
  tri   n14459;
  tri   n14458;
  tri   n14456;
  tri   n14461;
  tri   n14463;
  tri   n14462;
  tri   n14467;
  tri   n14465;
  tri   n14464;
  tri   n14469;
  tri   n14468;
  tri   n14466;
  tri   n14479;
  tri   n14471;
  tri   n14470;
  tri   n14475;
  tri   n14473;
  tri   n14472;
  tri   n14477;
  tri   n14476;
  tri   n14474;
  tri   n14481;
  tri   n14480;
  tri   n14478;
  tri   n14490;
  tri   n14483;
  tri   n14482;
  tri   n14487;
  tri   n14485;
  tri   n14484;
  tri   n14489;
  tri   n14488;
  tri   n14486;
  tri   n14491;
  tri   n14493;
  tri   n14492;
  tri   n14497;
  tri   n14495;
  tri   n14494;
  tri   n14499;
  tri   n14498;
  tri   n14496;
  tri   n14509;
  tri   n14501;
  tri   n14500;
  tri   n14505;
  tri   n14503;
  tri   n14502;
  tri   n14507;
  tri   n14506;
  tri   n14504;
  tri   n14511;
  tri   n14510;
  tri   n14508;
  tri   n14520;
  tri   n14514;
  tri   n14513;
  tri   n14517;
  tri   n14516;
  tri   n14512;
  tri   n14519;
  tri   n14515;
  tri   n14518;
  tri   P2_N4810;
  tri   P2_N4811;
  tri   P2_N4812;
  tri   P2_N4813;
  tri   P2_N4814;
  tri   P2_N4815;
  tri   P2_N4816;
  tri   P2_N4817;
  tri   P2_N4818;
  tri   P2_N4819;
  tri   P2_N4820;
  tri   P2_N4821;
  tri   P2_N4822;
  tri   P2_N4823;
  tri   P2_N4824;
  tri   P2_N4825;
  tri   P2_N4826;
  tri   P2_N4827;
  tri   P2_N4828;
  tri   P2_N4829;
  tri   P2_N4830;
  tri   P2_N4831;
  tri   P2_N4832;
  tri   P2_N4833;
  tri   P2_N4834;
  tri   P2_N4835;
  tri   P2_N4836;
  tri   P2_N4837;
  tri   n14068;
  tri   n14066;
  tri   n14071;
  tri   n14073;
  tri   n14072;
  tri   n14077;
  tri   n14075;
  tri   n14074;
  tri   n14079;
  tri   n14078;
  tri   n14076;
  tri   n14089;
  tri   n14081;
  tri   n14080;
  tri   n14085;
  tri   n14083;
  tri   n14082;
  tri   n14087;
  tri   n14086;
  tri   n14084;
  tri   n14091;
  tri   n14090;
  tri   n14088;
  tri   n14100;
  tri   n14093;
  tri   n14092;
  tri   n14097;
  tri   n14095;
  tri   n14094;
  tri   n14099;
  tri   n14098;
  tri   n14096;
  tri   n14101;
  tri   n14103;
  tri   n14102;
  tri   n14107;
  tri   n14105;
  tri   n14104;
  tri   n14109;
  tri   n14108;
  tri   n14106;
  tri   n14119;
  tri   n14111;
  tri   n14110;
  tri   n14115;
  tri   n14113;
  tri   n14112;
  tri   n14117;
  tri   n14116;
  tri   n14114;
  tri   n14121;
  tri   n14120;
  tri   n14118;
  tri   n14130;
  tri   n14123;
  tri   n14122;
  tri   n14127;
  tri   n14125;
  tri   n14124;
  tri   n14129;
  tri   n14128;
  tri   n14126;
  tri   n14131;
  tri   n14133;
  tri   n14132;
  tri   n14137;
  tri   n14135;
  tri   n14134;
  tri   n14139;
  tri   n14138;
  tri   n14136;
  tri   n14149;
  tri   n14141;
  tri   n14140;
  tri   n14145;
  tri   n14143;
  tri   n14142;
  tri   n14147;
  tri   n14146;
  tri   n14144;
  tri   n14151;
  tri   n14150;
  tri   n14148;
  tri   n14160;
  tri   n14153;
  tri   n14152;
  tri   n14157;
  tri   n14155;
  tri   n14154;
  tri   n14159;
  tri   n14158;
  tri   n14156;
  tri   n14161;
  tri   n14163;
  tri   n14162;
  tri   n14167;
  tri   n14165;
  tri   n14164;
  tri   n14169;
  tri   n14168;
  tri   n14166;
  tri   n14179;
  tri   n14171;
  tri   n14170;
  tri   n14175;
  tri   n14173;
  tri   n14172;
  tri   n14177;
  tri   n14176;
  tri   n14174;
  tri   n14181;
  tri   n14180;
  tri   n14178;
  tri   n14190;
  tri   n14183;
  tri   n14182;
  tri   n14187;
  tri   n14185;
  tri   n14184;
  tri   n14189;
  tri   n14188;
  tri   n14186;
  tri   n14191;
  tri   n14193;
  tri   n14192;
  tri   n14197;
  tri   n14195;
  tri   n14194;
  tri   n14199;
  tri   n14198;
  tri   n14196;
  tri   n14209;
  tri   n14201;
  tri   n14200;
  tri   n14205;
  tri   n14203;
  tri   n14202;
  tri   n14207;
  tri   n14206;
  tri   n14204;
  tri   n14211;
  tri   n14210;
  tri   n14208;
  tri   n14220;
  tri   n14213;
  tri   n14212;
  tri   n14217;
  tri   n14215;
  tri   n14214;
  tri   n14219;
  tri   n14218;
  tri   n14216;
  tri   n14221;
  tri   n14223;
  tri   n14222;
  tri   n14227;
  tri   n14225;
  tri   n14224;
  tri   n14229;
  tri   n14228;
  tri   n14226;
  tri   n14239;
  tri   n14231;
  tri   n14230;
  tri   n14235;
  tri   n14233;
  tri   n14232;
  tri   n14237;
  tri   n14236;
  tri   n14234;
  tri   n14241;
  tri   n14240;
  tri   n14238;
  tri   n14250;
  tri   n14243;
  tri   n14242;
  tri   n14247;
  tri   n14245;
  tri   n14244;
  tri   n14249;
  tri   n14248;
  tri   n14246;
  tri   n14251;
  tri   n14253;
  tri   n14252;
  tri   n14257;
  tri   n14255;
  tri   n14254;
  tri   n14259;
  tri   n14258;
  tri   n14256;
  tri   n14269;
  tri   n14261;
  tri   n14260;
  tri   n14265;
  tri   n14263;
  tri   n14262;
  tri   n14267;
  tri   n14266;
  tri   n14264;
  tri   n14271;
  tri   n14270;
  tri   n14268;
  tri   n14280;
  tri   n14273;
  tri   n14272;
  tri   n14277;
  tri   n14275;
  tri   n14274;
  tri   n14279;
  tri   n14278;
  tri   n14276;
  tri   n14281;
  tri   n14283;
  tri   n14282;
  tri   n14287;
  tri   n14285;
  tri   n14284;
  tri   n14289;
  tri   n14288;
  tri   n14286;
  tri   n14299;
  tri   n14291;
  tri   n14290;
  tri   n14295;
  tri   n14293;
  tri   n14292;
  tri   n14297;
  tri   n14296;
  tri   n14294;
  tri   n14301;
  tri   n14300;
  tri   n14298;
  tri   n14310;
  tri   n14303;
  tri   n14302;
  tri   n14307;
  tri   n14305;
  tri   n14304;
  tri   n14309;
  tri   n14308;
  tri   n14306;
  tri   n14311;
  tri   n14313;
  tri   n14312;
  tri   n14317;
  tri   n14315;
  tri   n14314;
  tri   n14319;
  tri   n14318;
  tri   n14316;
  tri   n14329;
  tri   n14321;
  tri   n14320;
  tri   n14325;
  tri   n14323;
  tri   n14322;
  tri   n14327;
  tri   n14326;
  tri   n14324;
  tri   n14331;
  tri   n14330;
  tri   n14328;
  tri   n14340;
  tri   n14333;
  tri   n14332;
  tri   n14337;
  tri   n14335;
  tri   n14334;
  tri   n14339;
  tri   n14338;
  tri   n14336;
  tri   n14341;
  tri   n14343;
  tri   n14342;
  tri   n14347;
  tri   n14345;
  tri   n14344;
  tri   n14349;
  tri   n13790;
  tri   n13789;
  tri   n13793;
  tri   n13792;
  tri   n13791;
  tri   n13794;
  tri   n13796;
  tri   n13795;
  tri   n13799;
  tri   n13798;
  tri   n13797;
  tri   n13800;
  tri   n13802;
  tri   n13801;
  tri   n13804;
  tri   n13805;
  tri   n13803;
  tri   n13816;
  tri   n13808;
  tri   n13807;
  tri   n13812;
  tri   n13810;
  tri   n13809;
  tri   n13814;
  tri   n13813;
  tri   n13811;
  tri   n13818;
  tri   n13817;
  tri   n13815;
  tri   n13830;
  tri   n13820;
  tri   n13819;
  tri   n13824;
  tri   n13822;
  tri   n13821;
  tri   n13826;
  tri   n13825;
  tri   n13823;
  tri   n13828;
  tri   n13829;
  tri   n13827;
  tri   n13831;
  tri   n13833;
  tri   n13832;
  tri   n13835;
  tri   n13836;
  tri   n13834;
  tri   n13846;
  tri   n13838;
  tri   n13837;
  tri   n13842;
  tri   n13840;
  tri   n13839;
  tri   n13844;
  tri   n13843;
  tri   n13841;
  tri   n13848;
  tri   n13847;
  tri   n13845;
  tri   n13860;
  tri   n13850;
  tri   n13849;
  tri   n13854;
  tri   n13852;
  tri   n13851;
  tri   n13856;
  tri   n13855;
  tri   n13853;
  tri   n13858;
  tri   n13859;
  tri   n13857;
  tri   n13861;
  tri   n13863;
  tri   n13862;
  tri   n13865;
  tri   n13866;
  tri   n13864;
  tri   n13876;
  tri   n13868;
  tri   n13867;
  tri   n13872;
  tri   n13870;
  tri   n13869;
  tri   n13874;
  tri   n13873;
  tri   n13871;
  tri   n13878;
  tri   n13877;
  tri   n13875;
  tri   n13890;
  tri   n13880;
  tri   n13879;
  tri   n13884;
  tri   n13882;
  tri   n13881;
  tri   n13886;
  tri   n13885;
  tri   n13883;
  tri   n13888;
  tri   n13889;
  tri   n13887;
  tri   n13891;
  tri   n13893;
  tri   n13892;
  tri   n13897;
  tri   n13895;
  tri   n13894;
  tri   n13899;
  tri   n13898;
  tri   n13896;
  tri   n13909;
  tri   n13901;
  tri   n13900;
  tri   n13905;
  tri   n13903;
  tri   n13902;
  tri   n13907;
  tri   n13906;
  tri   n13904;
  tri   n13911;
  tri   n13910;
  tri   n13908;
  tri   n13920;
  tri   n13913;
  tri   n13912;
  tri   n13917;
  tri   n13915;
  tri   n13914;
  tri   n13919;
  tri   n13918;
  tri   n13916;
  tri   n13921;
  tri   n13923;
  tri   n13922;
  tri   n13927;
  tri   n13925;
  tri   n13924;
  tri   n13929;
  tri   n13928;
  tri   n13926;
  tri   n13939;
  tri   n13931;
  tri   n13930;
  tri   n13935;
  tri   n13933;
  tri   n13932;
  tri   n13937;
  tri   n13936;
  tri   n13934;
  tri   n13941;
  tri   n13940;
  tri   n13938;
  tri   n13950;
  tri   n13943;
  tri   n13942;
  tri   n13947;
  tri   n13945;
  tri   n13944;
  tri   n13949;
  tri   n13948;
  tri   n13946;
  tri   n13951;
  tri   n13953;
  tri   n13952;
  tri   n13957;
  tri   n13955;
  tri   n13954;
  tri   n13959;
  tri   n13958;
  tri   n13956;
  tri   n13969;
  tri   n13961;
  tri   n13960;
  tri   n13965;
  tri   n13963;
  tri   n13962;
  tri   n13967;
  tri   n13966;
  tri   n13964;
  tri   n13971;
  tri   n13970;
  tri   n13968;
  tri   n13980;
  tri   n13973;
  tri   n13972;
  tri   n13977;
  tri   n13975;
  tri   n13974;
  tri   n13979;
  tri   n13978;
  tri   n13976;
  tri   n13981;
  tri   n13983;
  tri   n13982;
  tri   n13987;
  tri   n13985;
  tri   n13984;
  tri   n13989;
  tri   n13988;
  tri   n13986;
  tri   n13999;
  tri   n13991;
  tri   n13990;
  tri   n13995;
  tri   n13993;
  tri   n13992;
  tri   n13997;
  tri   n13996;
  tri   n13994;
  tri   n14001;
  tri   n14000;
  tri   n13998;
  tri   n14010;
  tri   n14003;
  tri   n14002;
  tri   n14007;
  tri   n14005;
  tri   n14004;
  tri   n14009;
  tri   n14008;
  tri   n14006;
  tri   n14011;
  tri   n14013;
  tri   n14012;
  tri   n14017;
  tri   n14015;
  tri   n14014;
  tri   n14019;
  tri   n14018;
  tri   n14016;
  tri   n14029;
  tri   n14021;
  tri   n14020;
  tri   n14025;
  tri   n14023;
  tri   n14022;
  tri   n14027;
  tri   n14026;
  tri   n14024;
  tri   n14031;
  tri   n14030;
  tri   n14028;
  tri   n14040;
  tri   n14033;
  tri   n14032;
  tri   n14037;
  tri   n14035;
  tri   n14034;
  tri   n14039;
  tri   n14038;
  tri   n14036;
  tri   n14041;
  tri   n14043;
  tri   n14042;
  tri   n14047;
  tri   n14045;
  tri   n14044;
  tri   n14049;
  tri   n14048;
  tri   n14046;
  tri   n14059;
  tri   n14051;
  tri   n14050;
  tri   n14055;
  tri   n14053;
  tri   n14052;
  tri   n14057;
  tri   n14056;
  tri   n14054;
  tri   n14061;
  tri   n14060;
  tri   n14058;
  tri   n14070;
  tri   n14063;
  tri   n14062;
  tri   n14067;
  tri   n14065;
  tri   n14064;
  tri   n14069;
  tri   n13510;
  tri   n13509;
  tri   n13514;
  tri   n13512;
  tri   n13511;
  tri   n13516;
  tri   n13515;
  tri   n13513;
  tri   n13519;
  tri   n13518;
  tri   n13517;
  tri   n13521;
  tri   n13523;
  tri   n13522;
  tri   n13527;
  tri   n13525;
  tri   n13524;
  tri   n13529;
  tri   n13528;
  tri   n13526;
  tri   n13539;
  tri   n13531;
  tri   n13530;
  tri   n13535;
  tri   n13533;
  tri   n13532;
  tri   n13537;
  tri   n13536;
  tri   n13534;
  tri   n13541;
  tri   n13540;
  tri   n13538;
  tri   n13553;
  tri   n13543;
  tri   n13542;
  tri   n13547;
  tri   n13545;
  tri   n13544;
  tri   n13549;
  tri   n13548;
  tri   n13546;
  tri   n13552;
  tri   n13551;
  tri   n13550;
  tri   n13554;
  tri   n13556;
  tri   n13555;
  tri   n13560;
  tri   n13558;
  tri   n13557;
  tri   n13562;
  tri   n13561;
  tri   n13559;
  tri   n13572;
  tri   n13564;
  tri   n13563;
  tri   n13568;
  tri   n13566;
  tri   n13565;
  tri   n13570;
  tri   n13569;
  tri   n13567;
  tri   n13574;
  tri   n13573;
  tri   n13571;
  tri   n13586;
  tri   n13576;
  tri   n13575;
  tri   n13580;
  tri   n13578;
  tri   n13577;
  tri   n13582;
  tri   n13581;
  tri   n13579;
  tri   n13585;
  tri   n13584;
  tri   n13583;
  tri   n13587;
  tri   n13589;
  tri   n13588;
  tri   n13593;
  tri   n13591;
  tri   n13590;
  tri   n13595;
  tri   n13594;
  tri   n13592;
  tri   n13605;
  tri   n13597;
  tri   n13596;
  tri   n13601;
  tri   n13599;
  tri   n13598;
  tri   n13603;
  tri   n13602;
  tri   n13600;
  tri   n13607;
  tri   n13606;
  tri   n13604;
  tri   n13619;
  tri   n13609;
  tri   n13608;
  tri   n13613;
  tri   n13611;
  tri   n13610;
  tri   n13615;
  tri   n13614;
  tri   n13612;
  tri   n13618;
  tri   n13617;
  tri   n13616;
  tri   n13620;
  tri   n13622;
  tri   n13621;
  tri   n13625;
  tri   n13624;
  tri   n13623;
  tri   n13626;
  tri   n13628;
  tri   n13627;
  tri   n13631;
  tri   n13630;
  tri   n13629;
  tri   n13632;
  tri   n13634;
  tri   n13633;
  tri   n13637;
  tri   n13636;
  tri   n13635;
  tri   n13638;
  tri   n13640;
  tri   n13639;
  tri   n13643;
  tri   n13642;
  tri   n13641;
  tri   n13644;
  tri   n13646;
  tri   n13645;
  tri   n13649;
  tri   n13648;
  tri   n13647;
  tri   n13650;
  tri   n13652;
  tri   n13651;
  tri   n13655;
  tri   n13654;
  tri   n13653;
  tri   n13656;
  tri   n13658;
  tri   n13657;
  tri   n13661;
  tri   n13660;
  tri   n13659;
  tri   n13662;
  tri   n13664;
  tri   n13663;
  tri   n13667;
  tri   n13666;
  tri   n13665;
  tri   n13668;
  tri   n13670;
  tri   n13669;
  tri   n13673;
  tri   n13672;
  tri   n13671;
  tri   n13674;
  tri   n13676;
  tri   n13675;
  tri   n13679;
  tri   n13678;
  tri   n13677;
  tri   n13680;
  tri   n13682;
  tri   n13681;
  tri   n13685;
  tri   n13684;
  tri   n13683;
  tri   n13686;
  tri   n13688;
  tri   n13687;
  tri   n13691;
  tri   n13690;
  tri   n13689;
  tri   n13692;
  tri   n13694;
  tri   n13693;
  tri   n13697;
  tri   n13696;
  tri   n13695;
  tri   n13698;
  tri   n13700;
  tri   n13699;
  tri   n13703;
  tri   n13702;
  tri   n13701;
  tri   n13704;
  tri   n13706;
  tri   n13705;
  tri   n13709;
  tri   n13708;
  tri   n13707;
  tri   n13710;
  tri   n13712;
  tri   n13711;
  tri   n13715;
  tri   n13714;
  tri   n13713;
  tri   n13716;
  tri   n13718;
  tri   n13717;
  tri   n13721;
  tri   n13720;
  tri   n13719;
  tri   n13722;
  tri   n13724;
  tri   n13723;
  tri   n13727;
  tri   n13726;
  tri   n13725;
  tri   n13728;
  tri   n13730;
  tri   n13729;
  tri   n13733;
  tri   n13732;
  tri   n13731;
  tri   n13734;
  tri   n13736;
  tri   n13735;
  tri   n13739;
  tri   n13738;
  tri   n13737;
  tri   n13740;
  tri   n13742;
  tri   n13741;
  tri   n13745;
  tri   n13744;
  tri   n13743;
  tri   n13746;
  tri   n13748;
  tri   n13747;
  tri   n13751;
  tri   n13750;
  tri   n13749;
  tri   n13752;
  tri   n13754;
  tri   n13753;
  tri   n13757;
  tri   n13756;
  tri   n13755;
  tri   n13758;
  tri   n13760;
  tri   n13759;
  tri   n13763;
  tri   n13762;
  tri   n13761;
  tri   n13764;
  tri   n13766;
  tri   n13765;
  tri   n13769;
  tri   n13768;
  tri   n13767;
  tri   n13770;
  tri   n13772;
  tri   n13771;
  tri   n13775;
  tri   n13774;
  tri   n13773;
  tri   n13776;
  tri   n13778;
  tri   n13777;
  tri   n13781;
  tri   n13780;
  tri   n13779;
  tri   n13782;
  tri   n13784;
  tri   n13783;
  tri   n13787;
  tri   n13786;
  tri   n13785;
  tri   n13788;
  tri   n13231;
  tri   n13229;
  tri   n13242;
  tri   n13234;
  tri   n13233;
  tri   n13238;
  tri   n13236;
  tri   n13235;
  tri   n13240;
  tri   n13239;
  tri   n13237;
  tri   n13244;
  tri   n13243;
  tri   n13241;
  tri   n13256;
  tri   n13246;
  tri   n13245;
  tri   n13250;
  tri   n13248;
  tri   n13247;
  tri   n13252;
  tri   n13251;
  tri   n13249;
  tri   n13255;
  tri   n13254;
  tri   n13253;
  tri   n13257;
  tri   n13259;
  tri   n13258;
  tri   n13263;
  tri   n13261;
  tri   n13260;
  tri   n13265;
  tri   n13264;
  tri   n13262;
  tri   n13275;
  tri   n13267;
  tri   n13266;
  tri   n13271;
  tri   n13269;
  tri   n13268;
  tri   n13273;
  tri   n13272;
  tri   n13270;
  tri   n13277;
  tri   n13276;
  tri   n13274;
  tri   n13289;
  tri   n13279;
  tri   n13278;
  tri   n13283;
  tri   n13281;
  tri   n13280;
  tri   n13285;
  tri   n13284;
  tri   n13282;
  tri   n13288;
  tri   n13287;
  tri   n13286;
  tri   n13290;
  tri   n13292;
  tri   n13291;
  tri   n13296;
  tri   n13294;
  tri   n13293;
  tri   n13298;
  tri   n13297;
  tri   n13295;
  tri   n13308;
  tri   n13300;
  tri   n13299;
  tri   n13304;
  tri   n13302;
  tri   n13301;
  tri   n13306;
  tri   n13305;
  tri   n13303;
  tri   n13310;
  tri   n13309;
  tri   n13307;
  tri   n13322;
  tri   n13312;
  tri   n13311;
  tri   n13316;
  tri   n13314;
  tri   n13313;
  tri   n13318;
  tri   n13317;
  tri   n13315;
  tri   n13321;
  tri   n13320;
  tri   n13319;
  tri   n13323;
  tri   n13325;
  tri   n13324;
  tri   n13329;
  tri   n13327;
  tri   n13326;
  tri   n13331;
  tri   n13330;
  tri   n13328;
  tri   n13341;
  tri   n13333;
  tri   n13332;
  tri   n13337;
  tri   n13335;
  tri   n13334;
  tri   n13339;
  tri   n13338;
  tri   n13336;
  tri   n13343;
  tri   n13342;
  tri   n13340;
  tri   n13355;
  tri   n13345;
  tri   n13344;
  tri   n13349;
  tri   n13347;
  tri   n13346;
  tri   n13351;
  tri   n13350;
  tri   n13348;
  tri   n13354;
  tri   n13353;
  tri   n13352;
  tri   n13356;
  tri   n13358;
  tri   n13357;
  tri   n13362;
  tri   n13360;
  tri   n13359;
  tri   n13364;
  tri   n13363;
  tri   n13361;
  tri   n13374;
  tri   n13366;
  tri   n13365;
  tri   n13370;
  tri   n13368;
  tri   n13367;
  tri   n13372;
  tri   n13371;
  tri   n13369;
  tri   n13376;
  tri   n13375;
  tri   n13373;
  tri   n13388;
  tri   n13378;
  tri   n13377;
  tri   n13382;
  tri   n13380;
  tri   n13379;
  tri   n13384;
  tri   n13383;
  tri   n13381;
  tri   n13387;
  tri   n13386;
  tri   n13385;
  tri   n13389;
  tri   n13391;
  tri   n13390;
  tri   n13395;
  tri   n13393;
  tri   n13392;
  tri   n13397;
  tri   n13396;
  tri   n13394;
  tri   n13407;
  tri   n13399;
  tri   n13398;
  tri   n13403;
  tri   n13401;
  tri   n13400;
  tri   n13405;
  tri   n13404;
  tri   n13402;
  tri   n13409;
  tri   n13408;
  tri   n13406;
  tri   n13421;
  tri   n13411;
  tri   n13410;
  tri   n13415;
  tri   n13413;
  tri   n13412;
  tri   n13417;
  tri   n13416;
  tri   n13414;
  tri   n13420;
  tri   n13419;
  tri   n13418;
  tri   n13422;
  tri   n13424;
  tri   n13423;
  tri   n13428;
  tri   n13426;
  tri   n13425;
  tri   n13430;
  tri   n13429;
  tri   n13427;
  tri   n13440;
  tri   n13432;
  tri   n13431;
  tri   n13436;
  tri   n13434;
  tri   n13433;
  tri   n13438;
  tri   n13437;
  tri   n13435;
  tri   n13442;
  tri   n13441;
  tri   n13439;
  tri   n13454;
  tri   n13444;
  tri   n13443;
  tri   n13448;
  tri   n13446;
  tri   n13445;
  tri   n13450;
  tri   n13449;
  tri   n13447;
  tri   n13453;
  tri   n13452;
  tri   n13451;
  tri   n13455;
  tri   n13457;
  tri   n13456;
  tri   n13461;
  tri   n13459;
  tri   n13458;
  tri   n13463;
  tri   n13462;
  tri   n13460;
  tri   n13473;
  tri   n13465;
  tri   n13464;
  tri   n13469;
  tri   n13467;
  tri   n13466;
  tri   n13471;
  tri   n13470;
  tri   n13468;
  tri   n13475;
  tri   n13474;
  tri   n13472;
  tri   n13487;
  tri   n13477;
  tri   n13476;
  tri   n13481;
  tri   n13479;
  tri   n13478;
  tri   n13483;
  tri   n13482;
  tri   n13480;
  tri   n13486;
  tri   n13485;
  tri   n13484;
  tri   n13488;
  tri   n13490;
  tri   n13489;
  tri   n13494;
  tri   n13492;
  tri   n13491;
  tri   n13496;
  tri   n13495;
  tri   n13493;
  tri   n13506;
  tri   n13498;
  tri   n13497;
  tri   n13502;
  tri   n13500;
  tri   n13499;
  tri   n13504;
  tri   n13503;
  tri   n13501;
  tri   n13508;
  tri   n13507;
  tri   n13505;
  tri   n13520;
  tri   n12951;
  tri   n12950;
  tri   n12955;
  tri   n12954;
  tri   n12952;
  tri   n12958;
  tri   n12957;
  tri   n12956;
  tri   n12960;
  tri   n12962;
  tri   n12961;
  tri   n12966;
  tri   n12964;
  tri   n12963;
  tri   n12968;
  tri   n12967;
  tri   n12965;
  tri   n12978;
  tri   n12970;
  tri   n12969;
  tri   n12974;
  tri   n12972;
  tri   n12971;
  tri   n12976;
  tri   n12975;
  tri   n12973;
  tri   n12980;
  tri   n12979;
  tri   n12977;
  tri   n12992;
  tri   n12982;
  tri   n12981;
  tri   n12986;
  tri   n12984;
  tri   n12983;
  tri   n12988;
  tri   n12987;
  tri   n12985;
  tri   n12991;
  tri   n12990;
  tri   n12989;
  tri   n12993;
  tri   n12995;
  tri   n12994;
  tri   n12999;
  tri   n12997;
  tri   n12996;
  tri   n13001;
  tri   n13000;
  tri   n12998;
  tri   n13011;
  tri   n13003;
  tri   n13002;
  tri   n13007;
  tri   n13005;
  tri   n13004;
  tri   n13009;
  tri   n13008;
  tri   n13006;
  tri   n13013;
  tri   n13012;
  tri   n13010;
  tri   n13025;
  tri   n13015;
  tri   n13014;
  tri   n13019;
  tri   n13017;
  tri   n13016;
  tri   n13021;
  tri   n13020;
  tri   n13018;
  tri   n13024;
  tri   n13023;
  tri   n13022;
  tri   n13026;
  tri   n13028;
  tri   n13027;
  tri   n13032;
  tri   n13030;
  tri   n13029;
  tri   n13034;
  tri   n13033;
  tri   n13031;
  tri   n13044;
  tri   n13036;
  tri   n13035;
  tri   n13040;
  tri   n13038;
  tri   n13037;
  tri   n13042;
  tri   n13041;
  tri   n13039;
  tri   n13046;
  tri   n13045;
  tri   n13043;
  tri   n13058;
  tri   n13048;
  tri   n13047;
  tri   n13052;
  tri   n13050;
  tri   n13049;
  tri   n13054;
  tri   n13053;
  tri   n13051;
  tri   n13057;
  tri   n13056;
  tri   n13055;
  tri   n13059;
  tri   n13061;
  tri   n13060;
  tri   n13065;
  tri   n13063;
  tri   n13062;
  tri   n13067;
  tri   n13066;
  tri   n13064;
  tri   n13077;
  tri   n13069;
  tri   n13068;
  tri   n13073;
  tri   n13071;
  tri   n13070;
  tri   n13075;
  tri   n13074;
  tri   n13072;
  tri   n13079;
  tri   n13078;
  tri   n13076;
  tri   n13091;
  tri   n13081;
  tri   n13080;
  tri   n13085;
  tri   n13083;
  tri   n13082;
  tri   n13087;
  tri   n13086;
  tri   n13084;
  tri   n13090;
  tri   n13089;
  tri   n13088;
  tri   n13092;
  tri   n13094;
  tri   n13093;
  tri   n13098;
  tri   n13096;
  tri   n13095;
  tri   n13100;
  tri   n13099;
  tri   n13097;
  tri   n13110;
  tri   n13102;
  tri   n13101;
  tri   n13106;
  tri   n13104;
  tri   n13103;
  tri   n13108;
  tri   n13107;
  tri   n13105;
  tri   n13112;
  tri   n13111;
  tri   n13109;
  tri   n13124;
  tri   n13114;
  tri   n13113;
  tri   n13118;
  tri   n13116;
  tri   n13115;
  tri   n13120;
  tri   n13119;
  tri   n13117;
  tri   n13123;
  tri   n13122;
  tri   n13121;
  tri   n13125;
  tri   n13127;
  tri   n13126;
  tri   n13131;
  tri   n13129;
  tri   n13128;
  tri   n13133;
  tri   n13132;
  tri   n13130;
  tri   n13143;
  tri   n13135;
  tri   n13134;
  tri   n13139;
  tri   n13137;
  tri   n13136;
  tri   n13141;
  tri   n13140;
  tri   n13138;
  tri   n13145;
  tri   n13144;
  tri   n13142;
  tri   n13157;
  tri   n13147;
  tri   n13146;
  tri   n13151;
  tri   n13149;
  tri   n13148;
  tri   n13153;
  tri   n13152;
  tri   n13150;
  tri   n13156;
  tri   n13155;
  tri   n13154;
  tri   n13158;
  tri   n13160;
  tri   n13159;
  tri   n13164;
  tri   n13162;
  tri   n13161;
  tri   n13166;
  tri   n13165;
  tri   n13163;
  tri   n13176;
  tri   n13168;
  tri   n13167;
  tri   n13172;
  tri   n13170;
  tri   n13169;
  tri   n13174;
  tri   n13173;
  tri   n13171;
  tri   n13178;
  tri   n13177;
  tri   n13175;
  tri   n13190;
  tri   n13180;
  tri   n13179;
  tri   n13184;
  tri   n13182;
  tri   n13181;
  tri   n13186;
  tri   n13185;
  tri   n13183;
  tri   n13189;
  tri   n13188;
  tri   n13187;
  tri   n13191;
  tri   n13193;
  tri   n13192;
  tri   n13197;
  tri   n13195;
  tri   n13194;
  tri   n13199;
  tri   n13198;
  tri   n13196;
  tri   n13209;
  tri   n13201;
  tri   n13200;
  tri   n13205;
  tri   n13203;
  tri   n13202;
  tri   n13207;
  tri   n13206;
  tri   n13204;
  tri   n13211;
  tri   n13210;
  tri   n13208;
  tri   n13223;
  tri   n13213;
  tri   n13212;
  tri   n13217;
  tri   n13215;
  tri   n13214;
  tri   n13219;
  tri   n13218;
  tri   n13216;
  tri   n13222;
  tri   n13221;
  tri   n13220;
  tri   n13224;
  tri   n13226;
  tri   n13225;
  tri   n13230;
  tri   n13228;
  tri   n13227;
  tri   n13232;
  tri   n12673;
  tri   n12672;
  tri   n12677;
  tri   n12675;
  tri   n12674;
  tri   n12679;
  tri   n12678;
  tri   n12676;
  tri   n12683;
  tri   n12682;
  tri   n12680;
  tri   n12695;
  tri   n12685;
  tri   n12684;
  tri   n12689;
  tri   n12687;
  tri   n12686;
  tri   n12691;
  tri   n12690;
  tri   n12688;
  tri   n12694;
  tri   n12693;
  tri   n12692;
  tri   n12696;
  tri   n12698;
  tri   n12697;
  tri   n12702;
  tri   n12700;
  tri   n12699;
  tri   n12704;
  tri   n12703;
  tri   n12701;
  tri   n12714;
  tri   n12706;
  tri   n12705;
  tri   n12710;
  tri   n12708;
  tri   n12707;
  tri   n12712;
  tri   n12711;
  tri   n12709;
  tri   n12716;
  tri   n12715;
  tri   n12713;
  tri   n12728;
  tri   n12718;
  tri   n12717;
  tri   n12722;
  tri   n12720;
  tri   n12719;
  tri   n12724;
  tri   n12723;
  tri   n12721;
  tri   n12727;
  tri   n12726;
  tri   n12725;
  tri   n12729;
  tri   n12731;
  tri   n12730;
  tri   n12735;
  tri   n12733;
  tri   n12732;
  tri   n12737;
  tri   n12736;
  tri   n12734;
  tri   n12747;
  tri   n12739;
  tri   n12738;
  tri   n12743;
  tri   n12741;
  tri   n12740;
  tri   n12745;
  tri   n12744;
  tri   n12742;
  tri   n12749;
  tri   n12748;
  tri   n12746;
  tri   n12761;
  tri   n12751;
  tri   n12750;
  tri   n12755;
  tri   n12753;
  tri   n12752;
  tri   n12757;
  tri   n12756;
  tri   n12754;
  tri   n12760;
  tri   n12759;
  tri   n12758;
  tri   n12762;
  tri   n12764;
  tri   n12763;
  tri   n12768;
  tri   n12766;
  tri   n12765;
  tri   n12770;
  tri   n12769;
  tri   n12767;
  tri   n12780;
  tri   n12772;
  tri   n12771;
  tri   n12776;
  tri   n12774;
  tri   n12773;
  tri   n12778;
  tri   n12777;
  tri   n12775;
  tri   n12782;
  tri   n12781;
  tri   n12779;
  tri   n12794;
  tri   n12784;
  tri   n12783;
  tri   n12788;
  tri   n12786;
  tri   n12785;
  tri   n12790;
  tri   n12789;
  tri   n12787;
  tri   n12793;
  tri   n12792;
  tri   n12791;
  tri   n12795;
  tri   n12797;
  tri   n12796;
  tri   n12801;
  tri   n12799;
  tri   n12798;
  tri   n12803;
  tri   n12802;
  tri   n12800;
  tri   n12813;
  tri   n12805;
  tri   n12804;
  tri   n12809;
  tri   n12807;
  tri   n12806;
  tri   n12811;
  tri   n12810;
  tri   n12808;
  tri   n12815;
  tri   n12814;
  tri   n12812;
  tri   n12827;
  tri   n12817;
  tri   n12816;
  tri   n12821;
  tri   n12819;
  tri   n12818;
  tri   n12823;
  tri   n12822;
  tri   n12820;
  tri   n12826;
  tri   n12825;
  tri   n12824;
  tri   n12828;
  tri   n12830;
  tri   n12829;
  tri   n12834;
  tri   n12832;
  tri   n12831;
  tri   n12836;
  tri   n12835;
  tri   n12833;
  tri   n12846;
  tri   n12838;
  tri   n12837;
  tri   n12842;
  tri   n12840;
  tri   n12839;
  tri   n12844;
  tri   n12843;
  tri   n12841;
  tri   n12848;
  tri   n12847;
  tri   n12845;
  tri   n12860;
  tri   n12850;
  tri   n12849;
  tri   n12854;
  tri   n12852;
  tri   n12851;
  tri   n12856;
  tri   n12855;
  tri   n12853;
  tri   n12859;
  tri   n12858;
  tri   n12857;
  tri   n12861;
  tri   n12863;
  tri   n12862;
  tri   n12867;
  tri   n12865;
  tri   n12864;
  tri   n12869;
  tri   n12868;
  tri   n12866;
  tri   n12879;
  tri   n12871;
  tri   n12870;
  tri   n12875;
  tri   n12873;
  tri   n12872;
  tri   n12877;
  tri   n12876;
  tri   n12874;
  tri   n12881;
  tri   n12880;
  tri   n12878;
  tri   n12893;
  tri   n12883;
  tri   n12882;
  tri   n12887;
  tri   n12885;
  tri   n12884;
  tri   n12889;
  tri   n12888;
  tri   n12886;
  tri   n12892;
  tri   n12891;
  tri   n12890;
  tri   n12894;
  tri   n12896;
  tri   n12895;
  tri   n12900;
  tri   n12898;
  tri   n12897;
  tri   n12902;
  tri   n12901;
  tri   n12899;
  tri   n12912;
  tri   n12904;
  tri   n12903;
  tri   n12908;
  tri   n12906;
  tri   n12905;
  tri   n12910;
  tri   n12909;
  tri   n12907;
  tri   n12914;
  tri   n12913;
  tri   n12911;
  tri   n12926;
  tri   n12916;
  tri   n12915;
  tri   n12920;
  tri   n12918;
  tri   n12917;
  tri   n12922;
  tri   n12921;
  tri   n12919;
  tri   n12925;
  tri   n12924;
  tri   n12923;
  tri   n12927;
  tri   n12929;
  tri   n12928;
  tri   n12933;
  tri   n12931;
  tri   n12930;
  tri   n12935;
  tri   n12934;
  tri   n12932;
  tri   n12945;
  tri   n12937;
  tri   n12936;
  tri   n12941;
  tri   n12939;
  tri   n12938;
  tri   n12943;
  tri   n12942;
  tri   n12940;
  tri   n12947;
  tri   n12946;
  tri   n12944;
  tri   n12959;
  tri   n12949;
  tri   n12948;
  tri   n12953;
  tri   n12393;
  tri   n12391;
  tri   n12398;
  tri   n12397;
  tri   n12395;
  tri   n12413;
  tri   n12400;
  tri   n12399;
  tri   n12404;
  tri   n12402;
  tri   n12401;
  tri   n12406;
  tri   n12405;
  tri   n12403;
  tri   n12410;
  tri   n12408;
  tri   n12407;
  tri   n12412;
  tri   n12411;
  tri   n12409;
  tri   n12414;
  tri   n12416;
  tri   n12415;
  tri   n12420;
  tri   n12418;
  tri   n12417;
  tri   n12422;
  tri   n12421;
  tri   n12419;
  tri   n12432;
  tri   n12424;
  tri   n12423;
  tri   n12428;
  tri   n12426;
  tri   n12425;
  tri   n12430;
  tri   n12429;
  tri   n12427;
  tri   n12434;
  tri   n12433;
  tri   n12431;
  tri   n12449;
  tri   n12436;
  tri   n12435;
  tri   n12440;
  tri   n12438;
  tri   n12437;
  tri   n12442;
  tri   n12441;
  tri   n12439;
  tri   n12446;
  tri   n12444;
  tri   n12443;
  tri   n12448;
  tri   n12447;
  tri   n12445;
  tri   n12450;
  tri   n12452;
  tri   n12451;
  tri   n12456;
  tri   n12454;
  tri   n12453;
  tri   n12458;
  tri   n12457;
  tri   n12455;
  tri   n12468;
  tri   n12460;
  tri   n12459;
  tri   n12464;
  tri   n12462;
  tri   n12461;
  tri   n12466;
  tri   n12465;
  tri   n12463;
  tri   n12470;
  tri   n12469;
  tri   n12467;
  tri   n12485;
  tri   n12472;
  tri   n12471;
  tri   n12476;
  tri   n12474;
  tri   n12473;
  tri   n12478;
  tri   n12477;
  tri   n12475;
  tri   n12482;
  tri   n12480;
  tri   n12479;
  tri   n12484;
  tri   n12483;
  tri   n12481;
  tri   n12486;
  tri   n12488;
  tri   n12487;
  tri   n12492;
  tri   n12490;
  tri   n12489;
  tri   n12494;
  tri   n12493;
  tri   n12491;
  tri   n12504;
  tri   n12496;
  tri   n12495;
  tri   n12500;
  tri   n12498;
  tri   n12497;
  tri   n12502;
  tri   n12501;
  tri   n12499;
  tri   n12506;
  tri   n12505;
  tri   n12503;
  tri   n12521;
  tri   n12508;
  tri   n12507;
  tri   n12512;
  tri   n12510;
  tri   n12509;
  tri   n12514;
  tri   n12513;
  tri   n12511;
  tri   n12518;
  tri   n12516;
  tri   n12515;
  tri   n12520;
  tri   n12519;
  tri   n12517;
  tri   n12522;
  tri   n12524;
  tri   n12523;
  tri   n12528;
  tri   n12526;
  tri   n12525;
  tri   n12530;
  tri   n12529;
  tri   n12527;
  tri   n12540;
  tri   n12532;
  tri   n12531;
  tri   n12536;
  tri   n12534;
  tri   n12533;
  tri   n12538;
  tri   n12537;
  tri   n12535;
  tri   n12542;
  tri   n12541;
  tri   n12539;
  tri   n12557;
  tri   n12544;
  tri   n12543;
  tri   n12548;
  tri   n12546;
  tri   n12545;
  tri   n12550;
  tri   n12549;
  tri   n12547;
  tri   n12554;
  tri   n12552;
  tri   n12551;
  tri   n12556;
  tri   n12555;
  tri   n12553;
  tri   n12558;
  tri   n12560;
  tri   n12559;
  tri   n12564;
  tri   n12562;
  tri   n12561;
  tri   n12566;
  tri   n12565;
  tri   n12563;
  tri   n12576;
  tri   n12568;
  tri   n12567;
  tri   n12572;
  tri   n12570;
  tri   n12569;
  tri   n12574;
  tri   n12573;
  tri   n12571;
  tri   n12578;
  tri   n12577;
  tri   n12575;
  tri   n12593;
  tri   n12580;
  tri   n12579;
  tri   n12584;
  tri   n12582;
  tri   n12581;
  tri   n12586;
  tri   n12585;
  tri   n12583;
  tri   n12590;
  tri   n12588;
  tri   n12587;
  tri   n12592;
  tri   n12591;
  tri   n12589;
  tri   n12594;
  tri   n12596;
  tri   n12595;
  tri   n12600;
  tri   n12598;
  tri   n12597;
  tri   n12602;
  tri   n12601;
  tri   n12599;
  tri   n12612;
  tri   n12604;
  tri   n12603;
  tri   n12608;
  tri   n12606;
  tri   n12605;
  tri   n12610;
  tri   n12609;
  tri   n12607;
  tri   n12614;
  tri   n12613;
  tri   n12611;
  tri   n12629;
  tri   n12616;
  tri   n12615;
  tri   n12620;
  tri   n12618;
  tri   n12617;
  tri   n12622;
  tri   n12621;
  tri   n12619;
  tri   n12626;
  tri   n12624;
  tri   n12623;
  tri   n12628;
  tri   n12627;
  tri   n12625;
  tri   n12630;
  tri   n12632;
  tri   n12631;
  tri   n12636;
  tri   n12634;
  tri   n12633;
  tri   n12638;
  tri   n12637;
  tri   n12635;
  tri   n12648;
  tri   n12640;
  tri   n12639;
  tri   n12644;
  tri   n12642;
  tri   n12641;
  tri   n12646;
  tri   n12645;
  tri   n12643;
  tri   n12650;
  tri   n12649;
  tri   n12647;
  tri   n12662;
  tri   n12652;
  tri   n12651;
  tri   n12656;
  tri   n12654;
  tri   n12653;
  tri   n12658;
  tri   n12657;
  tri   n12655;
  tri   n12661;
  tri   n12660;
  tri   n12659;
  tri   n12663;
  tri   n12665;
  tri   n12664;
  tri   n12669;
  tri   n12667;
  tri   n12666;
  tri   n12671;
  tri   n12670;
  tri   n12668;
  tri   n12681;
  tri   n12114;
  tri   n12113;
  tri   n12118;
  tri   n12117;
  tri   n12115;
  tri   n12122;
  tri   n12120;
  tri   n12119;
  tri   n12124;
  tri   n12123;
  tri   n12121;
  tri   n12126;
  tri   n12128;
  tri   n12127;
  tri   n12132;
  tri   n12130;
  tri   n12129;
  tri   n12134;
  tri   n12133;
  tri   n12131;
  tri   n12144;
  tri   n12136;
  tri   n12135;
  tri   n12140;
  tri   n12138;
  tri   n12137;
  tri   n12142;
  tri   n12141;
  tri   n12139;
  tri   n12146;
  tri   n12145;
  tri   n12143;
  tri   n12161;
  tri   n12148;
  tri   n12147;
  tri   n12152;
  tri   n12150;
  tri   n12149;
  tri   n12154;
  tri   n12153;
  tri   n12151;
  tri   n12158;
  tri   n12156;
  tri   n12155;
  tri   n12160;
  tri   n12159;
  tri   n12157;
  tri   n12162;
  tri   n12164;
  tri   n12163;
  tri   n12168;
  tri   n12166;
  tri   n12165;
  tri   n12170;
  tri   n12169;
  tri   n12167;
  tri   n12180;
  tri   n12172;
  tri   n12171;
  tri   n12176;
  tri   n12174;
  tri   n12173;
  tri   n12178;
  tri   n12177;
  tri   n12175;
  tri   n12182;
  tri   n12181;
  tri   n12179;
  tri   n12197;
  tri   n12184;
  tri   n12183;
  tri   n12188;
  tri   n12186;
  tri   n12185;
  tri   n12190;
  tri   n12189;
  tri   n12187;
  tri   n12194;
  tri   n12192;
  tri   n12191;
  tri   n12196;
  tri   n12195;
  tri   n12193;
  tri   n12198;
  tri   n12200;
  tri   n12199;
  tri   n12204;
  tri   n12202;
  tri   n12201;
  tri   n12206;
  tri   n12205;
  tri   n12203;
  tri   n12216;
  tri   n12208;
  tri   n12207;
  tri   n12212;
  tri   n12210;
  tri   n12209;
  tri   n12214;
  tri   n12213;
  tri   n12211;
  tri   n12218;
  tri   n12217;
  tri   n12215;
  tri   n12233;
  tri   n12220;
  tri   n12219;
  tri   n12224;
  tri   n12222;
  tri   n12221;
  tri   n12226;
  tri   n12225;
  tri   n12223;
  tri   n12230;
  tri   n12228;
  tri   n12227;
  tri   n12232;
  tri   n12231;
  tri   n12229;
  tri   n12234;
  tri   n12236;
  tri   n12235;
  tri   n12240;
  tri   n12238;
  tri   n12237;
  tri   n12242;
  tri   n12241;
  tri   n12239;
  tri   n12252;
  tri   n12244;
  tri   n12243;
  tri   n12248;
  tri   n12246;
  tri   n12245;
  tri   n12250;
  tri   n12249;
  tri   n12247;
  tri   n12254;
  tri   n12253;
  tri   n12251;
  tri   n12269;
  tri   n12256;
  tri   n12255;
  tri   n12260;
  tri   n12258;
  tri   n12257;
  tri   n12262;
  tri   n12261;
  tri   n12259;
  tri   n12266;
  tri   n12264;
  tri   n12263;
  tri   n12268;
  tri   n12267;
  tri   n12265;
  tri   n12270;
  tri   n12272;
  tri   n12271;
  tri   n12276;
  tri   n12274;
  tri   n12273;
  tri   n12278;
  tri   n12277;
  tri   n12275;
  tri   n12288;
  tri   n12280;
  tri   n12279;
  tri   n12284;
  tri   n12282;
  tri   n12281;
  tri   n12286;
  tri   n12285;
  tri   n12283;
  tri   n12290;
  tri   n12289;
  tri   n12287;
  tri   n12305;
  tri   n12292;
  tri   n12291;
  tri   n12296;
  tri   n12294;
  tri   n12293;
  tri   n12298;
  tri   n12297;
  tri   n12295;
  tri   n12302;
  tri   n12300;
  tri   n12299;
  tri   n12304;
  tri   n12303;
  tri   n12301;
  tri   n12306;
  tri   n12308;
  tri   n12307;
  tri   n12312;
  tri   n12310;
  tri   n12309;
  tri   n12314;
  tri   n12313;
  tri   n12311;
  tri   n12324;
  tri   n12316;
  tri   n12315;
  tri   n12320;
  tri   n12318;
  tri   n12317;
  tri   n12322;
  tri   n12321;
  tri   n12319;
  tri   n12326;
  tri   n12325;
  tri   n12323;
  tri   n12341;
  tri   n12328;
  tri   n12327;
  tri   n12332;
  tri   n12330;
  tri   n12329;
  tri   n12334;
  tri   n12333;
  tri   n12331;
  tri   n12338;
  tri   n12336;
  tri   n12335;
  tri   n12340;
  tri   n12339;
  tri   n12337;
  tri   n12342;
  tri   n12344;
  tri   n12343;
  tri   n12348;
  tri   n12346;
  tri   n12345;
  tri   n12350;
  tri   n12349;
  tri   n12347;
  tri   n12360;
  tri   n12352;
  tri   n12351;
  tri   n12356;
  tri   n12354;
  tri   n12353;
  tri   n12358;
  tri   n12357;
  tri   n12355;
  tri   n12362;
  tri   n12361;
  tri   n12359;
  tri   n12377;
  tri   n12364;
  tri   n12363;
  tri   n12368;
  tri   n12366;
  tri   n12365;
  tri   n12370;
  tri   n12369;
  tri   n12367;
  tri   n12374;
  tri   n12372;
  tri   n12371;
  tri   n12376;
  tri   n12375;
  tri   n12373;
  tri   n12378;
  tri   n12380;
  tri   n12379;
  tri   n12384;
  tri   n12382;
  tri   n12381;
  tri   n12386;
  tri   n12385;
  tri   n12383;
  tri   n12396;
  tri   n12388;
  tri   n12387;
  tri   n12392;
  tri   n12390;
  tri   n12389;
  tri   n12394;
  tri   n11835;
  tri   n11833;
  tri   n11838;
  tri   n11840;
  tri   n11839;
  tri   n11844;
  tri   n11842;
  tri   n11841;
  tri   n11846;
  tri   n11845;
  tri   n11843;
  tri   n11856;
  tri   n11848;
  tri   n11847;
  tri   n11852;
  tri   n11850;
  tri   n11849;
  tri   n11854;
  tri   n11853;
  tri   n11851;
  tri   n11858;
  tri   n11857;
  tri   n11855;
  tri   n11873;
  tri   n11860;
  tri   n11859;
  tri   n11864;
  tri   n11862;
  tri   n11861;
  tri   n11866;
  tri   n11865;
  tri   n11863;
  tri   n11870;
  tri   n11868;
  tri   n11867;
  tri   n11872;
  tri   n11871;
  tri   n11869;
  tri   n11874;
  tri   n11876;
  tri   n11875;
  tri   n11880;
  tri   n11878;
  tri   n11877;
  tri   n11882;
  tri   n11881;
  tri   n11879;
  tri   n11892;
  tri   n11884;
  tri   n11883;
  tri   n11888;
  tri   n11886;
  tri   n11885;
  tri   n11890;
  tri   n11889;
  tri   n11887;
  tri   n11894;
  tri   n11893;
  tri   n11891;
  tri   n11909;
  tri   n11896;
  tri   n11895;
  tri   n11900;
  tri   n11898;
  tri   n11897;
  tri   n11902;
  tri   n11901;
  tri   n11899;
  tri   n11906;
  tri   n11904;
  tri   n11903;
  tri   n11908;
  tri   n11907;
  tri   n11905;
  tri   n11910;
  tri   n11912;
  tri   n11911;
  tri   n11916;
  tri   n11914;
  tri   n11913;
  tri   n11918;
  tri   n11917;
  tri   n11915;
  tri   n11928;
  tri   n11920;
  tri   n11919;
  tri   n11924;
  tri   n11922;
  tri   n11921;
  tri   n11926;
  tri   n11925;
  tri   n11923;
  tri   n11930;
  tri   n11929;
  tri   n11927;
  tri   n11945;
  tri   n11932;
  tri   n11931;
  tri   n11936;
  tri   n11934;
  tri   n11933;
  tri   n11938;
  tri   n11937;
  tri   n11935;
  tri   n11942;
  tri   n11940;
  tri   n11939;
  tri   n11944;
  tri   n11943;
  tri   n11941;
  tri   n11946;
  tri   n11948;
  tri   n11947;
  tri   n11952;
  tri   n11950;
  tri   n11949;
  tri   n11954;
  tri   n11953;
  tri   n11951;
  tri   n11964;
  tri   n11956;
  tri   n11955;
  tri   n11960;
  tri   n11958;
  tri   n11957;
  tri   n11962;
  tri   n11961;
  tri   n11959;
  tri   n11966;
  tri   n11965;
  tri   n11963;
  tri   n11981;
  tri   n11968;
  tri   n11967;
  tri   n11972;
  tri   n11970;
  tri   n11969;
  tri   n11974;
  tri   n11973;
  tri   n11971;
  tri   n11978;
  tri   n11976;
  tri   n11975;
  tri   n11980;
  tri   n11979;
  tri   n11977;
  tri   n11982;
  tri   n11984;
  tri   n11983;
  tri   n11988;
  tri   n11986;
  tri   n11985;
  tri   n11990;
  tri   n11989;
  tri   n11987;
  tri   n12000;
  tri   n11992;
  tri   n11991;
  tri   n11996;
  tri   n11994;
  tri   n11993;
  tri   n11998;
  tri   n11997;
  tri   n11995;
  tri   n12002;
  tri   n12001;
  tri   n11999;
  tri   n12017;
  tri   n12004;
  tri   n12003;
  tri   n12008;
  tri   n12006;
  tri   n12005;
  tri   n12010;
  tri   n12009;
  tri   n12007;
  tri   n12014;
  tri   n12012;
  tri   n12011;
  tri   n12016;
  tri   n12015;
  tri   n12013;
  tri   n12018;
  tri   n12020;
  tri   n12019;
  tri   n12024;
  tri   n12022;
  tri   n12021;
  tri   n12026;
  tri   n12025;
  tri   n12023;
  tri   n12036;
  tri   n12028;
  tri   n12027;
  tri   n12032;
  tri   n12030;
  tri   n12029;
  tri   n12034;
  tri   n12033;
  tri   n12031;
  tri   n12038;
  tri   n12037;
  tri   n12035;
  tri   n12053;
  tri   n12040;
  tri   n12039;
  tri   n12044;
  tri   n12042;
  tri   n12041;
  tri   n12046;
  tri   n12045;
  tri   n12043;
  tri   n12050;
  tri   n12048;
  tri   n12047;
  tri   n12052;
  tri   n12051;
  tri   n12049;
  tri   n12054;
  tri   n12056;
  tri   n12055;
  tri   n12060;
  tri   n12058;
  tri   n12057;
  tri   n12062;
  tri   n12061;
  tri   n12059;
  tri   n12072;
  tri   n12064;
  tri   n12063;
  tri   n12068;
  tri   n12066;
  tri   n12065;
  tri   n12070;
  tri   n12069;
  tri   n12067;
  tri   n12074;
  tri   n12073;
  tri   n12071;
  tri   n12089;
  tri   n12076;
  tri   n12075;
  tri   n12080;
  tri   n12078;
  tri   n12077;
  tri   n12082;
  tri   n12081;
  tri   n12079;
  tri   n12086;
  tri   n12084;
  tri   n12083;
  tri   n12088;
  tri   n12087;
  tri   n12085;
  tri   n12090;
  tri   n12092;
  tri   n12091;
  tri   n12096;
  tri   n12094;
  tri   n12093;
  tri   n12098;
  tri   n12097;
  tri   n12095;
  tri   n12108;
  tri   n12100;
  tri   n12099;
  tri   n12104;
  tri   n12102;
  tri   n12101;
  tri   n12106;
  tri   n12105;
  tri   n12103;
  tri   n12110;
  tri   n12109;
  tri   n12107;
  tri   n12125;
  tri   n12112;
  tri   n12111;
  tri   n12116;
  tri   n11555;
  tri   n11554;
  tri   n11559;
  tri   n11558;
  tri   n11556;
  tri   n11563;
  tri   n11562;
  tri   n11560;
  tri   n11585;
  tri   n11565;
  tri   n11564;
  tri   n11569;
  tri   n11567;
  tri   n11566;
  tri   n11571;
  tri   n11570;
  tri   n11568;
  tri   n11581;
  tri   n11573;
  tri   n11572;
  tri   n11577;
  tri   n11575;
  tri   n11574;
  tri   n11579;
  tri   n11578;
  tri   n11576;
  tri   n11583;
  tri   n11582;
  tri   n11580;
  tri   n11586;
  tri   n11588;
  tri   n11587;
  tri   n11592;
  tri   n11590;
  tri   n11589;
  tri   n11594;
  tri   n11593;
  tri   n11591;
  tri   n11604;
  tri   n11596;
  tri   n11595;
  tri   n11600;
  tri   n11598;
  tri   n11597;
  tri   n11602;
  tri   n11601;
  tri   n11599;
  tri   n11606;
  tri   n11605;
  tri   n11603;
  tri   n11621;
  tri   n11608;
  tri   n11607;
  tri   n11612;
  tri   n11610;
  tri   n11609;
  tri   n11614;
  tri   n11613;
  tri   n11611;
  tri   n11618;
  tri   n11616;
  tri   n11615;
  tri   n11620;
  tri   n11619;
  tri   n11617;
  tri   n11622;
  tri   n11624;
  tri   n11623;
  tri   n11628;
  tri   n11626;
  tri   n11625;
  tri   n11630;
  tri   n11629;
  tri   n11627;
  tri   n11640;
  tri   n11632;
  tri   n11631;
  tri   n11636;
  tri   n11634;
  tri   n11633;
  tri   n11638;
  tri   n11637;
  tri   n11635;
  tri   n11642;
  tri   n11641;
  tri   n11639;
  tri   n11657;
  tri   n11644;
  tri   n11643;
  tri   n11648;
  tri   n11646;
  tri   n11645;
  tri   n11650;
  tri   n11649;
  tri   n11647;
  tri   n11654;
  tri   n11652;
  tri   n11651;
  tri   n11656;
  tri   n11655;
  tri   n11653;
  tri   n11658;
  tri   n11660;
  tri   n11659;
  tri   n11664;
  tri   n11662;
  tri   n11661;
  tri   n11666;
  tri   n11665;
  tri   n11663;
  tri   n11676;
  tri   n11668;
  tri   n11667;
  tri   n11672;
  tri   n11670;
  tri   n11669;
  tri   n11674;
  tri   n11673;
  tri   n11671;
  tri   n11678;
  tri   n11677;
  tri   n11675;
  tri   n11693;
  tri   n11680;
  tri   n11679;
  tri   n11684;
  tri   n11682;
  tri   n11681;
  tri   n11686;
  tri   n11685;
  tri   n11683;
  tri   n11690;
  tri   n11688;
  tri   n11687;
  tri   n11692;
  tri   n11691;
  tri   n11689;
  tri   n11694;
  tri   n11696;
  tri   n11695;
  tri   n11700;
  tri   n11698;
  tri   n11697;
  tri   n11702;
  tri   n11701;
  tri   n11699;
  tri   n11712;
  tri   n11704;
  tri   n11703;
  tri   n11708;
  tri   n11706;
  tri   n11705;
  tri   n11710;
  tri   n11709;
  tri   n11707;
  tri   n11714;
  tri   n11713;
  tri   n11711;
  tri   n11729;
  tri   n11716;
  tri   n11715;
  tri   n11720;
  tri   n11718;
  tri   n11717;
  tri   n11722;
  tri   n11721;
  tri   n11719;
  tri   n11726;
  tri   n11724;
  tri   n11723;
  tri   n11728;
  tri   n11727;
  tri   n11725;
  tri   n11730;
  tri   n11732;
  tri   n11731;
  tri   n11736;
  tri   n11734;
  tri   n11733;
  tri   n11738;
  tri   n11737;
  tri   n11735;
  tri   n11748;
  tri   n11740;
  tri   n11739;
  tri   n11744;
  tri   n11742;
  tri   n11741;
  tri   n11746;
  tri   n11745;
  tri   n11743;
  tri   n11750;
  tri   n11749;
  tri   n11747;
  tri   n11765;
  tri   n11752;
  tri   n11751;
  tri   n11756;
  tri   n11754;
  tri   n11753;
  tri   n11758;
  tri   n11757;
  tri   n11755;
  tri   n11762;
  tri   n11760;
  tri   n11759;
  tri   n11764;
  tri   n11763;
  tri   n11761;
  tri   n11766;
  tri   n11768;
  tri   n11767;
  tri   n11772;
  tri   n11770;
  tri   n11769;
  tri   n11774;
  tri   n11773;
  tri   n11771;
  tri   n11784;
  tri   n11776;
  tri   n11775;
  tri   n11780;
  tri   n11778;
  tri   n11777;
  tri   n11782;
  tri   n11781;
  tri   n11779;
  tri   n11786;
  tri   n11785;
  tri   n11783;
  tri   n11801;
  tri   n11788;
  tri   n11787;
  tri   n11792;
  tri   n11790;
  tri   n11789;
  tri   n11794;
  tri   n11793;
  tri   n11791;
  tri   n11798;
  tri   n11796;
  tri   n11795;
  tri   n11800;
  tri   n11799;
  tri   n11797;
  tri   n11802;
  tri   n11804;
  tri   n11803;
  tri   n11808;
  tri   n11806;
  tri   n11805;
  tri   n11810;
  tri   n11809;
  tri   n11807;
  tri   n11820;
  tri   n11812;
  tri   n11811;
  tri   n11816;
  tri   n11814;
  tri   n11813;
  tri   n11818;
  tri   n11817;
  tri   n11815;
  tri   n11822;
  tri   n11821;
  tri   n11819;
  tri   n11837;
  tri   n11824;
  tri   n11823;
  tri   n11828;
  tri   n11826;
  tri   n11825;
  tri   n11830;
  tri   n11829;
  tri   n11827;
  tri   n11834;
  tri   n11832;
  tri   n11831;
  tri   n11836;
  tri   n11537;
  tri   n11538;
  tri   n11539;
  tri   n11540;
  tri   n11541;
  tri   n11542;
  tri   n11543;
  tri   n11544;
  tri   n11546;
  tri   n11547;
  tri   n11545;
  tri   n11548;
  tri   n13806;
  tri   n11551;
  tri   n11549;
  tri   n11561;
  tri   n11553;
  tri   n11552;
  tri   n11557;
  tri   n11529;
  tri   n11530;
  tri   n11531;
  tri   n11532;
  tri   n11533;
  tri   n11534;
  tri   n11535;
  tri   n11536;
  tri   n11521;
  tri   n11522;
  tri   n11523;
  tri   n11524;
  tri   n11525;
  tri   n11526;
  tri   n11527;
  tri   n11528;
  tri   P1_N667;
  tri   n11513;
  tri   n11514;
  tri   n11515;
  tri   n11516;
  tri   n11517;
  tri   n11518;
  tri   n11519;
  tri   n11520;
  tri   n11504;
  tri   n11505;
  tri   n11506;
  tri   n11507;
  tri   n11508;
  tri   P1_N665;
  tri   n11509;
  tri   n11510;
  tri   n11511;
  tri   n11512;
  tri   n11483;
  tri   n11484;
  tri   P1_N1383;
  tri   n11485;
  tri   n11486;
  tri   P1_N1384;
  tri   n11487;
  tri   n11488;
  tri   P1_N1385;
  tri   n11489;
  tri   n11490;
  tri   P1_N1386;
  tri   n11491;
  tri   n11492;
  tri   n11493;
  tri   n11495;
  tri   n11496;
  tri   n11498;
  tri   n11497;
  tri   n11499;
  tri   n11500;
  tri   P1_N968;
  tri   P1_N1314;
  tri   n11502;
  tri   P1_N1942;
  tri   P1_N2688;
  tri   P1_N2315;
  tri   P1_N3061;
  tri   P1_N4180;
  tri   P1_N3807;
  tri   P1_N4553;
  tri   n11501;
  tri   n11503;
  tri   n11452;
  tri   P1_N1367;
  tri   n11453;
  tri   n11454;
  tri   P1_N1368;
  tri   n11455;
  tri   n11456;
  tri   P1_N1369;
  tri   n11457;
  tri   n11458;
  tri   P1_N1370;
  tri   n11459;
  tri   n11460;
  tri   P1_N1371;
  tri   n11461;
  tri   n11462;
  tri   P1_N1372;
  tri   n11463;
  tri   n11464;
  tri   P1_N1373;
  tri   n11465;
  tri   n11466;
  tri   P1_N1374;
  tri   n11467;
  tri   n11468;
  tri   P1_N1375;
  tri   n11469;
  tri   n11470;
  tri   P1_N1376;
  tri   n11471;
  tri   n11472;
  tri   P1_N1377;
  tri   n11473;
  tri   n11474;
  tri   P1_N1378;
  tri   n11475;
  tri   n11476;
  tri   P1_N1379;
  tri   n11477;
  tri   n11478;
  tri   P1_N1380;
  tri   n11479;
  tri   n11480;
  tri   P1_N1381;
  tri   n11481;
  tri   n11482;
  tri   P1_N1382;
  tri   P1_N4653;
  tri   n11429;
  tri   n11430;
  tri   P1_N1131;
  tri   P1_N4654;
  tri   n11431;
  tri   n11432;
  tri   P1_N1357;
  tri   n11433;
  tri   n11434;
  tri   P1_N1358;
  tri   n11435;
  tri   n11436;
  tri   P1_N1359;
  tri   n11437;
  tri   n11438;
  tri   P1_N1360;
  tri   n11439;
  tri   n11440;
  tri   P1_N1361;
  tri   n11441;
  tri   n11442;
  tri   P1_N1362;
  tri   n11443;
  tri   n11444;
  tri   P1_N1363;
  tri   n11445;
  tri   n11446;
  tri   P1_N1364;
  tri   n11447;
  tri   n11448;
  tri   P1_N1365;
  tri   n11449;
  tri   n11450;
  tri   P1_N1366;
  tri   n11451;
  tri   P1_N4649;
  tri   n11421;
  tri   n11422;
  tri   P1_N1127;
  tri   P1_N4650;
  tri   n11423;
  tri   n11424;
  tri   P1_N1128;
  tri   P1_N4651;
  tri   n11425;
  tri   n11426;
  tri   P1_N1129;
  tri   P1_N4652;
  tri   n11427;
  tri   n11428;
  tri   P1_N1130;
  tri   P1_N4645;
  tri   n11413;
  tri   n11414;
  tri   P1_N1123;
  tri   P1_N4646;
  tri   n11415;
  tri   n11416;
  tri   P1_N1124;
  tri   P1_N4647;
  tri   n11417;
  tri   n11418;
  tri   P1_N1125;
  tri   P1_N4648;
  tri   n11419;
  tri   n11420;
  tri   P1_N1126;
  tri   n11406;
  tri   P1_N1119;
  tri   P1_N4642;
  tri   n11407;
  tri   n11408;
  tri   P1_N1120;
  tri   P1_N4643;
  tri   n11409;
  tri   n11410;
  tri   P1_N1121;
  tri   P1_N4644;
  tri   n11411;
  tri   n11412;
  tri   P1_N1122;
  tri   P1_N4638;
  tri   n11399;
  tri   n11400;
  tri   P1_N1116;
  tri   P1_N4639;
  tri   n11401;
  tri   n11402;
  tri   P1_N1117;
  tri   P1_N4640;
  tri   n11403;
  tri   n11404;
  tri   P1_N1118;
  tri   P1_N4641;
  tri   n11405;
  tri   P1_N4634;
  tri   n11391;
  tri   n11392;
  tri   P1_N1112;
  tri   P1_N4635;
  tri   n11393;
  tri   n11394;
  tri   P1_N1113;
  tri   P1_N4636;
  tri   n11395;
  tri   n11396;
  tri   P1_N1114;
  tri   P1_N4637;
  tri   n11397;
  tri   n11398;
  tri   P1_N1115;
  tri   P1_N4630;
  tri   n11383;
  tri   n11384;
  tri   P1_N1108;
  tri   P1_N4631;
  tri   n11385;
  tri   n11386;
  tri   P1_N1109;
  tri   P1_N4632;
  tri   n11387;
  tri   n11388;
  tri   P1_N1110;
  tri   P1_N4633;
  tri   n11389;
  tri   n11390;
  tri   P1_N1111;
  tri   P1_N4626;
  tri   n11375;
  tri   n11376;
  tri   P1_N1104;
  tri   P1_N4627;
  tri   n11377;
  tri   n11378;
  tri   P1_N1105;
  tri   P1_N4628;
  tri   n11379;
  tri   n11380;
  tri   P1_N1106;
  tri   P1_N4629;
  tri   n11381;
  tri   n11382;
  tri   P1_N1107;
  tri   P1_N4813;
  tri   n11367;
  tri   n11368;
  tri   P1_N966;
  tri   P1_N1312;
  tri   P1_N1038;
  tri   P1_N1567;
  tri   P1_N1940;
  tri   P1_N2686;
  tri   P1_N2313;
  tri   P1_N3059;
  tri   P1_N3432;
  tri   P1_N4178;
  tri   P1_N3805;
  tri   P1_N4551;
  tri   P1_N4814;
  tri   n11369;
  tri   n11370;
  tri   P1_N967;
  tri   P1_N1313;
  tri   P1_N1039;
  tri   P1_N1568;
  tri   P1_N1941;
  tri   P1_N2687;
  tri   P1_N2314;
  tri   P1_N3060;
  tri   P1_N3433;
  tri   P1_N4179;
  tri   P1_N3806;
  tri   P1_N4552;
  tri   P1_N4815;
  tri   n11371;
  tri   n11372;
  tri   P1_N1102;
  tri   P1_N4625;
  tri   n11373;
  tri   n11374;
  tri   P1_N1103;
  tri   P1_N1936;
  tri   P1_N2682;
  tri   P1_N2309;
  tri   P1_N3055;
  tri   P1_N3428;
  tri   P1_N4174;
  tri   P1_N3801;
  tri   P1_N4547;
  tri   P1_N4810;
  tri   n11361;
  tri   n11362;
  tri   P1_N963;
  tri   P1_N1309;
  tri   P1_N1035;
  tri   P1_N1564;
  tri   P1_N1937;
  tri   P1_N2683;
  tri   P1_N2310;
  tri   P1_N3056;
  tri   P1_N3429;
  tri   P1_N4175;
  tri   P1_N3802;
  tri   P1_N4548;
  tri   P1_N4811;
  tri   n11363;
  tri   n11364;
  tri   P1_N964;
  tri   P1_N1310;
  tri   P1_N1036;
  tri   P1_N1565;
  tri   P1_N1938;
  tri   P1_N2684;
  tri   P1_N2311;
  tri   P1_N3057;
  tri   P1_N3430;
  tri   P1_N4176;
  tri   P1_N3803;
  tri   P1_N4549;
  tri   P1_N4812;
  tri   n11365;
  tri   n11366;
  tri   P1_N965;
  tri   P1_N1311;
  tri   P1_N1037;
  tri   P1_N1566;
  tri   P1_N1939;
  tri   P1_N2685;
  tri   P1_N2312;
  tri   P1_N3058;
  tri   P1_N3431;
  tri   P1_N4177;
  tri   P1_N3804;
  tri   P1_N4550;
  tri   P1_N3797;
  tri   P1_N4543;
  tri   P1_N4806;
  tri   n11353;
  tri   n11354;
  tri   P1_N959;
  tri   P1_N1305;
  tri   P1_N1031;
  tri   P1_N1560;
  tri   P1_N1933;
  tri   P1_N2679;
  tri   P1_N2306;
  tri   P1_N3052;
  tri   P1_N3425;
  tri   P1_N4171;
  tri   P1_N3798;
  tri   P1_N4544;
  tri   P1_N4807;
  tri   n11355;
  tri   n11356;
  tri   P1_N960;
  tri   P1_N1306;
  tri   P1_N1032;
  tri   P1_N1561;
  tri   P1_N1934;
  tri   P1_N2680;
  tri   P1_N2307;
  tri   P1_N3053;
  tri   P1_N3426;
  tri   P1_N4172;
  tri   P1_N3799;
  tri   P1_N4545;
  tri   P1_N4808;
  tri   n11357;
  tri   n11358;
  tri   P1_N961;
  tri   P1_N1307;
  tri   P1_N1033;
  tri   P1_N1562;
  tri   P1_N1935;
  tri   P1_N2681;
  tri   P1_N2308;
  tri   P1_N3054;
  tri   P1_N3427;
  tri   P1_N4173;
  tri   P1_N3800;
  tri   P1_N4546;
  tri   P1_N4809;
  tri   n11359;
  tri   n11360;
  tri   P1_N962;
  tri   P1_N1308;
  tri   P1_N1034;
  tri   P1_N1563;
  tri   P1_N1301;
  tri   P1_N1027;
  tri   P1_N1556;
  tri   P1_N1929;
  tri   P1_N2675;
  tri   P1_N2302;
  tri   P1_N3048;
  tri   P1_N3421;
  tri   P1_N4167;
  tri   P1_N3794;
  tri   P1_N4540;
  tri   P1_N4803;
  tri   n11347;
  tri   n11348;
  tri   P1_N956;
  tri   P1_N1302;
  tri   P1_N1028;
  tri   P1_N1557;
  tri   P1_N1930;
  tri   P1_N2676;
  tri   P1_N2303;
  tri   P1_N3049;
  tri   P1_N3422;
  tri   P1_N4168;
  tri   P1_N3795;
  tri   P1_N4541;
  tri   P1_N4804;
  tri   n11349;
  tri   n11350;
  tri   P1_N957;
  tri   P1_N1303;
  tri   P1_N1029;
  tri   P1_N1558;
  tri   P1_N1931;
  tri   P1_N2677;
  tri   P1_N2304;
  tri   P1_N3050;
  tri   P1_N3423;
  tri   P1_N4169;
  tri   P1_N3796;
  tri   P1_N4542;
  tri   P1_N4805;
  tri   n11351;
  tri   n11352;
  tri   P1_N958;
  tri   P1_N1304;
  tri   P1_N1030;
  tri   P1_N1559;
  tri   P1_N1932;
  tri   P1_N2678;
  tri   P1_N2305;
  tri   P1_N3051;
  tri   P1_N3424;
  tri   P1_N4170;
  tri   P1_N3417;
  tri   P1_N4163;
  tri   P1_N3790;
  tri   P1_N4536;
  tri   P1_N4799;
  tri   n11339;
  tri   n11340;
  tri   P1_N952;
  tri   P1_N1298;
  tri   P1_N1024;
  tri   P1_N1553;
  tri   P1_N1926;
  tri   P1_N2672;
  tri   P1_N2299;
  tri   P1_N3045;
  tri   P1_N3418;
  tri   P1_N4164;
  tri   P1_N3791;
  tri   P1_N4537;
  tri   P1_N4800;
  tri   n11341;
  tri   n11342;
  tri   P1_N953;
  tri   P1_N1299;
  tri   P1_N1025;
  tri   P1_N1554;
  tri   P1_N1927;
  tri   P1_N2673;
  tri   P1_N2300;
  tri   P1_N3046;
  tri   P1_N3419;
  tri   P1_N4165;
  tri   P1_N3792;
  tri   P1_N4538;
  tri   P1_N4801;
  tri   n11343;
  tri   n11344;
  tri   P1_N954;
  tri   P1_N1300;
  tri   P1_N1026;
  tri   P1_N1555;
  tri   P1_N1928;
  tri   P1_N2674;
  tri   P1_N2301;
  tri   P1_N3047;
  tri   P1_N3420;
  tri   P1_N4166;
  tri   P1_N3793;
  tri   P1_N4539;
  tri   P1_N4802;
  tri   n11345;
  tri   n11346;
  tri   P1_N955;
  tri   n11331;
  tri   n11332;
  tri   P1_N948;
  tri   P1_N1294;
  tri   P1_N1020;
  tri   P1_N1549;
  tri   P1_N1922;
  tri   P1_N2668;
  tri   P1_N2295;
  tri   P1_N3041;
  tri   P1_N3414;
  tri   P1_N4160;
  tri   P1_N3787;
  tri   P1_N4533;
  tri   P1_N4796;
  tri   n11333;
  tri   n11334;
  tri   P1_N949;
  tri   P1_N1295;
  tri   P1_N1021;
  tri   P1_N1550;
  tri   P1_N1923;
  tri   P1_N2669;
  tri   P1_N2296;
  tri   P1_N3042;
  tri   P1_N3415;
  tri   P1_N4161;
  tri   P1_N3788;
  tri   P1_N4534;
  tri   P1_N4797;
  tri   n11335;
  tri   n11336;
  tri   P1_N950;
  tri   P1_N1296;
  tri   P1_N1022;
  tri   P1_N1551;
  tri   P1_N1924;
  tri   P1_N2670;
  tri   P1_N2297;
  tri   P1_N3043;
  tri   P1_N3416;
  tri   P1_N4162;
  tri   P1_N3789;
  tri   P1_N4535;
  tri   P1_N4798;
  tri   n11337;
  tri   n11338;
  tri   P1_N951;
  tri   P1_N1297;
  tri   P1_N1023;
  tri   P1_N1552;
  tri   P1_N1925;
  tri   P1_N2671;
  tri   P1_N2298;
  tri   P1_N3044;
  tri   P1_N2291;
  tri   P1_N3037;
  tri   P1_N3410;
  tri   P1_N4156;
  tri   P1_N3783;
  tri   P1_N4529;
  tri   P1_N4792;
  tri   n11325;
  tri   n11326;
  tri   P1_N945;
  tri   P1_N1291;
  tri   P1_N1017;
  tri   P1_N1546;
  tri   P1_N1919;
  tri   P1_N2665;
  tri   P1_N2292;
  tri   P1_N3038;
  tri   P1_N3411;
  tri   P1_N4157;
  tri   P1_N3784;
  tri   P1_N4530;
  tri   P1_N4793;
  tri   n11327;
  tri   n11328;
  tri   P1_N946;
  tri   P1_N1292;
  tri   P1_N1018;
  tri   P1_N1547;
  tri   P1_N1920;
  tri   P1_N2666;
  tri   P1_N2293;
  tri   P1_N3039;
  tri   P1_N3412;
  tri   P1_N4158;
  tri   P1_N3785;
  tri   P1_N4531;
  tri   P1_N4794;
  tri   n11329;
  tri   n11330;
  tri   P1_N947;
  tri   P1_N1293;
  tri   P1_N1019;
  tri   P1_N1548;
  tri   P1_N1921;
  tri   P1_N2667;
  tri   P1_N2294;
  tri   P1_N3040;
  tri   P1_N3413;
  tri   P1_N4159;
  tri   P1_N3786;
  tri   P1_N4532;
  tri   P1_N4795;
  tri   P1_N4788;
  tri   n11317;
  tri   n11318;
  tri   P1_N941;
  tri   P1_N1287;
  tri   P1_N1013;
  tri   P1_N1542;
  tri   P1_N1915;
  tri   P1_N2661;
  tri   P1_N2288;
  tri   P1_N3034;
  tri   P1_N3407;
  tri   P1_N4153;
  tri   P1_N3780;
  tri   P1_N4526;
  tri   P1_N4789;
  tri   n11319;
  tri   n11320;
  tri   P1_N942;
  tri   P1_N1288;
  tri   P1_N1014;
  tri   P1_N1543;
  tri   P1_N1916;
  tri   P1_N2662;
  tri   P1_N2289;
  tri   P1_N3035;
  tri   P1_N3408;
  tri   P1_N4154;
  tri   P1_N3781;
  tri   P1_N4527;
  tri   P1_N4790;
  tri   n11321;
  tri   n11322;
  tri   P1_N943;
  tri   P1_N1289;
  tri   P1_N1015;
  tri   P1_N1544;
  tri   P1_N1917;
  tri   P1_N2663;
  tri   P1_N2290;
  tri   P1_N3036;
  tri   P1_N3409;
  tri   P1_N4155;
  tri   P1_N3782;
  tri   P1_N4528;
  tri   P1_N4791;
  tri   n11323;
  tri   n11324;
  tri   P1_N944;
  tri   P1_N1290;
  tri   P1_N1016;
  tri   P1_N1545;
  tri   P1_N1918;
  tri   P1_N2664;
  tri   P1_N4822;
  tri   P1_N4823;
  tri   P1_N4824;
  tri   P1_N4825;
  tri   P1_N4826;
  tri   P1_N4827;
  tri   P1_N4828;
  tri   P1_N4829;
  tri   P1_N4830;
  tri   P1_N4831;
  tri   P1_N4832;
  tri   P1_N4833;
  tri   P1_N4834;
  tri   P1_N4835;
  tri   P1_N4836;
  tri   P1_N4837;
  tri   P1_N4838;
  tri   P1_N4818;
  tri   n11311;
  tri   n11312;
  tri   P1_N5284;
  tri   P1_N5288;
  tri   P1_N5286;
  tri   P1_N5290;
  tri   P1_N5292;
  tri   P1_N5363;
  tri   P1_N5294;
  tri   P1_N5432;
  tri   n11313;
  tri   n11314;
  tri   P1_N939;
  tri   P1_N1285;
  tri   P1_N1011;
  tri   P1_N1540;
  tri   P1_N1913;
  tri   P1_N2659;
  tri   P1_N2286;
  tri   P1_N3032;
  tri   P1_N3405;
  tri   P1_N4151;
  tri   P1_N3778;
  tri   P1_N4524;
  tri   P1_N4787;
  tri   n11315;
  tri   n11316;
  tri   P1_N940;
  tri   P1_N1286;
  tri   P1_N1012;
  tri   P1_N1541;
  tri   P1_N1914;
  tri   P1_N2660;
  tri   P1_N2287;
  tri   P1_N3033;
  tri   P1_N3406;
  tri   P1_N4152;
  tri   P1_N3779;
  tri   P1_N4525;
  tri   P1_N4945;
  tri   P1_N4946;
  tri   P1_N4947;
  tri   P1_N4948;
  tri   P1_N4949;
  tri   P1_N4950;
  tri   P1_N4951;
  tri   P1_N4952;
  tri   P1_N4953;
  tri   P1_N4954;
  tri   P1_N4955;
  tri   P1_N4956;
  tri   P1_N4957;
  tri   P1_N4958;
  tri   P1_N4959;
  tri   P1_N4960;
  tri   P1_N4961;
  tri   P1_N4962;
  tri   P1_N4963;
  tri   P1_N4964;
  tri   P1_N4965;
  tri   P1_N4966;
  tri   P1_N4906;
  tri   P1_N4907;
  tri   P1_N4908;
  tri   P1_N4909;
  tri   P1_N4910;
  tri   P1_N4911;
  tri   P1_N4912;
  tri   P1_N4913;
  tri   P1_N4914;
  tri   P1_N4915;
  tri   P1_N4916;
  tri   P1_N4917;
  tri   P1_N4918;
  tri   P1_N4919;
  tri   P1_N4920;
  tri   P1_N4921;
  tri   P1_N4922;
  tri   P1_N4923;
  tri   P1_N4924;
  tri   P1_N4925;
  tri   P1_N4926;
  tri   P1_N4927;
  tri   P1_N4928;
  tri   P1_N4929;
  tri   P1_N4930;
  tri   P1_N4931;
  tri   P1_N4932;
  tri   P1_N4933;
  tri   P1_N4934;
  tri   P1_N4935;
  tri   P1_N4873;
  tri   P1_N4874;
  tri   P1_N4875;
  tri   P1_N4876;
  tri   P1_N4877;
  tri   P1_N4878;
  tri   P1_N4879;
  tri   P1_N4880;
  tri   P1_N4881;
  tri   P1_N4882;
  tri   P1_N4883;
  tri   P1_N4884;
  tri   P1_N4885;
  tri   P1_N4886;
  tri   P1_N4887;
  tri   P1_N4888;
  tri   P1_N4889;
  tri   P1_N4890;
  tri   P1_N4891;
  tri   P1_N4892;
  tri   P1_N4893;
  tri   P1_N4894;
  tri   P1_N4895;
  tri   P1_N4896;
  tri   P1_N4897;
  tri   P1_N4898;
  tri   P1_N4899;
  tri   P1_N4900;
  tri   P1_N4901;
  tri   P1_N4902;
  tri   P1_N4905;
  tri   P1_N4872;
  tri   P1_N4816;
  tri   P1_N1569;
  tri   P1_N4839;
  tri   P1_N4819;
  tri   P1_N4820;
  tri   P1_N4821;
  tri   P1_N4938;
  tri   P1_N4939;
  tri   P1_N4940;
  tri   P1_N4941;
  tri   P1_N4942;
  tri   P1_N4943;
  tri   P1_N4944;
  tri   n10368;
  tri   n10372;
  tri   n10376;
  tri   n10380;
  tri   n18190;
  tri   n10022;
  tri   n10026;
  tri   n10030;
  tri   n10034;
  tri   n10038;
  tri   n10042;
  tri   n10046;
  tri   n10050;
  tri   n10054;
  tri   n10058;
  tri   n10062;
  tri   n10066;
  tri   n10070;
  tri   n10074;
  tri   n10078;
  tri   n10082;
  tri   n10086;
  tri   n10090;
  tri   n10094;
  tri   n10098;
  tri   n18192;
  tri   n18193;
  tri   n10110;
  tri   n18191;
  tri   n10124;
  tri   n10128;
  tri   n10132;
  tri   n10136;
  tri   n10140;
  tri   n10144;
  tri   n10182;
  tri   n10186;
  tri   n10190;
  tri   n10194;
  tri   n9836;
  tri   n9841;
  tri   n9850;
  tri   n9854;
  tri   n9858;
  tri   n9862;
  tri   n9866;
  tri   n9870;
  tri   n9874;
  tri   n9878;
  tri   n9882;
  tri   n9886;
  tri   n9890;
  tri   n9894;
  tri   n9898;
  tri   n9902;
  tri   n9906;
  tri   n9910;
  tri   n9914;
  tri   n9918;
  tri   n9922;
  tri   n9926;
  tri   n9930;
  tri   n9934;
  tri   n9938;
  tri   n9942;
  tri   n9946;
  tri   n9950;
  tri   n9954;
  tri   n9958;
  tri   n9962;
  tri   n9966;
  tri   n9970;
  tri   n9974;
  tri   n9978;
  tri   n9982;
  tri   n9986;
  tri   n9990;
  tri   n9994;
  tri   n9998;
  tri   n10002;
  tri   n10006;
  tri   n10010;
  tri   n10014;
  tri   n10018;
  tri   n9648;
  tri   n9656;
  tri   n9660;
  tri   n9664;
  tri   n9668;
  tri   n9672;
  tri   n9676;
  tri   n9680;
  tri   n9684;
  tri   n9688;
  tri   n9692;
  tri   n9696;
  tri   n9700;
  tri   n9704;
  tri   n9708;
  tri   n9712;
  tri   n9716;
  tri   n9720;
  tri   n9724;
  tri   n9728;
  tri   n18187;
  tri   n9736;
  tri   n9740;
  tri   n9744;
  tri   n9748;
  tri   n9752;
  tri   n9756;
  tri   n9760;
  tri   n9764;
  tri   n9768;
  tri   n9772;
  tri   n9776;
  tri   n9780;
  tri   n9784;
  tri   n9788;
  tri   n9792;
  tri   n9796;
  tri   n9800;
  tri   n9804;
  tri   n9808;
  tri   n9812;
  tri   n9816;
  tri   n9820;
  tri   n9824;
  tri   n9828;
  tri   n9832;
  tri   n9464;
  tri   n9468;
  tri   n9472;
  tri   n9476;
  tri   n9480;
  tri   n9484;
  tri   n9488;
  tri   n9492;
  tri   n18188;
  tri   n9500;
  tri   n9504;
  tri   n9508;
  tri   n9512;
  tri   n9516;
  tri   n9520;
  tri   n9524;
  tri   n9528;
  tri   n9532;
  tri   n9536;
  tri   n9540;
  tri   n9544;
  tri   n9548;
  tri   n9552;
  tri   n9556;
  tri   n9564;
  tri   n9568;
  tri   n9572;
  tri   n9576;
  tri   n9580;
  tri   n9584;
  tri   n9588;
  tri   n9592;
  tri   n9596;
  tri   n18186;
  tri   n9604;
  tri   n9608;
  tri   n9612;
  tri   n9616;
  tri   n9620;
  tri   n9624;
  tri   n9628;
  tri   n9632;
  tri   n9636;
  tri   n9640;
  tri   n9644;
  tri   n9277;
  tri   n9278;
  tri   n9281;
  tri   n9282;
  tri   n9285;
  tri   n9286;
  tri   n9289;
  tri   n9290;
  tri   n9293;
  tri   n9294;
  tri   n9297;
  tri   n9298;
  tri   n9301;
  tri   n9302;
  tri   n9305;
  tri   n9306;
  tri   n9309;
  tri   n9313;
  tri   n9317;
  tri   n9321;
  tri   n9322;
  tri   n9325;
  tri   n18183;
  tri   n9328;
  tri   n9332;
  tri   n9336;
  tri   n9340;
  tri   n9344;
  tri   n9348;
  tri   n9352;
  tri   n9356;
  tri   n9360;
  tri   n9364;
  tri   n9368;
  tri   n9372;
  tri   n9376;
  tri   n9380;
  tri   n9384;
  tri   n9388;
  tri   n9396;
  tri   n9400;
  tri   n9404;
  tri   n9408;
  tri   n9412;
  tri   n9416;
  tri   n9420;
  tri   n9424;
  tri   n9428;
  tri   n9432;
  tri   n9436;
  tri   n9440;
  tri   n9444;
  tri   n9448;
  tri   n18185;
  tri   n9456;
  tri   n9460;
  tri   n9090;
  tri   n9089;
  tri   n9093;
  tri   n9094;
  tri   n9097;
  tri   n9098;
  tri   n9101;
  tri   n9102;
  tri   n9105;
  tri   n9106;
  tri   n9109;
  tri   n9110;
  tri   n9113;
  tri   n9114;
  tri   n9117;
  tri   n9118;
  tri   n9121;
  tri   n9122;
  tri   n9125;
  tri   n9126;
  tri   n9129;
  tri   n9130;
  tri   n9133;
  tri   n9134;
  tri   n9137;
  tri   n9138;
  tri   n9141;
  tri   n9142;
  tri   n9145;
  tri   n9146;
  tri   n9149;
  tri   n9150;
  tri   n9153;
  tri   n9154;
  tri   n9157;
  tri   n9158;
  tri   n9161;
  tri   n9162;
  tri   n9165;
  tri   n9166;
  tri   n9169;
  tri   n9170;
  tri   n9173;
  tri   n9174;
  tri   n9177;
  tri   n9178;
  tri   n9181;
  tri   n9182;
  tri   n9185;
  tri   n9186;
  tri   n9189;
  tri   n9190;
  tri   n9193;
  tri   n9194;
  tri   n9197;
  tri   n9198;
  tri   n9201;
  tri   n9202;
  tri   n9205;
  tri   n9206;
  tri   n9209;
  tri   n9210;
  tri   n9213;
  tri   n9214;
  tri   n9217;
  tri   n9218;
  tri   n9221;
  tri   n9222;
  tri   n9225;
  tri   n9226;
  tri   n9229;
  tri   n9230;
  tri   n9233;
  tri   n9234;
  tri   n9237;
  tri   n9238;
  tri   n9241;
  tri   n9242;
  tri   n9245;
  tri   n9246;
  tri   n9249;
  tri   n9250;
  tri   n9253;
  tri   n9254;
  tri   n9257;
  tri   n9258;
  tri   n9261;
  tri   n9262;
  tri   n9265;
  tri   n9266;
  tri   n9269;
  tri   n9270;
  tri   n9273;
  tri   n9274;
  tri   n8905;
  tri   n8906;
  tri   n8909;
  tri   n8910;
  tri   n8913;
  tri   n8914;
  tri   n8917;
  tri   n8918;
  tri   n8921;
  tri   n8922;
  tri   n8925;
  tri   n8926;
  tri   n8929;
  tri   n8930;
  tri   n8933;
  tri   n8934;
  tri   n8937;
  tri   n8938;
  tri   n8941;
  tri   n8942;
  tri   n8945;
  tri   n8946;
  tri   n8949;
  tri   n8950;
  tri   n8953;
  tri   n8954;
  tri   n8957;
  tri   n8958;
  tri   n8961;
  tri   n8962;
  tri   n8965;
  tri   n8966;
  tri   n8969;
  tri   n8970;
  tri   n8973;
  tri   n8974;
  tri   n8977;
  tri   n8978;
  tri   n8981;
  tri   n8982;
  tri   n8985;
  tri   n8986;
  tri   n8989;
  tri   n8990;
  tri   n8993;
  tri   n8994;
  tri   n8997;
  tri   n8998;
  tri   n9001;
  tri   n9002;
  tri   n9005;
  tri   n9006;
  tri   n9009;
  tri   n9010;
  tri   n9013;
  tri   n9014;
  tri   n9017;
  tri   n9018;
  tri   n9021;
  tri   n9022;
  tri   n9025;
  tri   n9026;
  tri   n9029;
  tri   n9030;
  tri   n9033;
  tri   n9034;
  tri   n9037;
  tri   n9038;
  tri   n9041;
  tri   n9042;
  tri   n9045;
  tri   n9046;
  tri   n9049;
  tri   n9050;
  tri   n9053;
  tri   n9054;
  tri   n9057;
  tri   n9058;
  tri   n9061;
  tri   n9062;
  tri   n9065;
  tri   n9066;
  tri   n9069;
  tri   n9070;
  tri   n9073;
  tri   n9074;
  tri   n9077;
  tri   n9078;
  tri   n9081;
  tri   n9082;
  tri   n9085;
  tri   n9086;
  tri   n6371;
  tri   P2_N196;
  tri   P2_N244;
  tri   n6370;
  tri   n6376;
  tri   n6369;
  tri   n6372;
  tri   n6374;
  tri   n6373;
  tri   P2_N246;
  tri   n6377;
  tri   n6378;
  tri   P2_N194;
  tri   n6380;
  tri   n6379;
  tri   P2_N247;
  tri   n6392;
  tri   P2_N252;
  tri   P2_N290;
  tri   n6391;
  tri   n6386;
  tri   P2_N251;
  tri   n6393;
  tri   n6387;
  tri   n6395;
  tri   n6394;
  tri   n6396;
  tri   P2_N249;
  tri   n6399;
  tri   P2_N190;
  tri   P2_N136;
  tri   n6402;
  tri   P2_N135;
  tri   n6405;
  tri   n6406;
  tri   P2_N504;
  tri   n6407;
  tri   P2_N508;
  tri   n6409;
  tri   P2_N511;
  tri   n6410;
  tri   P2_N514;
  tri   n6411;
  tri   P2_N517;
  tri   n6412;
  tri   P2_N519;
  tri   n6413;
  tri   P2_N455;
  tri   P2_N397;
  tri   n6416;
  tri   P2_N396;
  tri   P1_N247;
  tri   P1_N246;
  tri   n6419;
  tri   P1_N4969;
  tri   n6420;
  tri   P2_N4841;
  tri   n8869;
  tri   n8870;
  tri   n8873;
  tri   n8874;
  tri   n8877;
  tri   n8878;
  tri   n8881;
  tri   n8882;
  tri   n8885;
  tri   n8886;
  tri   n8889;
  tri   n8890;
  tri   n8893;
  tri   n8894;
  tri   n8897;
  tri   n8898;
  tri   n8901;
  tri   n8902;
  tri   n4145;
  tri   n4148;
  tri   n5944;
  tri   n4151;
  tri   n5947;
  tri   n4154;
  tri   n5950;
  tri   n6321;
  tri   P1_N196;
  tri   P1_N244;
  tri   n6320;
  tri   n6326;
  tri   n6319;
  tri   n6322;
  tri   n6324;
  tri   n6323;
  tri   n6327;
  tri   n6328;
  tri   P1_N194;
  tri   n6330;
  tri   n6329;
  tri   n6342;
  tri   P1_N252;
  tri   P1_N290;
  tri   n6341;
  tri   n6336;
  tri   P1_N251;
  tri   n6343;
  tri   n6337;
  tri   n6345;
  tri   n6344;
  tri   n6346;
  tri   P1_N249;
  tri   n6349;
  tri   P1_N190;
  tri   P1_N136;
  tri   n6352;
  tri   P1_N135;
  tri   n6355;
  tri   n6356;
  tri   P1_N504;
  tri   n6357;
  tri   P1_N508;
  tri   n6359;
  tri   P1_N511;
  tri   n6360;
  tri   P1_N514;
  tri   n6361;
  tri   P1_N517;
  tri   n6362;
  tri   P1_N519;
  tri   n6363;
  tri   P1_N455;
  tri   P1_N397;
  tri   n6366;
  tri   P1_N396;
  tri   n4097;
  tri   n4100;
  tri   n5896;
  tri   n4102;
  tri   n5897;
  tri   n5898;
  tri   n4103;
  tri   n5899;
  tri   n4105;
  tri   n5900;
  tri   n5901;
  tri   n4106;
  tri   n5902;
  tri   n4109;
  tri   n5905;
  tri   n5908;
  tri   n5911;
  tri   n5914;
  tri   n5917;
  tri   n5920;
  tri   n5923;
  tri   n4130;
  tri   n5926;
  tri   n4132;
  tri   n5927;
  tri   n5928;
  tri   n4133;
  tri   n5929;
  tri   n4135;
  tri   n5930;
  tri   n5931;
  tri   n5932;
  tri   n4139;
  tri   n5935;
  tri   n4142;
  tri   n5938;
  tri   n5941;
  tri   n5840;
  tri   n5841;
  tri   n5838;
  tri   n5842;
  tri   n5843;
  tri   n5844;
  tri   n5845;
  tri   n5846;
  tri   n5847;
  tri   n5848;
  tri   n5849;
  tri   n5850;
  tri   n5851;
  tri   n5852;
  tri   n5853;
  tri   n5854;
  tri   n5855;
  tri   n5856;
  tri   n5857;
  tri   n5858;
  tri   n5859;
  tri   n5860;
  tri   n5861;
  tri   n5862;
  tri   n5863;
  tri   n5864;
  tri   n5865;
  tri   n5866;
  tri   n5867;
  tri   n5868;
  tri   n5869;
  tri   n5870;
  tri   n5871;
  tri   n5872;
  tri   n5873;
  tri   n5875;
  tri   n5876;
  tri   n5877;
  tri   n5878;
  tri   n5879;
  tri   n5880;
  tri   n5881;
  tri   n5882;
  tri   n5883;
  tri   n5884;
  tri   n5885;
  tri   n5886;
  tri   n5887;
  tri   n5888;
  tri   n5889;
  tri   n5890;
  tri   n5891;
  tri   n5892;
  tri   n5893;
  tri   n5776;
  tri   n5777;
  tri   n5778;
  tri   n5779;
  tri   n5780;
  tri   n5781;
  tri   n5782;
  tri   n5783;
  tri   n5784;
  tri   n5785;
  tri   n5786;
  tri   n5787;
  tri   n5788;
  tri   n5789;
  tri   n5790;
  tri   n5791;
  tri   n5792;
  tri   n5793;
  tri   n5794;
  tri   n5795;
  tri   n5796;
  tri   n5797;
  tri   n5798;
  tri   n5799;
  tri   n5800;
  tri   n5801;
  tri   n5802;
  tri   n5803;
  tri   n5804;
  tri   n5805;
  tri   n5806;
  tri   n5807;
  tri   n5808;
  tri   n5809;
  tri   n5810;
  tri   n5811;
  tri   n5812;
  tri   n5813;
  tri   n5814;
  tri   n5815;
  tri   n5816;
  tri   n5817;
  tri   n5818;
  tri   n5819;
  tri   n5820;
  tri   n5821;
  tri   n5822;
  tri   n5823;
  tri   n5824;
  tri   n5825;
  tri   n5826;
  tri   n5827;
  tri   n5828;
  tri   n5829;
  tri   n5830;
  tri   n5831;
  tri   n5832;
  tri   n5833;
  tri   n5834;
  tri   n5835;
  tri   n5836;
  tri   n5837;
  tri   n5839;
  tri   n5721;
  tri   n5722;
  tri   P1_N5572;
  tri   n5723;
  tri   n5724;
  tri   n5725;
  tri   n5726;
  tri   n5727;
  tri   n5728;
  tri   n5729;
  tri   n5730;
  tri   n5731;
  tri   n5732;
  tri   n5733;
  tri   n5734;
  tri   n5735;
  tri   n5736;
  tri   n5737;
  tri   n5738;
  tri   n5739;
  tri   n5740;
  tri   n5741;
  tri   n5742;
  tri   n5743;
  tri   n5744;
  tri   n5745;
  tri   n5746;
  tri   n5747;
  tri   n5748;
  tri   n5749;
  tri   n5750;
  tri   n5751;
  tri   n5752;
  tri   n5753;
  tri   n5754;
  tri   n5755;
  tri   n5756;
  tri   n5757;
  tri   n5758;
  tri   n5759;
  tri   n5760;
  tri   n5761;
  tri   n5762;
  tri   n5763;
  tri   n5764;
  tri   n5765;
  tri   n5766;
  tri   n5769;
  tri   n5770;
  tri   n5772;
  tri   n5773;
  tri   n5774;
  tri   n5775;
  tri   P1_N5573;
  tri   n5667;
  tri   n5669;
  tri   n5670;
  tri   n5671;
  tri   n5672;
  tri   n5673;
  tri   n5674;
  tri   n5675;
  tri   n5676;
  tri   n5677;
  tri   n5678;
  tri   n5679;
  tri   n5680;
  tri   n5683;
  tri   n5684;
  tri   n5686;
  tri   n5687;
  tri   n5688;
  tri   n5689;
  tri   n5690;
  tri   n5691;
  tri   n5692;
  tri   n5693;
  tri   n5694;
  tri   n5695;
  tri   n5696;
  tri   n5697;
  tri   n5698;
  tri   n5699;
  tri   n5700;
  tri   n5701;
  tri   n5702;
  tri   n5703;
  tri   n5704;
  tri   n5705;
  tri   n5707;
  tri   n5708;
  tri   n5711;
  tri   n5712;
  tri   n5713;
  tri   n5714;
  tri   n5715;
  tri   n5716;
  tri   n5717;
  tri   n5718;
  tri   n5719;
  tri   n5720;
  tri   n5607;
  tri   n5608;
  tri   n5609;
  tri   n5610;
  tri   n5611;
  tri   n5612;
  tri   n5613;
  tri   n5614;
  tri   n5615;
  tri   n5616;
  tri   n5617;
  tri   n5618;
  tri   n5619;
  tri   n5621;
  tri   n5622;
  tri   n5625;
  tri   n5626;
  tri   n5627;
  tri   n5628;
  tri   n5629;
  tri   n5630;
  tri   n5631;
  tri   n5632;
  tri   n5633;
  tri   n5634;
  tri   n5635;
  tri   n5636;
  tri   n5637;
  tri   n5638;
  tri   n5639;
  tri   n5640;
  tri   n5641;
  tri   n5642;
  tri   n5643;
  tri   n5644;
  tri   n5645;
  tri   n5646;
  tri   n5647;
  tri   n5648;
  tri   n5649;
  tri   n5650;
  tri   n5651;
  tri   n5652;
  tri   n5653;
  tri   n5654;
  tri   n5655;
  tri   n5656;
  tri   n5657;
  tri   n5658;
  tri   n5659;
  tri   n5660;
  tri   n5661;
  tri   n5662;
  tri   n5663;
  tri   n5664;
  tri   n5665;
  tri   n5666;
  tri   n5668;
  tri   n5546;
  tri   P1_N5577;
  tri   n5545;
  tri   n5547;
  tri   n5548;
  tri   n5549;
  tri   n5550;
  tri   n5551;
  tri   n5552;
  tri   n5553;
  tri   n5554;
  tri   n5555;
  tri   n5556;
  tri   n5557;
  tri   n5558;
  tri   n5559;
  tri   n5560;
  tri   n5561;
  tri   n5562;
  tri   n5563;
  tri   n5564;
  tri   n5565;
  tri   n5566;
  tri   n5567;
  tri   n5568;
  tri   P1_N134;
  tri   n5571;
  tri   n5572;
  tri   n5573;
  tri   n5574;
  tri   n5575;
  tri   n5576;
  tri   n5577;
  tri   n5578;
  tri   n5579;
  tri   P1_N156;
  tri   P1_N155;
  tri   P1_N154;
  tri   P1_N153;
  tri   P1_N150;
  tri   n5580;
  tri   P1_N151;
  tri   P1_N152;
  tri   n5581;
  tri   n5582;
  tri   n5583;
  tri   n5584;
  tri   P1_N163;
  tri   P1_N162;
  tri   P1_N161;
  tri   P1_N160;
  tri   P1_N157;
  tri   n5585;
  tri   P1_N158;
  tri   P1_N159;
  tri   n5586;
  tri   n5587;
  tri   n5588;
  tri   n5589;
  tri   P1_N140;
  tri   n5590;
  tri   P1_N141;
  tri   P1_N142;
  tri   P1_N137;
  tri   n5591;
  tri   P1_N138;
  tri   P1_N139;
  tri   n5592;
  tri   n5593;
  tri   n5594;
  tri   n5595;
  tri   P1_N149;
  tri   P1_N148;
  tri   P1_N147;
  tri   P1_N146;
  tri   P1_N143;
  tri   n5596;
  tri   P1_N144;
  tri   P1_N145;
  tri   n5597;
  tri   n5598;
  tri   n5600;
  tri   n5601;
  tri   n5602;
  tri   n5603;
  tri   n5604;
  tri   n5605;
  tri   n5606;
  tri   n5488;
  tri   n5489;
  tri   n5490;
  tri   n5491;
  tri   n5492;
  tri   n5493;
  tri   n5494;
  tri   n5495;
  tri   n5496;
  tri   n5497;
  tri   n5498;
  tri   n5499;
  tri   n5500;
  tri   n5501;
  tri   n5502;
  tri   n5503;
  tri   n5504;
  tri   n5505;
  tri   n5506;
  tri   n5507;
  tri   n5509;
  tri   n5510;
  tri   n5513;
  tri   n5514;
  tri   n5515;
  tri   n5516;
  tri   n5517;
  tri   n5518;
  tri   n5519;
  tri   n5520;
  tri   n5521;
  tri   n5522;
  tri   n5523;
  tri   n5524;
  tri   n5525;
  tri   n5526;
  tri   n5527;
  tri   n5528;
  tri   n5529;
  tri   n5530;
  tri   n5531;
  tri   n5532;
  tri   n5533;
  tri   n5534;
  tri   n5535;
  tri   n5536;
  tri   n5537;
  tri   n5538;
  tri   n5539;
  tri   n5540;
  tri   n5541;
  tri   n5542;
  tri   n5543;
  tri   n5544;
  tri   n5431;
  tri   n5432;
  tri   P1_N5578;
  tri   n5433;
  tri   n5434;
  tri   n5435;
  tri   n5436;
  tri   n5437;
  tri   n5438;
  tri   n5439;
  tri   n5440;
  tri   n5441;
  tri   n5442;
  tri   n5443;
  tri   n5444;
  tri   n5445;
  tri   n5446;
  tri   n5447;
  tri   n5448;
  tri   n5449;
  tri   n5450;
  tri   n5451;
  tri   n5452;
  tri   n5453;
  tri   n5454;
  tri   n5455;
  tri   n5456;
  tri   n5457;
  tri   n5458;
  tri   n5459;
  tri   n5460;
  tri   n5461;
  tri   n5462;
  tri   n5463;
  tri   n5464;
  tri   n5465;
  tri   n5466;
  tri   n5467;
  tri   n5468;
  tri   n5469;
  tri   n5470;
  tri   n5471;
  tri   n5472;
  tri   n5473;
  tri   n5474;
  tri   n5475;
  tri   n5476;
  tri   n5477;
  tri   n5478;
  tri   n5479;
  tri   n5480;
  tri   n5481;
  tri   n5482;
  tri   n5485;
  tri   n5486;
  tri   P1_N5579;
  tri   n5370;
  tri   n5372;
  tri   n5373;
  tri   n5376;
  tri   n5377;
  tri   P1_N193;
  tri   n5378;
  tri   n5379;
  tri   n5380;
  tri   n5381;
  tri   n5382;
  tri   n5383;
  tri   n5384;
  tri   P1_N212;
  tri   n5385;
  tri   P1_N213;
  tri   P1_N214;
  tri   P1_N209;
  tri   n5386;
  tri   P1_N210;
  tri   P1_N211;
  tri   n5387;
  tri   n5388;
  tri   P1_N218;
  tri   n5389;
  tri   P1_N219;
  tri   P1_N220;
  tri   P1_N215;
  tri   n5390;
  tri   P1_N216;
  tri   P1_N217;
  tri   n5391;
  tri   n5392;
  tri   n5393;
  tri   n5394;
  tri   P1_N200;
  tri   n5395;
  tri   P1_N201;
  tri   P1_N202;
  tri   P1_N197;
  tri   n5396;
  tri   P1_N198;
  tri   P1_N199;
  tri   n5397;
  tri   n5398;
  tri   P1_N206;
  tri   n5399;
  tri   P1_N207;
  tri   P1_N208;
  tri   P1_N203;
  tri   n5400;
  tri   P1_N204;
  tri   P1_N205;
  tri   n5402;
  tri   n5403;
  tri   n5404;
  tri   n5405;
  tri   n5406;
  tri   n5407;
  tri   n5408;
  tri   n5409;
  tri   n5410;
  tri   n5411;
  tri   n5412;
  tri   n5413;
  tri   n5414;
  tri   n5415;
  tri   n5416;
  tri   n5417;
  tri   n5418;
  tri   n5419;
  tri   n5420;
  tri   n5421;
  tri   n5423;
  tri   n5424;
  tri   n5427;
  tri   n5428;
  tri   n5429;
  tri   n5430;
  tri   n5308;
  tri   n5309;
  tri   n5310;
  tri   n5311;
  tri   n5312;
  tri   n5314;
  tri   n5315;
  tri   n5318;
  tri   n5319;
  tri   n5320;
  tri   n5321;
  tri   n5322;
  tri   n5323;
  tri   n5324;
  tri   n5325;
  tri   n5326;
  tri   n5327;
  tri   n5328;
  tri   n5329;
  tri   n5330;
  tri   n5331;
  tri   n5332;
  tri   n5333;
  tri   n5334;
  tri   n5335;
  tri   n5336;
  tri   n5337;
  tri   n5338;
  tri   n5339;
  tri   n5340;
  tri   n5341;
  tri   n5342;
  tri   n5343;
  tri   n5344;
  tri   n5345;
  tri   n5346;
  tri   n5347;
  tri   n5348;
  tri   n5349;
  tri   n5350;
  tri   n5351;
  tri   n5352;
  tri   n5353;
  tri   n5354;
  tri   n5355;
  tri   n5356;
  tri   n5357;
  tri   n5358;
  tri   n5359;
  tri   n5360;
  tri   n5361;
  tri   n5362;
  tri   n5363;
  tri   n5364;
  tri   n5365;
  tri   n5366;
  tri   n5367;
  tri   n5368;
  tri   n5369;
  tri   n5371;
  tri   P1_N5580;
  tri   n5250;
  tri   n5252;
  tri   n5253;
  tri   n5254;
  tri   n5255;
  tri   n5256;
  tri   n5257;
  tri   n5258;
  tri   n5259;
  tri   n5260;
  tri   n5261;
  tri   n5262;
  tri   n5263;
  tri   n5264;
  tri   n5265;
  tri   n5266;
  tri   n5267;
  tri   n5268;
  tri   n5269;
  tri   P1_N248;
  tri   n5272;
  tri   n5273;
  tri   n5274;
  tri   n5275;
  tri   n5276;
  tri   n5277;
  tri   n5278;
  tri   P1_N264;
  tri   n5279;
  tri   P1_N265;
  tri   P1_N266;
  tri   P1_N263;
  tri   P1_N262;
  tri   n5280;
  tri   n5281;
  tri   P1_N269;
  tri   n5282;
  tri   P1_N270;
  tri   P1_N271;
  tri   P1_N268;
  tri   P1_N267;
  tri   n5283;
  tri   n5284;
  tri   n5285;
  tri   n5286;
  tri   P1_N256;
  tri   P1_N255;
  tri   P1_N254;
  tri   P1_N253;
  tri   n5287;
  tri   n5288;
  tri   P1_N259;
  tri   n5289;
  tri   P1_N260;
  tri   P1_N261;
  tri   P1_N258;
  tri   P1_N257;
  tri   n5290;
  tri   n5291;
  tri   n5293;
  tri   n5294;
  tri   n5295;
  tri   n5296;
  tri   n5297;
  tri   n5298;
  tri   n5299;
  tri   n5300;
  tri   n5301;
  tri   n5302;
  tri   n5303;
  tri   n5304;
  tri   n5305;
  tri   n5306;
  tri   n5307;
  tri   n5192;
  tri   n5193;
  tri   n5194;
  tri   n5195;
  tri   n5196;
  tri   n5197;
  tri   n5198;
  tri   n5199;
  tri   n5200;
  tri   n5201;
  tri   n5202;
  tri   n5203;
  tri   n5204;
  tri   n5205;
  tri   n5206;
  tri   n5207;
  tri   n5208;
  tri   n5210;
  tri   n5211;
  tri   n5214;
  tri   n5215;
  tri   n5216;
  tri   n5217;
  tri   n5218;
  tri   n5219;
  tri   n5220;
  tri   n5221;
  tri   n5222;
  tri   n5223;
  tri   n5224;
  tri   n5225;
  tri   n5226;
  tri   n5227;
  tri   n5228;
  tri   n5229;
  tri   n5230;
  tri   n5231;
  tri   n5232;
  tri   n5233;
  tri   n5234;
  tri   n5235;
  tri   n5236;
  tri   n5237;
  tri   n5238;
  tri   n5239;
  tri   n5240;
  tri   n5241;
  tri   n5242;
  tri   n5243;
  tri   n5244;
  tri   n5245;
  tri   n5246;
  tri   n5247;
  tri   n5248;
  tri   n5249;
  tri   n5251;
  tri   n5130;
  tri   n5131;
  tri   P1_N295;
  tri   n5132;
  tri   P1_N342;
  tri   n5133;
  tri   n5134;
  tri   n5135;
  tri   n5136;
  tri   n5137;
  tri   n5138;
  tri   P1_N311;
  tri   n5139;
  tri   P1_N312;
  tri   P1_N313;
  tri   P1_N308;
  tri   n5140;
  tri   P1_N309;
  tri   P1_N310;
  tri   n5141;
  tri   n5142;
  tri   P1_N317;
  tri   n5143;
  tri   P1_N318;
  tri   P1_N319;
  tri   P1_N314;
  tri   n5144;
  tri   P1_N315;
  tri   P1_N316;
  tri   n5145;
  tri   n5146;
  tri   n5147;
  tri   n5148;
  tri   P1_N299;
  tri   n5149;
  tri   P1_N300;
  tri   P1_N301;
  tri   P1_N298;
  tri   P1_N297;
  tri   n5150;
  tri   n5151;
  tri   P1_N305;
  tri   n5152;
  tri   P1_N306;
  tri   P1_N307;
  tri   P1_N302;
  tri   n5153;
  tri   P1_N303;
  tri   P1_N304;
  tri   n5154;
  tri   n5155;
  tri   n5156;
  tri   n5157;
  tri   n5158;
  tri   n5159;
  tri   n5160;
  tri   n5161;
  tri   n5162;
  tri   n5163;
  tri   n5164;
  tri   n5165;
  tri   n5166;
  tri   n5167;
  tri   n5168;
  tri   n5169;
  tri   n5170;
  tri   n5171;
  tri   n5172;
  tri   n5173;
  tri   n5174;
  tri   n5175;
  tri   n5176;
  tri   n5177;
  tri   n5178;
  tri   n5179;
  tri   n5180;
  tri   n5181;
  tri   n5182;
  tri   n5183;
  tri   n5186;
  tri   n5187;
  tri   n5189;
  tri   n5190;
  tri   n5191;
  tri   n5079;
  tri   n5078;
  tri   n5081;
  tri   n5082;
  tri   n5083;
  tri   n5084;
  tri   n5085;
  tri   n5086;
  tri   n5087;
  tri   n5088;
  tri   n5089;
  tri   n5090;
  tri   n5091;
  tri   n5092;
  tri   n5093;
  tri   n5094;
  tri   n5095;
  tri   n5096;
  tri   n5097;
  tri   n5098;
  tri   n5099;
  tri   n5100;
  tri   n5102;
  tri   n5103;
  tri   n5106;
  tri   n5107;
  tri   n5108;
  tri   n5109;
  tri   n5110;
  tri   n5111;
  tri   n5112;
  tri   n5113;
  tri   n5114;
  tri   n5115;
  tri   n5116;
  tri   n5117;
  tri   n5118;
  tri   n5119;
  tri   n5120;
  tri   n5121;
  tri   n5122;
  tri   n5123;
  tri   n5124;
  tri   n5125;
  tri   n5126;
  tri   n5127;
  tri   n5128;
  tri   n5129;
  tri   n5013;
  tri   n5014;
  tri   n5016;
  tri   n5017;
  tri   P1_N5582;
  tri   n5020;
  tri   n5021;
  tri   n5022;
  tri   n5023;
  tri   n5024;
  tri   n5025;
  tri   n5026;
  tri   n5027;
  tri   n5028;
  tri   n5029;
  tri   n5030;
  tri   n5031;
  tri   n5032;
  tri   n5033;
  tri   n5034;
  tri   n5035;
  tri   n5036;
  tri   n5037;
  tri   n5038;
  tri   n5039;
  tri   n5040;
  tri   n5041;
  tri   n5042;
  tri   n5043;
  tri   n5044;
  tri   n5045;
  tri   n5046;
  tri   n5047;
  tri   n5048;
  tri   n5049;
  tri   n5050;
  tri   n5051;
  tri   n5052;
  tri   n5053;
  tri   n5054;
  tri   n5055;
  tri   n5056;
  tri   n5057;
  tri   n5058;
  tri   n5059;
  tri   n5060;
  tri   n5061;
  tri   n5062;
  tri   n5063;
  tri   n5064;
  tri   n5065;
  tri   n5066;
  tri   n5067;
  tri   n5068;
  tri   n5069;
  tri   n5070;
  tri   n5071;
  tri   n5072;
  tri   n5073;
  tri   n5074;
  tri   n5075;
  tri   n4963;
  tri   P1_N5583;
  tri   n4962;
  tri   n4964;
  tri   n4965;
  tri   n4966;
  tri   n4967;
  tri   n4968;
  tri   n4969;
  tri   n4970;
  tri   n4971;
  tri   n4972;
  tri   n4973;
  tri   n4974;
  tri   n4975;
  tri   n4976;
  tri   n4977;
  tri   n4978;
  tri   n4979;
  tri   n4980;
  tri   n4981;
  tri   n4982;
  tri   n4983;
  tri   n4984;
  tri   n4985;
  tri   n4986;
  tri   n4987;
  tri   n4988;
  tri   n4989;
  tri   n4992;
  tri   n4993;
  tri   n4995;
  tri   n4996;
  tri   n4997;
  tri   n4998;
  tri   n4999;
  tri   n5000;
  tri   n5001;
  tri   n5002;
  tri   n5003;
  tri   n5004;
  tri   n5005;
  tri   n5006;
  tri   n5007;
  tri   n5008;
  tri   n5009;
  tri   n5010;
  tri   n5011;
  tri   n5012;
  tri   n4909;
  tri   n4910;
  tri   n4911;
  tri   n4912;
  tri   n4913;
  tri   n4914;
  tri   n4915;
  tri   n4916;
  tri   n4917;
  tri   n4918;
  tri   n4919;
  tri   n4920;
  tri   n4921;
  tri   n4922;
  tri   n4923;
  tri   n4924;
  tri   n4925;
  tri   n4926;
  tri   n4927;
  tri   n4928;
  tri   n4930;
  tri   n4931;
  tri   n4934;
  tri   n4935;
  tri   n4936;
  tri   n4937;
  tri   n4938;
  tri   n4939;
  tri   n4940;
  tri   n4941;
  tri   n4942;
  tri   n4943;
  tri   n4944;
  tri   n4945;
  tri   n4946;
  tri   n4947;
  tri   n4948;
  tri   n4949;
  tri   n4950;
  tri   n4951;
  tri   n4952;
  tri   n4953;
  tri   n4954;
  tri   n4955;
  tri   n4956;
  tri   n4957;
  tri   n4958;
  tri   n4959;
  tri   n4960;
  tri   n4961;
  tri   n4847;
  tri   n4848;
  tri   n4840;
  tri   n4849;
  tri   n4850;
  tri   P1_N411;
  tri   P1_N410;
  tri   P1_N409;
  tri   P1_N408;
  tri   P1_N405;
  tri   n4851;
  tri   P1_N406;
  tri   P1_N407;
  tri   n4852;
  tri   n4853;
  tri   P1_N5584;
  tri   n4854;
  tri   n4855;
  tri   n4856;
  tri   n4857;
  tri   n4858;
  tri   n4859;
  tri   n4860;
  tri   n4861;
  tri   n4862;
  tri   n4863;
  tri   n4864;
  tri   n4865;
  tri   n4866;
  tri   n4867;
  tri   n4868;
  tri   n4869;
  tri   n4870;
  tri   n4871;
  tri   n4872;
  tri   n4873;
  tri   n4874;
  tri   n4875;
  tri   n4876;
  tri   n4877;
  tri   n4878;
  tri   n4879;
  tri   n4880;
  tri   n4881;
  tri   n4882;
  tri   n4883;
  tri   n4884;
  tri   n4885;
  tri   n4886;
  tri   n4887;
  tri   n4888;
  tri   n4889;
  tri   n4890;
  tri   n4891;
  tri   n4892;
  tri   n4893;
  tri   n4894;
  tri   n4895;
  tri   n4896;
  tri   n4897;
  tri   n4898;
  tri   n4899;
  tri   n4900;
  tri   n4901;
  tri   n4902;
  tri   n4903;
  tri   n4906;
  tri   n4907;
  tri   n4772;
  tri   n4771;
  tri   n4773;
  tri   n4774;
  tri   n4775;
  tri   n4776;
  tri   n4777;
  tri   n4778;
  tri   n4584;
  tri   P1_N5571;
  tri   n4780;
  tri   n4779;
  tri   n4781;
  tri   n4782;
  tri   n4783;
  tri   n4784;
  tri   n4785;
  tri   n4786;
  tri   n4788;
  tri   n4787;
  tri   n4789;
  tri   n4790;
  tri   n4791;
  tri   n4792;
  tri   n4793;
  tri   n4794;
  tri   n4796;
  tri   n4795;
  tri   n4797;
  tri   n4798;
  tri   n4799;
  tri   n4800;
  tri   n4801;
  tri   n4802;
  tri   n4806;
  tri   n4807;
  tri   n4808;
  tri   n4809;
  tri   n4811;
  tri   n4812;
  tri   n4813;
  tri   n4816;
  tri   n4817;
  tri   n4820;
  tri   n4821;
  tri   n4822;
  tri   n4823;
  tri   P1_N395;
  tri   n4824;
  tri   n4825;
  tri   n4826;
  tri   n4827;
  tri   n4828;
  tri   n4829;
  tri   n4830;
  tri   n4831;
  tri   n4832;
  tri   P1_N418;
  tri   P1_N417;
  tri   P1_N416;
  tri   P1_N415;
  tri   P1_N412;
  tri   n4833;
  tri   P1_N413;
  tri   P1_N414;
  tri   n4835;
  tri   n4834;
  tri   n4836;
  tri   n4837;
  tri   P1_N422;
  tri   P1_N421;
  tri   P1_N420;
  tri   P1_N419;
  tri   n4838;
  tri   n4839;
  tri   P1_N426;
  tri   P1_N425;
  tri   P1_N424;
  tri   P1_N423;
  tri   n4841;
  tri   n4842;
  tri   n4843;
  tri   n4844;
  tri   n4845;
  tri   P1_N404;
  tri   P1_N403;
  tri   P1_N402;
  tri   P1_N401;
  tri   P1_N398;
  tri   n4846;
  tri   P1_N399;
  tri   P1_N400;
  tri   n4697;
  tri   n4698;
  tri   n4700;
  tri   n4699;
  tri   n4701;
  tri   n4702;
  tri   n4703;
  tri   n4704;
  tri   n4705;
  tri   n4706;
  tri   n4708;
  tri   n4707;
  tri   n4709;
  tri   n4710;
  tri   n4711;
  tri   n4712;
  tri   n4713;
  tri   n4714;
  tri   n4716;
  tri   n4715;
  tri   n4717;
  tri   n4718;
  tri   n4719;
  tri   n4720;
  tri   n4721;
  tri   n4722;
  tri   n4724;
  tri   n4723;
  tri   n4725;
  tri   n4726;
  tri   n4727;
  tri   n4728;
  tri   n4729;
  tri   n4730;
  tri   n4732;
  tri   n4731;
  tri   n4733;
  tri   n4734;
  tri   n4735;
  tri   n4736;
  tri   n4737;
  tri   n4738;
  tri   n4740;
  tri   n4739;
  tri   n4741;
  tri   n4742;
  tri   n4743;
  tri   n4744;
  tri   n4745;
  tri   n4746;
  tri   n4748;
  tri   n4747;
  tri   n4749;
  tri   n4750;
  tri   n4751;
  tri   n4752;
  tri   n4753;
  tri   n4754;
  tri   n4756;
  tri   n4755;
  tri   n4757;
  tri   n4758;
  tri   n4759;
  tri   n4760;
  tri   n4761;
  tri   n4762;
  tri   n4764;
  tri   n4763;
  tri   n4765;
  tri   n4766;
  tri   n4767;
  tri   n4768;
  tri   n4769;
  tri   n4770;
  tri   n4623;
  tri   n4624;
  tri   n4619;
  tri   n4625;
  tri   n4626;
  tri   n4628;
  tri   n4627;
  tri   n4629;
  tri   n4630;
  tri   n4631;
  tri   n4632;
  tri   n4633;
  tri   n4634;
  tri   n4636;
  tri   n4635;
  tri   n4637;
  tri   n4638;
  tri   n4639;
  tri   n4640;
  tri   n4641;
  tri   n4642;
  tri   n4644;
  tri   n4643;
  tri   n4645;
  tri   n4646;
  tri   n4647;
  tri   n4648;
  tri   n4649;
  tri   n4650;
  tri   n4652;
  tri   n4651;
  tri   n4653;
  tri   n4654;
  tri   n4655;
  tri   n4656;
  tri   n4657;
  tri   n4658;
  tri   n4660;
  tri   n4659;
  tri   n4661;
  tri   n4662;
  tri   n4663;
  tri   n4664;
  tri   n4665;
  tri   n4666;
  tri   n4668;
  tri   n4667;
  tri   n4669;
  tri   n4670;
  tri   n4671;
  tri   n4672;
  tri   n4673;
  tri   n4674;
  tri   n4676;
  tri   n4675;
  tri   n4677;
  tri   n4678;
  tri   n4679;
  tri   n4680;
  tri   n4681;
  tri   n4682;
  tri   n4684;
  tri   n4683;
  tri   n4685;
  tri   n4686;
  tri   n4687;
  tri   n4688;
  tri   n4689;
  tri   n4690;
  tri   n4692;
  tri   n4691;
  tri   n4693;
  tri   n4694;
  tri   n4695;
  tri   n4696;
  tri   n4551;
  tri   P1_N5574;
  tri   n4550;
  tri   n4552;
  tri   n4553;
  tri   n4554;
  tri   n4555;
  tri   n4556;
  tri   n4557;
  tri   n4558;
  tri   n4559;
  tri   n4560;
  tri   n4561;
  tri   n4562;
  tri   n4563;
  tri   n4564;
  tri   n4565;
  tri   n4566;
  tri   n4567;
  tri   n4570;
  tri   n4571;
  tri   n4572;
  tri   n4573;
  tri   n4574;
  tri   n4506;
  tri   n4575;
  tri   n4577;
  tri   n4576;
  tri   n4578;
  tri   n4579;
  tri   n4580;
  tri   n4581;
  tri   n4582;
  tri   n4583;
  tri   n4586;
  tri   n4585;
  tri   n4587;
  tri   n4588;
  tri   n4589;
  tri   n4590;
  tri   n4591;
  tri   n4592;
  tri   n4594;
  tri   n4593;
  tri   n4595;
  tri   n4596;
  tri   n4597;
  tri   n4598;
  tri   n4599;
  tri   n4600;
  tri   n4602;
  tri   n4601;
  tri   n4603;
  tri   n4604;
  tri   n4605;
  tri   n4606;
  tri   n4607;
  tri   n4608;
  tri   n4610;
  tri   n4609;
  tri   n4611;
  tri   n4612;
  tri   n4613;
  tri   n4614;
  tri   n4617;
  tri   n4618;
  tri   n4620;
  tri   n4621;
  tri   n4622;
  tri   n4483;
  tri   n4484;
  tri   n4482;
  tri   n4485;
  tri   n4486;
  tri   n4481;
  tri   P1_N543;
  tri   n4492;
  tri   n4493;
  tri   n4084;
  tri   n4494;
  tri   n4175;
  tri   n4495;
  tri   n4496;
  tri   n4497;
  tri   P1_N542;
  tri   P1_N541;
  tri   n4500;
  tri   n4501;
  tri   n4086;
  tri   n4502;
  tri   n4503;
  tri   n4178;
  tri   n4504;
  tri   n4505;
  tri   n4508;
  tri   n4509;
  tri   n4512;
  tri   n4513;
  tri   n4514;
  tri   n4515;
  tri   n4516;
  tri   n4517;
  tri   n4518;
  tri   n4519;
  tri   n4520;
  tri   n4521;
  tri   n4522;
  tri   n4523;
  tri   n4524;
  tri   n4525;
  tri   n4526;
  tri   n4527;
  tri   n4528;
  tri   n4529;
  tri   n4530;
  tri   n4531;
  tri   n4532;
  tri   n4533;
  tri   n4534;
  tri   n4535;
  tri   n4536;
  tri   n4537;
  tri   n4538;
  tri   n4539;
  tri   n4540;
  tri   n4541;
  tri   n4542;
  tri   n4543;
  tri   n4544;
  tri   n4545;
  tri   n4546;
  tri   n4547;
  tri   n4548;
  tri   n4549;
  tri   n4429;
  tri   n4431;
  tri   n4432;
  tri   n4433;
  tri   n4434;
  tri   n4435;
  tri   n4436;
  tri   n4437;
  tri   n4438;
  tri   n4439;
  tri   n4440;
  tri   n4441;
  tri   n4442;
  tri   n4443;
  tri   n4444;
  tri   n4445;
  tri   n4446;
  tri   n4447;
  tri   n4448;
  tri   n4449;
  tri   n4450;
  tri   n4451;
  tri   n4452;
  tri   n4453;
  tri   n4454;
  tri   n4455;
  tri   n4456;
  tri   n4457;
  tri   n4458;
  tri   n4459;
  tri   n4460;
  tri   n4461;
  tri   n4462;
  tri   n4463;
  tri   n4464;
  tri   n4465;
  tri   n4466;
  tri   n4467;
  tri   n4468;
  tri   n4470;
  tri   n4471;
  tri   P1_N4977;
  tri   P1_N4971;
  tri   n4472;
  tri   n4473;
  tri   P1_N5570;
  tri   P1_N4970;
  tri   n4475;
  tri   n4476;
  tri   n4477;
  tri   n4363;
  tri   n4359;
  tri   n4360;
  tri   n4370;
  tri   n4371;
  tri   P1_N531;
  tri   n4372;
  tri   P1_N530;
  tri   n4373;
  tri   n4374;
  tri   n4377;
  tri   n4378;
  tri   n4379;
  tri   n4380;
  tri   n4381;
  tri   n4382;
  tri   n4383;
  tri   n4384;
  tri   n4385;
  tri   n4387;
  tri   n4388;
  tri   n4389;
  tri   n4390;
  tri   n4391;
  tri   n4392;
  tri   n4393;
  tri   n4394;
  tri   n4395;
  tri   n4396;
  tri   n4397;
  tri   n4398;
  tri   n4399;
  tri   n4400;
  tri   n4401;
  tri   n4402;
  tri   n4403;
  tri   n4404;
  tri   n4405;
  tri   n4406;
  tri   n4407;
  tri   n4408;
  tri   n4409;
  tri   n4410;
  tri   n4411;
  tri   n4412;
  tri   n4413;
  tri   n4414;
  tri   n4415;
  tri   n4416;
  tri   n4417;
  tri   n4418;
  tri   n4419;
  tri   n4420;
  tri   n4421;
  tri   n4422;
  tri   n4423;
  tri   n4424;
  tri   n4425;
  tri   n4426;
  tri   n4427;
  tri   n4428;
  tri   n4430;
  tri   n4272;
  tri   P1_N5513;
  tri   n4273;
  tri   n4274;
  tri   n4277;
  tri   P1_N5512;
  tri   n4278;
  tri   n4279;
  tri   n4282;
  tri   P1_N5511;
  tri   n4283;
  tri   n4284;
  tri   n4287;
  tri   P1_N5510;
  tri   n4288;
  tri   n4289;
  tri   n4292;
  tri   P1_N5509;
  tri   n4293;
  tri   n4294;
  tri   n4297;
  tri   P1_N5508;
  tri   n4298;
  tri   n4299;
  tri   n4302;
  tri   P1_N5507;
  tri   n4303;
  tri   n4304;
  tri   n4307;
  tri   P1_N5506;
  tri   n4308;
  tri   n4309;
  tri   n4312;
  tri   P1_N5505;
  tri   n4313;
  tri   n4314;
  tri   n4317;
  tri   P1_N5504;
  tri   n4318;
  tri   n4319;
  tri   n4323;
  tri   P1_N5503;
  tri   n4324;
  tri   n4325;
  tri   n4329;
  tri   n4328;
  tri   P1_N5502;
  tri   n4330;
  tri   n4331;
  tri   n4332;
  tri   n4333;
  tri   n4172;
  tri   n4335;
  tri   P1_N5501;
  tri   n4336;
  tri   n4337;
  tri   n4341;
  tri   n4340;
  tri   P1_N5500;
  tri   n4342;
  tri   n4343;
  tri   n4344;
  tri   n4345;
  tri   n4347;
  tri   P1_N5499;
  tri   n4348;
  tri   n4349;
  tri   n4353;
  tri   P1_N5498;
  tri   n4354;
  tri   n4355;
  tri   n4361;
  tri   P1_N5518;
  tri   n4362;
  tri   n4364;
  tri   n4198;
  tri   n4197;
  tri   n4200;
  tri   n4201;
  tri   P1_N5543;
  tri   n4203;
  tri   n4204;
  tri   P1_N5542;
  tri   n4206;
  tri   n4207;
  tri   P1_N5541;
  tri   n4209;
  tri   n4210;
  tri   P1_N5540;
  tri   n4211;
  tri   n4212;
  tri   P1_N5539;
  tri   n4213;
  tri   n4214;
  tri   P1_N5538;
  tri   n4215;
  tri   n4216;
  tri   P1_N5537;
  tri   n4217;
  tri   n4218;
  tri   P1_N5536;
  tri   n4219;
  tri   n4220;
  tri   P1_N5535;
  tri   n4221;
  tri   n4222;
  tri   P1_N5534;
  tri   n4223;
  tri   n4224;
  tri   P1_N5532;
  tri   n4225;
  tri   n4226;
  tri   P1_N5531;
  tri   n4227;
  tri   n4228;
  tri   P1_N5530;
  tri   n4229;
  tri   n4230;
  tri   P1_N5529;
  tri   n4231;
  tri   n4232;
  tri   P1_N5528;
  tri   n4233;
  tri   n4234;
  tri   P1_N5527;
  tri   n4235;
  tri   n4236;
  tri   P1_N5526;
  tri   n4237;
  tri   n4238;
  tri   P1_N5525;
  tri   n4239;
  tri   n4240;
  tri   P1_N5524;
  tri   n4241;
  tri   n4242;
  tri   P1_N5523;
  tri   n4243;
  tri   n4244;
  tri   P1_N5522;
  tri   n4245;
  tri   n4246;
  tri   P1_N5521;
  tri   n4247;
  tri   n4248;
  tri   P1_N5520;
  tri   n4251;
  tri   P1_N5517;
  tri   n4252;
  tri   n4253;
  tri   n4257;
  tri   P1_N5516;
  tri   n4258;
  tri   n4259;
  tri   n4262;
  tri   P1_N5515;
  tri   n4263;
  tri   n4264;
  tri   n4267;
  tri   P1_N5514;
  tri   n4268;
  tri   n4269;
  tri   n4098;
  tri   n4101;
  tri   n4104;
  tri   n4107;
  tri   n4110;
  tri   n4113;
  tri   n4116;
  tri   n4119;
  tri   n4122;
  tri   n4125;
  tri   n4128;
  tri   n4131;
  tri   n4134;
  tri   n4137;
  tri   n4140;
  tri   n4143;
  tri   n4146;
  tri   n4149;
  tri   n4152;
  tri   n4155;
  tri   n4166;
  tri   P1_N5561;
  tri   n4167;
  tri   n4168;
  tri   P1_N5560;
  tri   n4173;
  tri   n4174;
  tri   P1_N5553;
  tri   n4176;
  tri   n4177;
  tri   P1_N5552;
  tri   n4179;
  tri   n4180;
  tri   P1_N5551;
  tri   n4182;
  tri   n4183;
  tri   P1_N5550;
  tri   n4185;
  tri   n4186;
  tri   P1_N5549;
  tri   n4188;
  tri   n4189;
  tri   P1_N5547;
  tri   n4191;
  tri   n4192;
  tri   P1_N5546;
  tri   n4194;
  tri   n4195;
  tri   P1_N5545;
  tri   P1_N5544;
  tri   n4020;
  tri   n4021;
  tri   P1_N5576;
  tri   n4024;
  tri   n4025;
  tri   n4026;
  tri   n4027;
  tri   n4028;
  tri   n4029;
  tri   n4030;
  tri   n4031;
  tri   n4032;
  tri   n4033;
  tri   n4034;
  tri   n4035;
  tri   n4036;
  tri   n4037;
  tri   n4038;
  tri   n4039;
  tri   n4040;
  tri   n4041;
  tri   n4042;
  tri   n4043;
  tri   n4044;
  tri   n4045;
  tri   n4046;
  tri   n4047;
  tri   n4048;
  tri   n4049;
  tri   n4050;
  tri   n4051;
  tri   n4052;
  tri   n4053;
  tri   n4054;
  tri   n4055;
  tri   n4056;
  tri   n4057;
  tri   n4058;
  tri   n4059;
  tri   n4060;
  tri   n4061;
  tri   n4062;
  tri   n4063;
  tri   n4064;
  tri   n4065;
  tri   n4066;
  tri   n4067;
  tri   n4068;
  tri   n4069;
  tri   n4070;
  tri   n4071;
  tri   n4072;
  tri   n4073;
  tri   n4074;
  tri   n4075;
  tri   n4076;
  tri   n4077;
  tri   n4078;
  tri   n4079;
  tri   n4082;
  tri   n4083;
  tri   n3957;
  tri   n3958;
  tri   n3955;
  tri   n3959;
  tri   n3960;
  tri   n3961;
  tri   n3962;
  tri   n3965;
  tri   n3966;
  tri   n3967;
  tri   n3968;
  tri   n3969;
  tri   n3970;
  tri   n3971;
  tri   n3972;
  tri   n3973;
  tri   n3974;
  tri   n3975;
  tri   n3976;
  tri   n3977;
  tri   n3978;
  tri   n3979;
  tri   n3980;
  tri   n3981;
  tri   n3982;
  tri   n3983;
  tri   n3984;
  tri   n3985;
  tri   n3986;
  tri   n3987;
  tri   n3988;
  tri   n3989;
  tri   n3990;
  tri   n3991;
  tri   n3992;
  tri   n3993;
  tri   n3994;
  tri   n3995;
  tri   n3996;
  tri   n3997;
  tri   n3998;
  tri   n3999;
  tri   n4000;
  tri   n4001;
  tri   n4002;
  tri   n4003;
  tri   n4004;
  tri   n4005;
  tri   n4006;
  tri   n4007;
  tri   n4008;
  tri   n4009;
  tri   n4010;
  tri   n4011;
  tri   n4012;
  tri   n4013;
  tri   n4014;
  tri   n4015;
  tri   n4016;
  tri   n4017;
  tri   n4018;
  tri   n2048;
  tri   P2_N5495;
  tri   n3893;
  tri   n3898;
  tri   n3899;
  tri   n2051;
  tri   n3900;
  tri   n2053;
  tri   n3901;
  tri   n3902;
  tri   n3903;
  tri   n3904;
  tri   n2054;
  tri   n3905;
  tri   n2056;
  tri   n3906;
  tri   n3907;
  tri   n3908;
  tri   n3909;
  tri   n2057;
  tri   n3910;
  tri   n2059;
  tri   n3911;
  tri   n3912;
  tri   n3913;
  tri   n3914;
  tri   n2060;
  tri   n3915;
  tri   n2062;
  tri   n3916;
  tri   n3917;
  tri   n3918;
  tri   n3919;
  tri   n2063;
  tri   n3920;
  tri   n2065;
  tri   n3921;
  tri   n3922;
  tri   n3925;
  tri   n3926;
  tri   n3927;
  tri   n3928;
  tri   n3929;
  tri   n3930;
  tri   n3931;
  tri   n3932;
  tri   n3933;
  tri   n3934;
  tri   n3935;
  tri   n3936;
  tri   n3937;
  tri   n3938;
  tri   n3939;
  tri   n3940;
  tri   n3941;
  tri   n3942;
  tri   n3943;
  tri   n3944;
  tri   n3945;
  tri   n3946;
  tri   n3949;
  tri   n3950;
  tri   n3953;
  tri   n3954;
  tri   n3956;
  tri   n2018;
  tri   n3843;
  tri   n3848;
  tri   n3849;
  tri   n2021;
  tri   n3850;
  tri   n3853;
  tri   n3854;
  tri   n3855;
  tri   n3858;
  tri   n3859;
  tri   n3860;
  tri   n3863;
  tri   n3864;
  tri   n3865;
  tri   n2032;
  tri   n3866;
  tri   n3867;
  tri   n3868;
  tri   n3869;
  tri   n2033;
  tri   n3870;
  tri   n2035;
  tri   n3871;
  tri   n3872;
  tri   n3873;
  tri   n3874;
  tri   n2036;
  tri   n3875;
  tri   n2038;
  tri   n3876;
  tri   n3877;
  tri   n3878;
  tri   n3879;
  tri   n2039;
  tri   n3880;
  tri   n3883;
  tri   n3884;
  tri   n2042;
  tri   n3885;
  tri   n3888;
  tri   n3889;
  tri   n2045;
  tri   n3890;
  tri   n2047;
  tri   n3891;
  tri   n3892;
  tri   n3894;
  tri   n3895;
  tri   n2050;
  tri   n3896;
  tri   n3897;
  tri   n3790;
  tri   n3791;
  tri   n3792;
  tri   n3794;
  tri   n3795;
  tri   n3798;
  tri   n3799;
  tri   n3800;
  tri   n3801;
  tri   n3802;
  tri   n3803;
  tri   n3804;
  tri   n3805;
  tri   n3806;
  tri   n3807;
  tri   n3809;
  tri   n3810;
  tri   n3811;
  tri   n3812;
  tri   n3813;
  tri   n3814;
  tri   n3815;
  tri   n3816;
  tri   n3817;
  tri   n3818;
  tri   n3819;
  tri   n3820;
  tri   n3821;
  tri   n3822;
  tri   n3823;
  tri   n3824;
  tri   n2006;
  tri   n3825;
  tri   n3828;
  tri   n3829;
  tri   n2009;
  tri   n3830;
  tri   n3833;
  tri   n3834;
  tri   n2012;
  tri   n3835;
  tri   n3838;
  tri   n3839;
  tri   n2015;
  tri   n3840;
  tri   n3844;
  tri   n3845;
  tri   P2_N5496;
  tri   n3738;
  tri   n3740;
  tri   n3741;
  tri   n3742;
  tri   n3743;
  tri   n3744;
  tri   n3745;
  tri   n3746;
  tri   n3747;
  tri   n3748;
  tri   n3749;
  tri   n3750;
  tri   n3751;
  tri   n3752;
  tri   n3753;
  tri   n3754;
  tri   n3755;
  tri   n3756;
  tri   n3757;
  tri   n3758;
  tri   n3759;
  tri   n3760;
  tri   n3761;
  tri   n3762;
  tri   n3763;
  tri   n3764;
  tri   n3765;
  tri   n3766;
  tri   n3767;
  tri   n3770;
  tri   n3771;
  tri   n3773;
  tri   n3774;
  tri   n3775;
  tri   n3776;
  tri   n3777;
  tri   n3778;
  tri   n3779;
  tri   n3780;
  tri   n3781;
  tri   n3782;
  tri   n3783;
  tri   n3784;
  tri   n3785;
  tri   n3786;
  tri   n3787;
  tri   n3788;
  tri   n3789;
  tri   n3687;
  tri   n3688;
  tri   n3689;
  tri   n3690;
  tri   n3691;
  tri   n3692;
  tri   n3693;
  tri   n3694;
  tri   n3695;
  tri   n3696;
  tri   n3697;
  tri   n3698;
  tri   n3699;
  tri   n3700;
  tri   n3701;
  tri   n3702;
  tri   n3703;
  tri   n3704;
  tri   n3705;
  tri   n3706;
  tri   n3708;
  tri   n3709;
  tri   n3712;
  tri   n3713;
  tri   n3714;
  tri   n3715;
  tri   n3716;
  tri   n3717;
  tri   n3718;
  tri   n3719;
  tri   n3720;
  tri   n3721;
  tri   n3722;
  tri   n3723;
  tri   n3724;
  tri   n3725;
  tri   n3726;
  tri   n3727;
  tri   n3728;
  tri   n3729;
  tri   n3730;
  tri   n3731;
  tri   n3732;
  tri   n3733;
  tri   n3734;
  tri   n3735;
  tri   n3736;
  tri   n3737;
  tri   n3739;
  tri   n3623;
  tri   P2_N5502;
  tri   n3622;
  tri   n3626;
  tri   n3627;
  tri   n3628;
  tri   n3629;
  tri   n3630;
  tri   n3631;
  tri   n3632;
  tri   n3633;
  tri   n3634;
  tri   n3635;
  tri   n3636;
  tri   n3637;
  tri   n3638;
  tri   n3639;
  tri   n3640;
  tri   n3641;
  tri   n3642;
  tri   n3643;
  tri   n3644;
  tri   n3645;
  tri   n3646;
  tri   n3647;
  tri   n3648;
  tri   n3649;
  tri   n3650;
  tri   n3651;
  tri   n3652;
  tri   n3653;
  tri   n3654;
  tri   n3655;
  tri   n3656;
  tri   n3657;
  tri   n3658;
  tri   n3659;
  tri   n3660;
  tri   n3661;
  tri   n3662;
  tri   n3663;
  tri   n3664;
  tri   n3665;
  tri   n3666;
  tri   n3667;
  tri   n3668;
  tri   n3669;
  tri   n3670;
  tri   n3671;
  tri   n3672;
  tri   n3673;
  tri   n3674;
  tri   n3675;
  tri   n3676;
  tri   n3677;
  tri   n3678;
  tri   n3679;
  tri   n3680;
  tri   n3681;
  tri   n3684;
  tri   n3685;
  tri   n3564;
  tri   n3565;
  tri   P2_N5503;
  tri   n3566;
  tri   n3567;
  tri   n3568;
  tri   n3569;
  tri   n3572;
  tri   n3573;
  tri   P2_N134;
  tri   n3574;
  tri   n3575;
  tri   n3576;
  tri   n3577;
  tri   n3578;
  tri   n3579;
  tri   n3580;
  tri   n3581;
  tri   n3582;
  tri   P2_N156;
  tri   P2_N155;
  tri   P2_N154;
  tri   P2_N153;
  tri   P2_N150;
  tri   n3583;
  tri   P2_N151;
  tri   P2_N152;
  tri   n3584;
  tri   n3585;
  tri   n3586;
  tri   n3587;
  tri   P2_N163;
  tri   P2_N162;
  tri   P2_N161;
  tri   P2_N160;
  tri   P2_N157;
  tri   n3588;
  tri   P2_N158;
  tri   P2_N159;
  tri   n3589;
  tri   n3590;
  tri   n3591;
  tri   n3592;
  tri   P2_N140;
  tri   n3593;
  tri   P2_N141;
  tri   P2_N142;
  tri   P2_N137;
  tri   n3594;
  tri   P2_N138;
  tri   P2_N139;
  tri   n3595;
  tri   n3596;
  tri   n3597;
  tri   n3598;
  tri   P2_N149;
  tri   P2_N148;
  tri   P2_N147;
  tri   P2_N146;
  tri   P2_N143;
  tri   n3599;
  tri   P2_N144;
  tri   P2_N145;
  tri   n3601;
  tri   n3602;
  tri   n3603;
  tri   n3604;
  tri   n3605;
  tri   n3606;
  tri   n3607;
  tri   n3608;
  tri   n3609;
  tri   n3610;
  tri   n3611;
  tri   n3612;
  tri   n3613;
  tri   n3614;
  tri   n3615;
  tri   n3616;
  tri   n3617;
  tri   n3618;
  tri   n3619;
  tri   n3620;
  tri   n3501;
  tri   n3502;
  tri   n3503;
  tri   n3504;
  tri   n3505;
  tri   n3506;
  tri   n3507;
  tri   n3508;
  tri   n3510;
  tri   n3511;
  tri   n3514;
  tri   n3515;
  tri   n3516;
  tri   n3517;
  tri   n3518;
  tri   n3519;
  tri   n3520;
  tri   n3521;
  tri   n3522;
  tri   n3523;
  tri   n3524;
  tri   n3525;
  tri   n3526;
  tri   n3527;
  tri   n3528;
  tri   n3529;
  tri   n3530;
  tri   n3531;
  tri   n3532;
  tri   n3533;
  tri   n3534;
  tri   n3535;
  tri   n3536;
  tri   n3537;
  tri   n3538;
  tri   n3539;
  tri   n3540;
  tri   n3541;
  tri   n3542;
  tri   n3543;
  tri   n3544;
  tri   n3545;
  tri   n3546;
  tri   n3547;
  tri   n3548;
  tri   n3549;
  tri   n3550;
  tri   n3551;
  tri   n3552;
  tri   n3553;
  tri   n3554;
  tri   n3555;
  tri   n3556;
  tri   n3557;
  tri   n3558;
  tri   n3559;
  tri   n3560;
  tri   n3561;
  tri   n3562;
  tri   n3563;
  tri   P2_N5504;
  tri   n3441;
  tri   n3443;
  tri   n3444;
  tri   n3445;
  tri   n3446;
  tri   n3447;
  tri   n3448;
  tri   n3449;
  tri   n3450;
  tri   n3451;
  tri   n3452;
  tri   n3453;
  tri   n3454;
  tri   n3455;
  tri   n3456;
  tri   n3457;
  tri   n3458;
  tri   n3459;
  tri   n3460;
  tri   P2_N193;
  tri   n3463;
  tri   n3464;
  tri   n3465;
  tri   n3466;
  tri   n3467;
  tri   n3468;
  tri   n3469;
  tri   P2_N212;
  tri   n3470;
  tri   P2_N213;
  tri   P2_N214;
  tri   P2_N209;
  tri   n3471;
  tri   P2_N210;
  tri   P2_N211;
  tri   n3472;
  tri   n3473;
  tri   P2_N218;
  tri   n3474;
  tri   P2_N219;
  tri   P2_N220;
  tri   P2_N215;
  tri   n3475;
  tri   P2_N216;
  tri   P2_N217;
  tri   n3476;
  tri   n3477;
  tri   n3478;
  tri   n3479;
  tri   P2_N200;
  tri   n3480;
  tri   P2_N201;
  tri   P2_N202;
  tri   P2_N197;
  tri   n3481;
  tri   P2_N198;
  tri   P2_N199;
  tri   n3482;
  tri   n3483;
  tri   P2_N206;
  tri   n3484;
  tri   P2_N207;
  tri   P2_N208;
  tri   P2_N203;
  tri   n3485;
  tri   P2_N204;
  tri   P2_N205;
  tri   n3486;
  tri   n3487;
  tri   n3489;
  tri   n3490;
  tri   n3491;
  tri   n3492;
  tri   n3493;
  tri   n3494;
  tri   n3495;
  tri   n3496;
  tri   n3497;
  tri   n3498;
  tri   n3499;
  tri   n3500;
  tri   n3383;
  tri   n3384;
  tri   n3385;
  tri   n3386;
  tri   n3387;
  tri   n3388;
  tri   n3389;
  tri   n3390;
  tri   n3391;
  tri   n3392;
  tri   n3393;
  tri   n3394;
  tri   n3395;
  tri   n3396;
  tri   n3397;
  tri   n3398;
  tri   n3399;
  tri   n3401;
  tri   n3402;
  tri   n3405;
  tri   n3406;
  tri   n3407;
  tri   n3408;
  tri   n3409;
  tri   n3410;
  tri   n3411;
  tri   n3412;
  tri   n3413;
  tri   n3414;
  tri   n3415;
  tri   n3416;
  tri   n3417;
  tri   n3418;
  tri   n3419;
  tri   n3420;
  tri   n3421;
  tri   n3422;
  tri   n3423;
  tri   n3424;
  tri   n3425;
  tri   n3426;
  tri   n3427;
  tri   n3428;
  tri   n3429;
  tri   n3430;
  tri   n3431;
  tri   n3432;
  tri   n3433;
  tri   n3434;
  tri   n3435;
  tri   n3436;
  tri   n3437;
  tri   n3438;
  tri   n3439;
  tri   n3440;
  tri   n3442;
  tri   P2_N5505;
  tri   n3321;
  tri   n3323;
  tri   n3324;
  tri   n3325;
  tri   n3326;
  tri   n3327;
  tri   n3328;
  tri   n3329;
  tri   n3330;
  tri   n3331;
  tri   n3332;
  tri   n3333;
  tri   n3334;
  tri   n3335;
  tri   n3336;
  tri   n3337;
  tri   n3338;
  tri   n3339;
  tri   n3340;
  tri   n3341;
  tri   n3342;
  tri   n3343;
  tri   n3344;
  tri   n3345;
  tri   n3346;
  tri   n3347;
  tri   n3348;
  tri   n3349;
  tri   n3350;
  tri   n3351;
  tri   n3352;
  tri   n3353;
  tri   n3354;
  tri   n3355;
  tri   n3356;
  tri   P2_N248;
  tri   n3359;
  tri   n3360;
  tri   n3361;
  tri   n3362;
  tri   n3363;
  tri   n3364;
  tri   n3365;
  tri   P2_N264;
  tri   n3366;
  tri   P2_N265;
  tri   P2_N266;
  tri   P2_N263;
  tri   P2_N262;
  tri   n3367;
  tri   n3368;
  tri   P2_N269;
  tri   n3369;
  tri   P2_N270;
  tri   P2_N271;
  tri   P2_N268;
  tri   P2_N267;
  tri   n3370;
  tri   n3371;
  tri   n3372;
  tri   n3373;
  tri   P2_N256;
  tri   P2_N255;
  tri   P2_N254;
  tri   P2_N253;
  tri   n3374;
  tri   n3375;
  tri   P2_N259;
  tri   n3376;
  tri   P2_N260;
  tri   P2_N261;
  tri   P2_N258;
  tri   P2_N257;
  tri   n3377;
  tri   n3378;
  tri   n3380;
  tri   n3381;
  tri   n3382;
  tri   n3270;
  tri   P2_N5506;
  tri   n3269;
  tri   n3273;
  tri   n3274;
  tri   n3276;
  tri   n3277;
  tri   n3278;
  tri   n3279;
  tri   n3280;
  tri   n3281;
  tri   n3282;
  tri   n3283;
  tri   n3284;
  tri   n3285;
  tri   n3286;
  tri   n3287;
  tri   n3288;
  tri   n3289;
  tri   n3290;
  tri   n3291;
  tri   n3292;
  tri   n3293;
  tri   n3294;
  tri   n3295;
  tri   n3297;
  tri   n3298;
  tri   n3301;
  tri   n3302;
  tri   n3303;
  tri   n3304;
  tri   n3305;
  tri   n3306;
  tri   n3307;
  tri   n3308;
  tri   n3309;
  tri   n3310;
  tri   n3311;
  tri   n3312;
  tri   n3313;
  tri   n3314;
  tri   n3315;
  tri   n3316;
  tri   n3317;
  tri   n3318;
  tri   n3319;
  tri   n3320;
  tri   n3322;
  tri   n3206;
  tri   n3207;
  tri   n3208;
  tri   n3209;
  tri   n3211;
  tri   n3212;
  tri   n3215;
  tri   n3216;
  tri   n3217;
  tri   n3218;
  tri   n3219;
  tri   n3220;
  tri   n3221;
  tri   n3222;
  tri   n3223;
  tri   n3224;
  tri   n3225;
  tri   n3226;
  tri   n3227;
  tri   n3228;
  tri   n3229;
  tri   n3230;
  tri   n3231;
  tri   n3232;
  tri   n3233;
  tri   n3234;
  tri   n3235;
  tri   n3236;
  tri   n3237;
  tri   n3238;
  tri   n3239;
  tri   n3240;
  tri   n3241;
  tri   n3242;
  tri   n3243;
  tri   n3244;
  tri   n3245;
  tri   n3246;
  tri   n3247;
  tri   n3248;
  tri   n3249;
  tri   n3250;
  tri   n3251;
  tri   n3252;
  tri   n3253;
  tri   n3254;
  tri   n3255;
  tri   n3256;
  tri   n3257;
  tri   n3258;
  tri   n3259;
  tri   n3260;
  tri   n3261;
  tri   n3262;
  tri   n3263;
  tri   n3264;
  tri   n3265;
  tri   n3266;
  tri   n3267;
  tri   n3268;
  tri   P2_N5507;
  tri   n3147;
  tri   n3149;
  tri   n3150;
  tri   n3151;
  tri   n3152;
  tri   n3153;
  tri   n3154;
  tri   n3155;
  tri   n3156;
  tri   n3157;
  tri   n3158;
  tri   n3159;
  tri   n3160;
  tri   n3161;
  tri   n3162;
  tri   n3165;
  tri   n3166;
  tri   P2_N295;
  tri   n3167;
  tri   P2_N342;
  tri   n3168;
  tri   n3169;
  tri   n3170;
  tri   n3171;
  tri   n3172;
  tri   n3173;
  tri   P2_N311;
  tri   n3174;
  tri   P2_N312;
  tri   P2_N313;
  tri   P2_N308;
  tri   n3175;
  tri   P2_N309;
  tri   P2_N310;
  tri   n3176;
  tri   n3177;
  tri   P2_N317;
  tri   n3178;
  tri   P2_N318;
  tri   P2_N319;
  tri   P2_N314;
  tri   n3179;
  tri   P2_N315;
  tri   P2_N316;
  tri   n3180;
  tri   n3181;
  tri   n3182;
  tri   n3183;
  tri   P2_N299;
  tri   n3184;
  tri   P2_N300;
  tri   P2_N301;
  tri   P2_N298;
  tri   P2_N297;
  tri   n3185;
  tri   n3186;
  tri   P2_N305;
  tri   n3187;
  tri   P2_N306;
  tri   P2_N307;
  tri   P2_N302;
  tri   n3188;
  tri   P2_N303;
  tri   P2_N304;
  tri   n3190;
  tri   n3191;
  tri   n3192;
  tri   n3193;
  tri   n3194;
  tri   n3195;
  tri   n3196;
  tri   n3197;
  tri   n3198;
  tri   n3199;
  tri   n3200;
  tri   n3201;
  tri   n3202;
  tri   n3203;
  tri   n3204;
  tri   n3205;
  tri   n3088;
  tri   n3089;
  tri   n3090;
  tri   n3091;
  tri   n3092;
  tri   n3093;
  tri   n3094;
  tri   n3095;
  tri   n3096;
  tri   n3097;
  tri   n3098;
  tri   n3099;
  tri   n3100;
  tri   n3101;
  tri   n3103;
  tri   n3104;
  tri   n3107;
  tri   n3108;
  tri   n3109;
  tri   n3110;
  tri   n3111;
  tri   n3112;
  tri   n3113;
  tri   n3114;
  tri   n3115;
  tri   n3116;
  tri   n3117;
  tri   n3118;
  tri   n3119;
  tri   n3120;
  tri   n3121;
  tri   n3122;
  tri   n3123;
  tri   n3124;
  tri   n3125;
  tri   n3126;
  tri   n3127;
  tri   n3128;
  tri   n3129;
  tri   n3130;
  tri   n3131;
  tri   n3132;
  tri   n3133;
  tri   n3134;
  tri   n3135;
  tri   n3136;
  tri   n3137;
  tri   n3138;
  tri   n3139;
  tri   n3140;
  tri   n3141;
  tri   n3142;
  tri   n3143;
  tri   n3144;
  tri   n3145;
  tri   n3146;
  tri   n3148;
  tri   n3034;
  tri   P2_N5508;
  tri   n3033;
  tri   n3035;
  tri   n3036;
  tri   n3037;
  tri   n3038;
  tri   n3039;
  tri   n3040;
  tri   n3041;
  tri   n3042;
  tri   n3043;
  tri   n3044;
  tri   n3045;
  tri   n3046;
  tri   n3047;
  tri   n3048;
  tri   n3049;
  tri   n3050;
  tri   n3051;
  tri   n3052;
  tri   n3053;
  tri   n3054;
  tri   n3055;
  tri   n3056;
  tri   n3057;
  tri   n3058;
  tri   n3059;
  tri   n3060;
  tri   n3061;
  tri   n3062;
  tri   n3063;
  tri   n3064;
  tri   n3065;
  tri   n3066;
  tri   n3067;
  tri   n3068;
  tri   n3069;
  tri   n3070;
  tri   n3071;
  tri   n3072;
  tri   n3073;
  tri   n3074;
  tri   n3075;
  tri   n3076;
  tri   n3079;
  tri   n3080;
  tri   n3082;
  tri   n3083;
  tri   n3084;
  tri   n3085;
  tri   n3086;
  tri   n3087;
  tri   n2980;
  tri   n2982;
  tri   n2983;
  tri   n2984;
  tri   n2985;
  tri   n2986;
  tri   n2987;
  tri   n2988;
  tri   n2989;
  tri   n2990;
  tri   n2991;
  tri   n2996;
  tri   n2997;
  tri   n2998;
  tri   n2999;
  tri   n3000;
  tri   n3001;
  tri   n3002;
  tri   n3003;
  tri   n3004;
  tri   n3005;
  tri   n3006;
  tri   n3007;
  tri   n3008;
  tri   n3009;
  tri   n3010;
  tri   n3011;
  tri   n3012;
  tri   n3013;
  tri   n3014;
  tri   n3015;
  tri   n3017;
  tri   n3018;
  tri   n3021;
  tri   n3022;
  tri   n3023;
  tri   n3024;
  tri   n3025;
  tri   n3026;
  tri   n3027;
  tri   n3028;
  tri   n3029;
  tri   n3030;
  tri   n3031;
  tri   n3032;
  tri   P2_N5493;
  tri   n2917;
  tri   n2702;
  tri   n2922;
  tri   n2923;
  tri   n2924;
  tri   n2925;
  tri   n2926;
  tri   n2927;
  tri   n2928;
  tri   n2929;
  tri   n2567;
  tri   n2930;
  tri   n2932;
  tri   n2933;
  tri   n2936;
  tri   n2937;
  tri   n2938;
  tri   n2939;
  tri   n2940;
  tri   n2941;
  tri   n2942;
  tri   n2943;
  tri   n2944;
  tri   n2945;
  tri   n2946;
  tri   n2947;
  tri   n2948;
  tri   n2949;
  tri   n2950;
  tri   n2951;
  tri   n2952;
  tri   n2953;
  tri   n2954;
  tri   n2955;
  tri   n2956;
  tri   n2957;
  tri   n2958;
  tri   n2959;
  tri   n2960;
  tri   n2961;
  tri   n2962;
  tri   n2963;
  tri   n2964;
  tri   n2965;
  tri   n2966;
  tri   n2967;
  tri   n2968;
  tri   n2969;
  tri   n2970;
  tri   n2971;
  tri   n2972;
  tri   n2973;
  tri   n2974;
  tri   n2975;
  tri   n2976;
  tri   n2977;
  tri   n2978;
  tri   n2979;
  tri   n2981;
  tri   n2843;
  tri   n2845;
  tri   n2846;
  tri   n2848;
  tri   n2847;
  tri   n2849;
  tri   n2850;
  tri   n2851;
  tri   n2852;
  tri   n2853;
  tri   n2854;
  tri   n2856;
  tri   n2855;
  tri   n2857;
  tri   n2858;
  tri   n2859;
  tri   n2860;
  tri   n2861;
  tri   n2862;
  tri   n2864;
  tri   n2863;
  tri   n2865;
  tri   n2866;
  tri   n2867;
  tri   n2868;
  tri   n2869;
  tri   n2870;
  tri   n2872;
  tri   n2871;
  tri   n2873;
  tri   n2874;
  tri   n2875;
  tri   n2876;
  tri   n2877;
  tri   n2878;
  tri   n2880;
  tri   n2879;
  tri   n2881;
  tri   n2882;
  tri   n2883;
  tri   n2884;
  tri   n2885;
  tri   n2886;
  tri   n2888;
  tri   n2887;
  tri   n2889;
  tri   n2890;
  tri   n2891;
  tri   n2892;
  tri   n2893;
  tri   n2894;
  tri   n2896;
  tri   n2895;
  tri   n2897;
  tri   n2898;
  tri   n2899;
  tri   n2900;
  tri   n2901;
  tri   n2902;
  tri   n2904;
  tri   n2903;
  tri   n2905;
  tri   n2906;
  tri   n2907;
  tri   n2908;
  tri   n2909;
  tri   n2910;
  tri   n2912;
  tri   n2911;
  tri   n2913;
  tri   n2914;
  tri   n2915;
  tri   n2916;
  tri   n2918;
  tri   n2769;
  tri   n2771;
  tri   n2772;
  tri   n2767;
  tri   n2773;
  tri   n2774;
  tri   n2776;
  tri   n2775;
  tri   n2777;
  tri   n2778;
  tri   n2779;
  tri   n2780;
  tri   n2781;
  tri   n2782;
  tri   n2784;
  tri   n2783;
  tri   n2785;
  tri   n2786;
  tri   n2787;
  tri   n2788;
  tri   n2789;
  tri   n2790;
  tri   n2792;
  tri   n2791;
  tri   n2793;
  tri   n2794;
  tri   n2795;
  tri   n2796;
  tri   n2797;
  tri   n2798;
  tri   n2800;
  tri   n2799;
  tri   n2801;
  tri   n2802;
  tri   n2803;
  tri   n2804;
  tri   n2805;
  tri   n2806;
  tri   n2808;
  tri   n2807;
  tri   n2809;
  tri   n2810;
  tri   n2811;
  tri   n2812;
  tri   n2813;
  tri   n2814;
  tri   n2816;
  tri   n2815;
  tri   n2817;
  tri   n2818;
  tri   n2819;
  tri   n2820;
  tri   n2821;
  tri   n2822;
  tri   n2824;
  tri   n2823;
  tri   n2825;
  tri   n2826;
  tri   n2827;
  tri   n2828;
  tri   n2829;
  tri   n2830;
  tri   n2832;
  tri   n2831;
  tri   n2833;
  tri   n2834;
  tri   n2835;
  tri   n2836;
  tri   n2837;
  tri   n2838;
  tri   n2840;
  tri   n2839;
  tri   n2841;
  tri   n2842;
  tri   n2844;
  tri   n2695;
  tri   n2694;
  tri   n2696;
  tri   n2697;
  tri   n2698;
  tri   n2699;
  tri   n2700;
  tri   n2701;
  tri   n2704;
  tri   n2703;
  tri   n2705;
  tri   n2706;
  tri   n2707;
  tri   n2708;
  tri   n2709;
  tri   n2710;
  tri   n2712;
  tri   n2711;
  tri   n2713;
  tri   n2714;
  tri   n2715;
  tri   n2716;
  tri   n2717;
  tri   n2718;
  tri   n2720;
  tri   n2719;
  tri   n2721;
  tri   n2722;
  tri   n2723;
  tri   n2724;
  tri   n2725;
  tri   n2726;
  tri   n2728;
  tri   n2727;
  tri   n2729;
  tri   n2730;
  tri   n2731;
  tri   n2732;
  tri   n2733;
  tri   n2734;
  tri   n2736;
  tri   n2735;
  tri   n2737;
  tri   n2738;
  tri   n2739;
  tri   n2740;
  tri   n2741;
  tri   n2742;
  tri   n2744;
  tri   n2743;
  tri   n2745;
  tri   n2746;
  tri   n2747;
  tri   n2748;
  tri   n2749;
  tri   n2750;
  tri   n2752;
  tri   n2751;
  tri   n2753;
  tri   n2754;
  tri   n2755;
  tri   n2756;
  tri   n2757;
  tri   n2758;
  tri   n2760;
  tri   n2759;
  tri   n2761;
  tri   n2762;
  tri   n2763;
  tri   n2764;
  tri   n2765;
  tri   n2766;
  tri   n2768;
  tri   n2770;
  tri   n2599;
  tri   n2624;
  tri   n2623;
  tri   n2625;
  tri   n2626;
  tri   n2627;
  tri   n2628;
  tri   n2629;
  tri   n2630;
  tri   n2631;
  tri   n2632;
  tri   n2633;
  tri   n2634;
  tri   n2635;
  tri   n2636;
  tri   n2637;
  tri   n2638;
  tri   n2639;
  tri   n2640;
  tri   n2641;
  tri   n2642;
  tri   n2643;
  tri   n2644;
  tri   n2645;
  tri   n2646;
  tri   n2647;
  tri   n2648;
  tri   n2649;
  tri   n2650;
  tri   n2651;
  tri   n2652;
  tri   n2653;
  tri   n2654;
  tri   n2655;
  tri   n2656;
  tri   P2_N395;
  tri   n2662;
  tri   n2663;
  tri   n2664;
  tri   n2665;
  tri   n2666;
  tri   n2667;
  tri   n2668;
  tri   n2669;
  tri   n2670;
  tri   P2_N418;
  tri   P2_N417;
  tri   P2_N416;
  tri   P2_N415;
  tri   P2_N412;
  tri   n2671;
  tri   P2_N413;
  tri   P2_N414;
  tri   n2673;
  tri   n2672;
  tri   n2674;
  tri   n2675;
  tri   P2_N422;
  tri   P2_N421;
  tri   P2_N420;
  tri   P2_N419;
  tri   n2676;
  tri   n2677;
  tri   P2_N426;
  tri   P2_N425;
  tri   P2_N424;
  tri   P2_N423;
  tri   n2678;
  tri   n2679;
  tri   n2680;
  tri   n2681;
  tri   n2682;
  tri   n2683;
  tri   P2_N404;
  tri   P2_N403;
  tri   P2_N402;
  tri   P2_N401;
  tri   P2_N398;
  tri   n2684;
  tri   P2_N399;
  tri   P2_N400;
  tri   n2685;
  tri   n2686;
  tri   n2687;
  tri   n2688;
  tri   P2_N411;
  tri   P2_N410;
  tri   P2_N409;
  tri   P2_N408;
  tri   P2_N405;
  tri   n2689;
  tri   P2_N406;
  tri   P2_N407;
  tri   n2690;
  tri   n2691;
  tri   n2589;
  tri   n2692;
  tri   n2554;
  tri   n2555;
  tri   n2556;
  tri   n2557;
  tri   n2558;
  tri   n2559;
  tri   n2560;
  tri   n2561;
  tri   n2564;
  tri   n2563;
  tri   n2565;
  tri   n2566;
  tri   n2568;
  tri   n2571;
  tri   n2570;
  tri   n2572;
  tri   n2573;
  tri   n2574;
  tri   n2575;
  tri   n2576;
  tri   P2_N4809;
  tri   P2_N4808;
  tri   n2581;
  tri   n2582;
  tri   n2172;
  tri   n2583;
  tri   n2584;
  tri   n2588;
  tri   n2175;
  tri   n2590;
  tri   n2591;
  tri   n2592;
  tri   n2593;
  tri   n2594;
  tri   n2595;
  tri   P2_N543;
  tri   P2_N542;
  tri   P2_N541;
  tri   n2597;
  tri   n2598;
  tri   n2601;
  tri   n2602;
  tri   n2603;
  tri   n2604;
  tri   n2605;
  tri   n2606;
  tri   n2607;
  tri   n2608;
  tri   n2609;
  tri   n2610;
  tri   n2611;
  tri   n2612;
  tri   n2613;
  tri   n2614;
  tri   n2615;
  tri   n2616;
  tri   n2617;
  tri   n2618;
  tri   n2619;
  tri   n2620;
  tri   n2621;
  tri   n2622;
  tri   n2505;
  tri   n2504;
  tri   n2506;
  tri   n2507;
  tri   n2508;
  tri   n2509;
  tri   n2510;
  tri   n2511;
  tri   n2512;
  tri   n2513;
  tri   n2514;
  tri   n2515;
  tri   n2516;
  tri   n2517;
  tri   n2518;
  tri   n2519;
  tri   n2520;
  tri   n2521;
  tri   n2522;
  tri   n2523;
  tri   n2524;
  tri   n2525;
  tri   n2526;
  tri   n2527;
  tri   n2528;
  tri   n2529;
  tri   n2530;
  tri   n2531;
  tri   n2532;
  tri   n2533;
  tri   n2534;
  tri   n2535;
  tri   n2536;
  tri   n2537;
  tri   n2538;
  tri   n2539;
  tri   n2540;
  tri   n2541;
  tri   n2542;
  tri   n2543;
  tri   n2544;
  tri   n2545;
  tri   n2546;
  tri   n2547;
  tri   n2548;
  tri   n2549;
  tri   n2550;
  tri   n2551;
  tri   n2552;
  tri   n2553;
  tri   n2252;
  tri   n2434;
  tri   n2253;
  tri   n2433;
  tri   n2254;
  tri   n2431;
  tri   n2429;
  tri   n2435;
  tri   n2436;
  tri   n2437;
  tri   n2438;
  tri   n2161;
  tri   n2439;
  tri   n2440;
  tri   P2_N5420;
  tri   n2441;
  tri   n2442;
  tri   n2443;
  tri   n2444;
  tri   n2445;
  tri   P2_N5492;
  tri   n2169;
  tri   n2447;
  tri   n2448;
  tri   n2449;
  tri   n2450;
  tri   n2451;
  tri   n2453;
  tri   n2454;
  tri   P2_N5440;
  tri   n2455;
  tri   n2456;
  tri   n2457;
  tri   n2463;
  tri   n2464;
  tri   P2_N531;
  tri   n2465;
  tri   P2_N530;
  tri   n2466;
  tri   n2467;
  tri   n2470;
  tri   n2471;
  tri   n2472;
  tri   n2473;
  tri   n2474;
  tri   n2475;
  tri   n2476;
  tri   n2477;
  tri   n2478;
  tri   n2480;
  tri   n2481;
  tri   n2482;
  tri   n2483;
  tri   n2484;
  tri   n2485;
  tri   n2486;
  tri   n2487;
  tri   n2488;
  tri   n2489;
  tri   n2490;
  tri   n2491;
  tri   n2492;
  tri   n2493;
  tri   n2494;
  tri   n2495;
  tri   n2496;
  tri   n2497;
  tri   n2498;
  tri   n2499;
  tri   n2500;
  tri   n2501;
  tri   n2502;
  tri   n2503;
  tri   n2347;
  tri   n2345;
  tri   n2349;
  tri   n2350;
  tri   P2_N5429;
  tri   n2351;
  tri   n2352;
  tri   n2353;
  tri   n2354;
  tri   n2355;
  tri   n2356;
  tri   n2357;
  tri   n2358;
  tri   n2359;
  tri   n2360;
  tri   P2_N5428;
  tri   n2361;
  tri   n2362;
  tri   n2363;
  tri   n2364;
  tri   n2365;
  tri   n2366;
  tri   n2367;
  tri   n2368;
  tri   n2369;
  tri   n2370;
  tri   P2_N5427;
  tri   n2371;
  tri   n2372;
  tri   n2373;
  tri   n2374;
  tri   n2375;
  tri   n2376;
  tri   n2377;
  tri   n2378;
  tri   n2379;
  tri   n2380;
  tri   P2_N5426;
  tri   n2381;
  tri   n2382;
  tri   n2383;
  tri   n2384;
  tri   n2385;
  tri   n2386;
  tri   n2387;
  tri   n2388;
  tri   n2389;
  tri   n2390;
  tri   P2_N5425;
  tri   n2391;
  tri   n2392;
  tri   n2393;
  tri   n2394;
  tri   n2395;
  tri   n2396;
  tri   n2397;
  tri   n2398;
  tri   n2399;
  tri   n2400;
  tri   P2_N5424;
  tri   n2401;
  tri   n2402;
  tri   n2403;
  tri   n2404;
  tri   n2405;
  tri   n2406;
  tri   n2407;
  tri   n2408;
  tri   n2409;
  tri   n2410;
  tri   P2_N5423;
  tri   n2411;
  tri   n2412;
  tri   n2413;
  tri   n2414;
  tri   n2415;
  tri   n2416;
  tri   n2417;
  tri   n2418;
  tri   n2419;
  tri   n2420;
  tri   P2_N5422;
  tri   n2421;
  tri   n2422;
  tri   n2423;
  tri   n2424;
  tri   n2425;
  tri   n2426;
  tri   n2427;
  tri   n2428;
  tri   n2430;
  tri   P2_N5421;
  tri   n2432;
  tri   n2263;
  tri   n2261;
  tri   n2259;
  tri   n2265;
  tri   n2266;
  tri   n2267;
  tri   n2268;
  tri   n2269;
  tri   n2270;
  tri   P2_N5437;
  tri   n2271;
  tri   n2272;
  tri   n2273;
  tri   n2274;
  tri   n2275;
  tri   n2276;
  tri   n2277;
  tri   n2278;
  tri   n2279;
  tri   n2280;
  tri   P2_N5436;
  tri   n2281;
  tri   n2282;
  tri   n2283;
  tri   n2284;
  tri   n2285;
  tri   n2286;
  tri   n2287;
  tri   n2288;
  tri   n2289;
  tri   n2290;
  tri   P2_N5435;
  tri   n2291;
  tri   n2292;
  tri   n2293;
  tri   n2294;
  tri   n2295;
  tri   n2296;
  tri   n2297;
  tri   n2298;
  tri   n2299;
  tri   n2300;
  tri   P2_N5434;
  tri   n2301;
  tri   n2302;
  tri   n2303;
  tri   n2304;
  tri   n2305;
  tri   n2306;
  tri   n2307;
  tri   n2308;
  tri   n2309;
  tri   n2310;
  tri   P2_N5433;
  tri   n2311;
  tri   n2312;
  tri   n2313;
  tri   n2314;
  tri   n2315;
  tri   n2316;
  tri   n2317;
  tri   n2318;
  tri   n2319;
  tri   n2320;
  tri   P2_N5432;
  tri   n2321;
  tri   n2322;
  tri   n2323;
  tri   n2324;
  tri   n2325;
  tri   n2326;
  tri   n2327;
  tri   n2328;
  tri   n2329;
  tri   n2330;
  tri   P2_N5431;
  tri   n2331;
  tri   n2332;
  tri   n2333;
  tri   n2334;
  tri   n2335;
  tri   n2336;
  tri   n2337;
  tri   n2338;
  tri   n2339;
  tri   n2340;
  tri   P2_N5430;
  tri   n2341;
  tri   n2342;
  tri   n2343;
  tri   n2344;
  tri   n2346;
  tri   n2348;
  tri   n2192;
  tri   n2191;
  tri   n2194;
  tri   n2195;
  tri   P2_N5466;
  tri   n2197;
  tri   n2198;
  tri   P2_N5465;
  tri   n2200;
  tri   n2201;
  tri   P2_N5464;
  tri   n2203;
  tri   n2204;
  tri   P2_N5463;
  tri   n2206;
  tri   n2207;
  tri   P2_N5462;
  tri   n2208;
  tri   n2209;
  tri   P2_N5461;
  tri   n2210;
  tri   n2211;
  tri   P2_N5460;
  tri   n2212;
  tri   n2213;
  tri   P2_N5459;
  tri   n2214;
  tri   n2215;
  tri   P2_N5458;
  tri   n2216;
  tri   n2217;
  tri   P2_N5457;
  tri   n2218;
  tri   n2219;
  tri   P2_N5456;
  tri   n2220;
  tri   n2221;
  tri   P2_N5454;
  tri   n2222;
  tri   n2223;
  tri   P2_N5453;
  tri   n2224;
  tri   n2225;
  tri   P2_N5452;
  tri   n2226;
  tri   n2227;
  tri   P2_N5451;
  tri   n2228;
  tri   n2229;
  tri   P2_N5450;
  tri   n2230;
  tri   n2231;
  tri   P2_N5449;
  tri   n2232;
  tri   n2233;
  tri   P2_N5448;
  tri   n2234;
  tri   n2235;
  tri   P2_N5447;
  tri   n2236;
  tri   n2237;
  tri   P2_N5446;
  tri   n2238;
  tri   n2239;
  tri   P2_N5445;
  tri   n2240;
  tri   n2241;
  tri   P2_N5444;
  tri   n2242;
  tri   n2243;
  tri   P2_N5443;
  tri   n2244;
  tri   n2245;
  tri   P2_N5442;
  tri   n2246;
  tri   n2247;
  tri   P2_N5439;
  tri   n2248;
  tri   n2249;
  tri   n2250;
  tri   n2251;
  tri   n2255;
  tri   n2256;
  tri   n2257;
  tri   n2258;
  tri   n2260;
  tri   P2_N5438;
  tri   n2262;
  tri   n2264;
  tri   n2130;
  tri   n2133;
  tri   n2134;
  tri   n2135;
  tri   n2136;
  tri   n2137;
  tri   n2138;
  tri   n2139;
  tri   n2140;
  tri   n2141;
  tri   n2142;
  tri   n2143;
  tri   n2144;
  tri   n2145;
  tri   n2146;
  tri   n2147;
  tri   n2148;
  tri   n2149;
  tri   n2150;
  tri   n2151;
  tri   n2152;
  tri   n2163;
  tri   P2_N5483;
  tri   n2164;
  tri   n2165;
  tri   P2_N5482;
  tri   n2170;
  tri   n2171;
  tri   P2_N5475;
  tri   n2173;
  tri   n2174;
  tri   P2_N5474;
  tri   n2176;
  tri   n2177;
  tri   P2_N5473;
  tri   n2179;
  tri   n2180;
  tri   P2_N5472;
  tri   n2182;
  tri   n2183;
  tri   P2_N5471;
  tri   n2185;
  tri   n2186;
  tri   P2_N5469;
  tri   n2188;
  tri   n2189;
  tri   P2_N5468;
  tri   P2_N5467;
  tri   n2064;
  tri   n2067;
  tri   n2068;
  tri   P2_N5494;
  tri   n2071;
  tri   n2072;
  tri   n2073;
  tri   n2074;
  tri   n2075;
  tri   n2076;
  tri   n2077;
  tri   n2078;
  tri   n2079;
  tri   n2080;
  tri   n2081;
  tri   n2082;
  tri   n2083;
  tri   n2084;
  tri   n2085;
  tri   n2086;
  tri   n2087;
  tri   n2088;
  tri   n2089;
  tri   n2090;
  tri   n2091;
  tri   n2092;
  tri   n2093;
  tri   n2094;
  tri   n2095;
  tri   n2096;
  tri   n2097;
  tri   n2098;
  tri   n2099;
  tri   n2100;
  tri   n2101;
  tri   n2102;
  tri   n2103;
  tri   n2104;
  tri   n2105;
  tri   n2106;
  tri   n2107;
  tri   n2108;
  tri   n2109;
  tri   n2110;
  tri   n2111;
  tri   n2112;
  tri   n2113;
  tri   n2114;
  tri   n2115;
  tri   n2116;
  tri   n2117;
  tri   n2118;
  tri   n2119;
  tri   n2120;
  tri   n2121;
  tri   n2122;
  tri   n2123;
  tri   n2124;
  tri   n2125;
  tri   n2126;
  tri   n2129;
  tri   n1478;
  tri   n1482;
  tri   n1483;
  tri   n1484;
  tri   n1486;
  tri   n1487;
  tri   n1488;
  tri   n1489;
  tri   n1490;
  tri   n1491;
  tri   n1492;
  tri   n1493;
  tri   n1494;
  tri   n1495;
  tri   n1497;
  tri   n1498;
  tri   n1500;
  tri   n1501;
  tri   n2007;
  tri   n2010;
  tri   n2013;
  tri   n2016;
  tri   n2019;
  tri   n2022;
  tri   n2025;
  tri   n2028;
  tri   n2031;
  tri   n2034;
  tri   n2037;
  tri   n2040;
  tri   n2043;
  tri   n2046;
  tri   n2049;
  tri   n2052;
  tri   n2055;
  tri   n2058;
  tri   n2061;
  tri   n1423;
  tri   n1422;
  tri   n1424;
  tri   n1425;
  tri   n6298;
  tri   n1426;
  tri   n1427;
  tri   n6299;
  tri   n1428;
  tri   n1429;
  tri   n6300;
  tri   n1430;
  tri   n1431;
  tri   n6301;
  tri   n1432;
  tri   n1433;
  tri   n6302;
  tri   n1434;
  tri   n1435;
  tri   n6303;
  tri   n1436;
  tri   n1437;
  tri   n6304;
  tri   n1438;
  tri   n1439;
  tri   n6305;
  tri   n1440;
  tri   n1441;
  tri   n6306;
  tri   n1442;
  tri   n1443;
  tri   n6307;
  tri   n1444;
  tri   n1445;
  tri   n6308;
  tri   n1446;
  tri   n1447;
  tri   n6309;
  tri   n1448;
  tri   n1449;
  tri   n6310;
  tri   n1450;
  tri   n1451;
  tri   n6311;
  tri   n1452;
  tri   n1453;
  tri   n6312;
  tri   n1454;
  tri   n1455;
  tri   n6313;
  tri   n1456;
  tri   n1457;
  tri   n6314;
  tri   n1458;
  tri   n1459;
  tri   n6315;
  tri   n1460;
  tri   n1461;
  tri   n6316;
  tri   n1462;
  tri   n1463;
  tri   n6317;
  tri   n1464;
  tri   n1465;
  tri   n6318;
  tri   n1467;
  tri   n1468;
  tri   n1469;
  tri   n1470;
  tri   n1471;
  tri   n1472;
  tri   n1473;
  tri   n1475;
  tri   n1476;
  tri   n1477;
  tri   n1479;
  tri   n1360;
  tri   n1362;
  tri   n1363;
  tri   n6267;
  tri   n1364;
  tri   n1365;
  tri   n6268;
  tri   n1366;
  tri   n1367;
  tri   n6269;
  tri   n1368;
  tri   n1369;
  tri   n6270;
  tri   n1370;
  tri   n1371;
  tri   n6271;
  tri   n1372;
  tri   n1373;
  tri   n6272;
  tri   n1374;
  tri   n1375;
  tri   n6273;
  tri   n1376;
  tri   n1377;
  tri   n6274;
  tri   n1378;
  tri   n1379;
  tri   n6275;
  tri   n1380;
  tri   n1381;
  tri   n6276;
  tri   n1382;
  tri   n1383;
  tri   n6277;
  tri   n1384;
  tri   n1385;
  tri   n6278;
  tri   n1386;
  tri   n1387;
  tri   n6279;
  tri   n1388;
  tri   n1389;
  tri   n6280;
  tri   n1390;
  tri   n1391;
  tri   n6281;
  tri   n1392;
  tri   n1393;
  tri   n6282;
  tri   n1394;
  tri   n1395;
  tri   n6283;
  tri   n1396;
  tri   n1397;
  tri   n6284;
  tri   n1398;
  tri   n1399;
  tri   n6285;
  tri   n1400;
  tri   n1401;
  tri   n6286;
  tri   n1402;
  tri   n1403;
  tri   n6287;
  tri   n1404;
  tri   n1405;
  tri   n6288;
  tri   n1406;
  tri   n1407;
  tri   n6289;
  tri   n1408;
  tri   n1409;
  tri   n6290;
  tri   n1410;
  tri   n1411;
  tri   n6291;
  tri   n1412;
  tri   n1413;
  tri   n6292;
  tri   n1414;
  tri   n1415;
  tri   n6293;
  tri   n1416;
  tri   n1417;
  tri   n6294;
  tri   n1418;
  tri   n1419;
  tri   n6295;
  tri   n1420;
  tri   n1421;
  tri   n6296;
  tri   n6297;
  tri   n1300;
  tri   n1301;
  tri   n6236;
  tri   n1302;
  tri   n1303;
  tri   n6237;
  tri   n1304;
  tri   n1305;
  tri   n6238;
  tri   n1306;
  tri   n1307;
  tri   n6239;
  tri   n1308;
  tri   n1309;
  tri   n6240;
  tri   n1310;
  tri   n1311;
  tri   n6241;
  tri   n1312;
  tri   n1313;
  tri   n6242;
  tri   n1314;
  tri   n1315;
  tri   n6243;
  tri   n1316;
  tri   n1317;
  tri   n6244;
  tri   n1318;
  tri   n1319;
  tri   n6245;
  tri   n1320;
  tri   n1321;
  tri   n6246;
  tri   n1322;
  tri   n1323;
  tri   n6247;
  tri   n1324;
  tri   n1325;
  tri   n6248;
  tri   n1326;
  tri   n1327;
  tri   n6249;
  tri   n1328;
  tri   n1329;
  tri   n6250;
  tri   n1330;
  tri   n1331;
  tri   n6251;
  tri   n1332;
  tri   n1333;
  tri   n6252;
  tri   n1334;
  tri   n1335;
  tri   n6253;
  tri   n1336;
  tri   n1337;
  tri   n6254;
  tri   n1338;
  tri   n1339;
  tri   n6255;
  tri   n1340;
  tri   n1341;
  tri   n6256;
  tri   n1342;
  tri   n1343;
  tri   n6257;
  tri   n1344;
  tri   n1345;
  tri   n6258;
  tri   n1346;
  tri   n1347;
  tri   n6259;
  tri   n1348;
  tri   n1349;
  tri   n6260;
  tri   n1350;
  tri   n1351;
  tri   n6261;
  tri   n1352;
  tri   n1353;
  tri   n6262;
  tri   n1354;
  tri   n1355;
  tri   n6263;
  tri   n1356;
  tri   n1357;
  tri   n6264;
  tri   n1358;
  tri   n1359;
  tri   n6265;
  tri   n1361;
  tri   n6266;
  tri   n1239;
  tri   n1238;
  tri   n1240;
  tri   n1241;
  tri   n6206;
  tri   n1242;
  tri   n1243;
  tri   n6207;
  tri   n1244;
  tri   n1245;
  tri   n6208;
  tri   n1246;
  tri   n1247;
  tri   n6209;
  tri   n1248;
  tri   n1249;
  tri   n6210;
  tri   n1250;
  tri   n1251;
  tri   n6211;
  tri   n1252;
  tri   n1253;
  tri   n6212;
  tri   n1254;
  tri   n1255;
  tri   n6213;
  tri   n1256;
  tri   n1257;
  tri   n6214;
  tri   n1258;
  tri   n1259;
  tri   n6215;
  tri   n1260;
  tri   n1261;
  tri   n6216;
  tri   n1262;
  tri   n1263;
  tri   n6217;
  tri   n1264;
  tri   n1265;
  tri   n6218;
  tri   n1266;
  tri   n1267;
  tri   n6219;
  tri   n1268;
  tri   n1269;
  tri   n6220;
  tri   n1270;
  tri   n1271;
  tri   n6221;
  tri   n1272;
  tri   n1273;
  tri   n6222;
  tri   n1274;
  tri   n1275;
  tri   n6223;
  tri   n1276;
  tri   n1277;
  tri   n6224;
  tri   n1278;
  tri   n1279;
  tri   n6225;
  tri   n1280;
  tri   n1281;
  tri   n6226;
  tri   n1282;
  tri   n1283;
  tri   n6227;
  tri   n1284;
  tri   n1285;
  tri   n6228;
  tri   n1286;
  tri   n1287;
  tri   n6229;
  tri   n1288;
  tri   n1289;
  tri   n6230;
  tri   n1290;
  tri   n1291;
  tri   n6231;
  tri   n1292;
  tri   n1293;
  tri   n6232;
  tri   n1294;
  tri   n1295;
  tri   n6233;
  tri   n1296;
  tri   n1297;
  tri   n6234;
  tri   n1298;
  tri   n1299;
  tri   n6235;
  tri   n1176;
  tri   n1177;
  tri   n6175;
  tri   n1178;
  tri   n1179;
  tri   n6176;
  tri   n1180;
  tri   n1181;
  tri   n6177;
  tri   n1183;
  tri   n1184;
  tri   n6178;
  tri   n1186;
  tri   n1187;
  tri   n6179;
  tri   n1188;
  tri   n1189;
  tri   n6180;
  tri   n1190;
  tri   n1191;
  tri   n6181;
  tri   n1192;
  tri   n1193;
  tri   n6182;
  tri   n1194;
  tri   n1195;
  tri   n6183;
  tri   n1196;
  tri   n1197;
  tri   n6184;
  tri   n1198;
  tri   n1199;
  tri   n6185;
  tri   n1200;
  tri   n1201;
  tri   n6186;
  tri   n1202;
  tri   n1203;
  tri   n6187;
  tri   n1204;
  tri   n1205;
  tri   n6188;
  tri   n1206;
  tri   n1207;
  tri   n6189;
  tri   n1208;
  tri   n1209;
  tri   n6190;
  tri   n1210;
  tri   n1211;
  tri   n6191;
  tri   n1212;
  tri   n1213;
  tri   n6192;
  tri   n1214;
  tri   n1215;
  tri   n6193;
  tri   n1216;
  tri   n1217;
  tri   n6194;
  tri   n1218;
  tri   n1219;
  tri   n6195;
  tri   n1220;
  tri   n1221;
  tri   n6196;
  tri   n1222;
  tri   n1223;
  tri   n6197;
  tri   n1224;
  tri   n1225;
  tri   n6198;
  tri   n1226;
  tri   n1227;
  tri   n6199;
  tri   n1228;
  tri   n1229;
  tri   n6200;
  tri   n1230;
  tri   n1231;
  tri   n6201;
  tri   n1232;
  tri   n1233;
  tri   n6202;
  tri   n1234;
  tri   n1235;
  tri   n6203;
  tri   n1236;
  tri   n1237;
  tri   n6204;
  tri   n6205;
  tri   n1112;
  tri   n1114;
  tri   n1115;
  tri   n6145;
  tri   n1116;
  tri   n1117;
  tri   n1118;
  tri   n6146;
  tri   n1119;
  tri   n1120;
  tri   n6147;
  tri   n1121;
  tri   n1122;
  tri   n1123;
  tri   n6148;
  tri   n1124;
  tri   n1125;
  tri   n6149;
  tri   n1126;
  tri   n1127;
  tri   n6150;
  tri   n1128;
  tri   n1129;
  tri   n6151;
  tri   n1130;
  tri   n1131;
  tri   n6152;
  tri   n1132;
  tri   n1133;
  tri   n6153;
  tri   n1134;
  tri   n1135;
  tri   n6154;
  tri   n1136;
  tri   n1137;
  tri   n6155;
  tri   n1138;
  tri   n1139;
  tri   n6156;
  tri   n1140;
  tri   n1141;
  tri   n6157;
  tri   n1142;
  tri   n1143;
  tri   n6158;
  tri   n1144;
  tri   n1145;
  tri   n6159;
  tri   n1146;
  tri   n1147;
  tri   n6160;
  tri   n1148;
  tri   n1149;
  tri   n6161;
  tri   n1150;
  tri   n1151;
  tri   n6162;
  tri   n1152;
  tri   n1153;
  tri   n6163;
  tri   n1154;
  tri   n1155;
  tri   n6164;
  tri   n1156;
  tri   n1157;
  tri   n6165;
  tri   n1158;
  tri   n1159;
  tri   n6166;
  tri   n1160;
  tri   n1161;
  tri   n6167;
  tri   n1162;
  tri   n1163;
  tri   n6168;
  tri   n1164;
  tri   n1165;
  tri   n6169;
  tri   n1166;
  tri   n1167;
  tri   n6170;
  tri   n1168;
  tri   n1169;
  tri   n6171;
  tri   n1170;
  tri   n1171;
  tri   n6172;
  tri   n1172;
  tri   n1173;
  tri   n6173;
  tri   n1174;
  tri   n1175;
  tri   n6174;
  tri   n1051;
  tri   n1052;
  tri   n6114;
  tri   n1053;
  tri   n1054;
  tri   n6115;
  tri   n1055;
  tri   n1056;
  tri   n6116;
  tri   n1057;
  tri   n1058;
  tri   n6117;
  tri   n1059;
  tri   n1060;
  tri   n6118;
  tri   n1061;
  tri   n1062;
  tri   n6119;
  tri   n1063;
  tri   n1064;
  tri   n6120;
  tri   n1065;
  tri   n1066;
  tri   n6121;
  tri   n1067;
  tri   n1068;
  tri   n6122;
  tri   n1069;
  tri   n1070;
  tri   n6123;
  tri   n1071;
  tri   n1072;
  tri   n6124;
  tri   n1073;
  tri   n1074;
  tri   n6125;
  tri   n1075;
  tri   n1076;
  tri   n6126;
  tri   n1077;
  tri   n1078;
  tri   n6127;
  tri   n1079;
  tri   n1080;
  tri   n6128;
  tri   n1081;
  tri   n1082;
  tri   n6129;
  tri   n1083;
  tri   n1084;
  tri   n6130;
  tri   n1085;
  tri   n1086;
  tri   n6131;
  tri   n1087;
  tri   n1088;
  tri   n6132;
  tri   n1089;
  tri   n1090;
  tri   n6133;
  tri   n1091;
  tri   n1092;
  tri   n6134;
  tri   n1093;
  tri   n1094;
  tri   n6135;
  tri   n1095;
  tri   n1096;
  tri   n6136;
  tri   n1097;
  tri   n1098;
  tri   n6137;
  tri   n1099;
  tri   n1100;
  tri   n6138;
  tri   n1101;
  tri   n1102;
  tri   n6139;
  tri   n1103;
  tri   n1104;
  tri   n6140;
  tri   n1105;
  tri   n1106;
  tri   n6141;
  tri   n1107;
  tri   n1108;
  tri   n6142;
  tri   n1110;
  tri   n1111;
  tri   n6143;
  tri   n1113;
  tri   n6144;
  tri   n989;
  tri   n988;
  tri   n990;
  tri   n991;
  tri   n6084;
  tri   n992;
  tri   n993;
  tri   n6085;
  tri   n994;
  tri   n995;
  tri   n6086;
  tri   n996;
  tri   n997;
  tri   n6087;
  tri   n998;
  tri   n999;
  tri   n6088;
  tri   n1000;
  tri   n1001;
  tri   n6089;
  tri   n1002;
  tri   n1003;
  tri   n6090;
  tri   n1004;
  tri   n1005;
  tri   n6091;
  tri   n1006;
  tri   n1007;
  tri   n6092;
  tri   n1008;
  tri   n1009;
  tri   n6093;
  tri   n1010;
  tri   n1011;
  tri   n6094;
  tri   n1012;
  tri   n1013;
  tri   n6095;
  tri   n1014;
  tri   n1015;
  tri   n6096;
  tri   n1016;
  tri   n1017;
  tri   n6097;
  tri   n1018;
  tri   n1019;
  tri   n6098;
  tri   n1020;
  tri   n1021;
  tri   n6099;
  tri   n1022;
  tri   n1023;
  tri   n6100;
  tri   n1024;
  tri   n1025;
  tri   n6101;
  tri   n1026;
  tri   n1027;
  tri   n6102;
  tri   n1028;
  tri   n1029;
  tri   n6103;
  tri   n1030;
  tri   n1031;
  tri   n6104;
  tri   n1032;
  tri   n1033;
  tri   n6105;
  tri   n1034;
  tri   n1035;
  tri   n6106;
  tri   n1036;
  tri   n1037;
  tri   n6107;
  tri   n1038;
  tri   n1039;
  tri   n6108;
  tri   n1040;
  tri   n1041;
  tri   n6109;
  tri   n1042;
  tri   n1043;
  tri   n6110;
  tri   n1045;
  tri   n1046;
  tri   n6111;
  tri   n1047;
  tri   n1048;
  tri   n6112;
  tri   n1049;
  tri   n1050;
  tri   n6113;
  tri   n925;
  tri   n927;
  tri   n928;
  tri   n6053;
  tri   n929;
  tri   n930;
  tri   n6054;
  tri   n931;
  tri   n932;
  tri   n6055;
  tri   n933;
  tri   n934;
  tri   n6056;
  tri   n935;
  tri   n936;
  tri   n6057;
  tri   n937;
  tri   n938;
  tri   n6058;
  tri   n939;
  tri   n940;
  tri   n6059;
  tri   n941;
  tri   n942;
  tri   n6060;
  tri   n943;
  tri   n944;
  tri   n6061;
  tri   n945;
  tri   n946;
  tri   n6062;
  tri   n947;
  tri   n948;
  tri   n6063;
  tri   n949;
  tri   n950;
  tri   n6064;
  tri   n951;
  tri   n952;
  tri   n6065;
  tri   n953;
  tri   n954;
  tri   n6066;
  tri   n955;
  tri   n956;
  tri   n6067;
  tri   n957;
  tri   n958;
  tri   n6068;
  tri   n959;
  tri   n960;
  tri   n6069;
  tri   n961;
  tri   n962;
  tri   n6070;
  tri   n963;
  tri   n964;
  tri   n6071;
  tri   n965;
  tri   n966;
  tri   n6072;
  tri   n967;
  tri   n968;
  tri   n6073;
  tri   n969;
  tri   n970;
  tri   n6074;
  tri   n971;
  tri   n972;
  tri   n6075;
  tri   n973;
  tri   n974;
  tri   n6076;
  tri   n975;
  tri   n976;
  tri   n6077;
  tri   n977;
  tri   n978;
  tri   n6078;
  tri   n979;
  tri   n980;
  tri   n6079;
  tri   n982;
  tri   n983;
  tri   n6080;
  tri   n984;
  tri   n985;
  tri   n6081;
  tri   n986;
  tri   n987;
  tri   n6082;
  tri   n6083;
  tri   n864;
  tri   n865;
  tri   n6022;
  tri   n866;
  tri   n867;
  tri   n6023;
  tri   n868;
  tri   n869;
  tri   n6024;
  tri   n870;
  tri   n871;
  tri   n6025;
  tri   n872;
  tri   n873;
  tri   n6026;
  tri   n874;
  tri   n875;
  tri   n6027;
  tri   n876;
  tri   n877;
  tri   n6028;
  tri   n878;
  tri   n879;
  tri   n6029;
  tri   n880;
  tri   n881;
  tri   n6030;
  tri   n882;
  tri   n883;
  tri   n6031;
  tri   n884;
  tri   n885;
  tri   n6032;
  tri   n886;
  tri   n887;
  tri   n6033;
  tri   n888;
  tri   n889;
  tri   n6034;
  tri   n890;
  tri   n891;
  tri   n6035;
  tri   n892;
  tri   n893;
  tri   n6036;
  tri   n894;
  tri   n895;
  tri   n6037;
  tri   n896;
  tri   n897;
  tri   n6038;
  tri   n898;
  tri   n899;
  tri   n6039;
  tri   n900;
  tri   n901;
  tri   n6040;
  tri   n902;
  tri   n903;
  tri   n6041;
  tri   n904;
  tri   n905;
  tri   n6042;
  tri   n906;
  tri   n907;
  tri   n6043;
  tri   n908;
  tri   n909;
  tri   n6044;
  tri   n910;
  tri   n911;
  tri   n6045;
  tri   n912;
  tri   n913;
  tri   n6046;
  tri   n914;
  tri   n915;
  tri   n6047;
  tri   n916;
  tri   n917;
  tri   n6048;
  tri   n918;
  tri   n919;
  tri   n6049;
  tri   n921;
  tri   n922;
  tri   n6050;
  tri   n923;
  tri   n924;
  tri   n6051;
  tri   n926;
  tri   n6052;
  tri   n801;
  tri   n803;
  tri   n804;
  tri   n5992;
  tri   n805;
  tri   n806;
  tri   n5993;
  tri   n807;
  tri   n808;
  tri   n5994;
  tri   n809;
  tri   n810;
  tri   n5995;
  tri   n811;
  tri   n812;
  tri   n5996;
  tri   n813;
  tri   n814;
  tri   n5997;
  tri   n815;
  tri   n816;
  tri   n5998;
  tri   n817;
  tri   n818;
  tri   n5999;
  tri   n819;
  tri   n820;
  tri   n6000;
  tri   n822;
  tri   n823;
  tri   n6001;
  tri   n824;
  tri   n825;
  tri   n6002;
  tri   n826;
  tri   n827;
  tri   n6003;
  tri   n828;
  tri   n829;
  tri   n6004;
  tri   n830;
  tri   n831;
  tri   n6005;
  tri   n832;
  tri   n833;
  tri   n6006;
  tri   n834;
  tri   n835;
  tri   n6007;
  tri   n836;
  tri   n837;
  tri   n6008;
  tri   n838;
  tri   n839;
  tri   n6009;
  tri   n840;
  tri   n841;
  tri   n6010;
  tri   n842;
  tri   n843;
  tri   n6011;
  tri   n844;
  tri   n845;
  tri   n6012;
  tri   n846;
  tri   n847;
  tri   n6013;
  tri   n848;
  tri   n849;
  tri   n6014;
  tri   n850;
  tri   n851;
  tri   n6015;
  tri   n852;
  tri   n853;
  tri   n6016;
  tri   n854;
  tri   n855;
  tri   n6017;
  tri   n856;
  tri   n857;
  tri   n6018;
  tri   n858;
  tri   n859;
  tri   n6019;
  tri   n860;
  tri   n861;
  tri   n6020;
  tri   n862;
  tri   n863;
  tri   n6021;
  tri   n738;
  tri   n739;
  tri   n5962;
  tri   n741;
  tri   n742;
  tri   n5963;
  tri   n744;
  tri   n745;
  tri   n5964;
  tri   n746;
  tri   n747;
  tri   n5965;
  tri   n749;
  tri   n750;
  tri   n5966;
  tri   n751;
  tri   n752;
  tri   n5967;
  tri   n753;
  tri   n754;
  tri   n5968;
  tri   n755;
  tri   n756;
  tri   n757;
  tri   n5969;
  tri   n758;
  tri   n759;
  tri   n5970;
  tri   n760;
  tri   n761;
  tri   n762;
  tri   n5971;
  tri   n763;
  tri   n764;
  tri   n5972;
  tri   n765;
  tri   n766;
  tri   n5973;
  tri   n767;
  tri   n768;
  tri   n5974;
  tri   n769;
  tri   n770;
  tri   n5975;
  tri   n771;
  tri   n772;
  tri   n5976;
  tri   n773;
  tri   n774;
  tri   n5977;
  tri   n775;
  tri   n776;
  tri   n5978;
  tri   n777;
  tri   n778;
  tri   n5979;
  tri   n779;
  tri   n780;
  tri   n5980;
  tri   n781;
  tri   n782;
  tri   n5981;
  tri   n783;
  tri   n784;
  tri   n5982;
  tri   n785;
  tri   n786;
  tri   n5983;
  tri   n787;
  tri   n788;
  tri   n5984;
  tri   n789;
  tri   n790;
  tri   n5985;
  tri   n791;
  tri   n792;
  tri   n5986;
  tri   n793;
  tri   n794;
  tri   n5987;
  tri   n795;
  tri   n796;
  tri   n5988;
  tri   n797;
  tri   n798;
  tri   n5989;
  tri   n799;
  tri   n800;
  tri   n5990;
  tri   n802;
  tri   n5991;
  tri   n666;
  tri   n667;
  tri   n664;
  tri   n668;
  tri   n669;
  tri   n1865;
  tri   n670;
  tri   n671;
  tri   n672;
  tri   n673;
  tri   n1867;
  tri   n674;
  tri   n675;
  tri   n676;
  tri   n677;
  tri   n1869;
  tri   n678;
  tri   n679;
  tri   n680;
  tri   n681;
  tri   n1871;
  tri   n682;
  tri   n683;
  tri   n684;
  tri   n685;
  tri   n1873;
  tri   n686;
  tri   n687;
  tri   n688;
  tri   n689;
  tri   n1875;
  tri   n690;
  tri   n691;
  tri   n692;
  tri   n693;
  tri   n1877;
  tri   n694;
  tri   n695;
  tri   n696;
  tri   n697;
  tri   n1879;
  tri   n698;
  tri   n699;
  tri   n700;
  tri   n701;
  tri   n1881;
  tri   n702;
  tri   n703;
  tri   n704;
  tri   n705;
  tri   n1883;
  tri   n706;
  tri   n707;
  tri   n708;
  tri   n709;
  tri   n1885;
  tri   n710;
  tri   n711;
  tri   n712;
  tri   n713;
  tri   n5953;
  tri   n715;
  tri   n716;
  tri   n5954;
  tri   n717;
  tri   n718;
  tri   n5955;
  tri   n720;
  tri   n721;
  tri   n722;
  tri   n5956;
  tri   n724;
  tri   n725;
  tri   n5957;
  tri   n726;
  tri   n727;
  tri   n728;
  tri   n5958;
  tri   n729;
  tri   n730;
  tri   n5959;
  tri   n732;
  tri   n733;
  tri   n5960;
  tri   n734;
  tri   n735;
  tri   n5961;
  tri   n591;
  tri   n592;
  tri   n593;
  tri   n590;
  tri   n594;
  tri   n595;
  tri   n1829;
  tri   n596;
  tri   n597;
  tri   n600;
  tri   n601;
  tri   n1831;
  tri   n602;
  tri   n603;
  tri   n604;
  tri   n605;
  tri   n1833;
  tri   n606;
  tri   n607;
  tri   n608;
  tri   n609;
  tri   n1835;
  tri   n610;
  tri   n611;
  tri   n612;
  tri   n613;
  tri   n1837;
  tri   n614;
  tri   n615;
  tri   n616;
  tri   n617;
  tri   n1839;
  tri   n618;
  tri   n619;
  tri   n620;
  tri   n621;
  tri   n1841;
  tri   n622;
  tri   n623;
  tri   n624;
  tri   n625;
  tri   n1843;
  tri   n626;
  tri   n627;
  tri   n628;
  tri   n629;
  tri   n1845;
  tri   n630;
  tri   n631;
  tri   n632;
  tri   n633;
  tri   n1847;
  tri   n634;
  tri   n635;
  tri   n636;
  tri   n637;
  tri   n1849;
  tri   n638;
  tri   n639;
  tri   n640;
  tri   n641;
  tri   n1851;
  tri   n642;
  tri   n643;
  tri   n644;
  tri   n645;
  tri   n1853;
  tri   n646;
  tri   n647;
  tri   n648;
  tri   n649;
  tri   n1855;
  tri   n650;
  tri   n651;
  tri   n652;
  tri   n653;
  tri   n1857;
  tri   n654;
  tri   n655;
  tri   n656;
  tri   n657;
  tri   n1859;
  tri   n658;
  tri   n659;
  tri   n660;
  tri   n661;
  tri   n1861;
  tri   n662;
  tri   n663;
  tri   n665;
  tri   n1863;
  tri   n517;
  tri   n516;
  tri   n518;
  tri   n519;
  tri   n1618;
  tri   n520;
  tri   n521;
  tri   n522;
  tri   n523;
  tri   n1621;
  tri   n524;
  tri   n525;
  tri   n526;
  tri   n527;
  tri   n1624;
  tri   n528;
  tri   n529;
  tri   n530;
  tri   n531;
  tri   n1627;
  tri   n532;
  tri   n533;
  tri   n534;
  tri   n535;
  tri   n1630;
  tri   n536;
  tri   n537;
  tri   n538;
  tri   n539;
  tri   n1633;
  tri   n540;
  tri   n541;
  tri   n542;
  tri   n543;
  tri   n1636;
  tri   n544;
  tri   n545;
  tri   n546;
  tri   n547;
  tri   n1639;
  tri   n548;
  tri   n549;
  tri   n550;
  tri   n551;
  tri   n1642;
  tri   n552;
  tri   n553;
  tri   n554;
  tri   n555;
  tri   n1645;
  tri   n556;
  tri   n557;
  tri   n558;
  tri   n559;
  tri   n1648;
  tri   n560;
  tri   n561;
  tri   n562;
  tri   n563;
  tri   n1651;
  tri   n564;
  tri   n565;
  tri   n566;
  tri   n567;
  tri   n1654;
  tri   n568;
  tri   n569;
  tri   n570;
  tri   n571;
  tri   n1657;
  tri   n572;
  tri   n573;
  tri   n574;
  tri   n575;
  tri   n1660;
  tri   n576;
  tri   n577;
  tri   n578;
  tri   n579;
  tri   n1663;
  tri   n580;
  tri   n581;
  tri   n582;
  tri   n583;
  tri   n1666;
  tri   n584;
  tri   n585;
  tri   n586;
  tri   n587;
  tri   n1669;
  tri   n588;
  tri   n589;
  tri   n1673;
  tri   n470;
  tri   n471;
  tri   n18189;
  tri   n473;
  tri   n474;
  tri   n476;
  tri   n477;
  tri   n1559;
  tri   n478;
  tri   n479;
  tri   n482;
  tri   n483;
  tri   n1591;
  tri   n484;
  tri   n485;
  tri   n486;
  tri   n487;
  tri   n1594;
  tri   n488;
  tri   n489;
  tri   n490;
  tri   n491;
  tri   n1597;
  tri   n492;
  tri   n493;
  tri   n494;
  tri   n495;
  tri   n1600;
  tri   n496;
  tri   n497;
  tri   n498;
  tri   n499;
  tri   n1603;
  tri   n500;
  tri   n501;
  tri   n502;
  tri   n503;
  tri   n1606;
  tri   n504;
  tri   n505;
  tri   n506;
  tri   n507;
  tri   n1609;
  tri   n508;
  tri   n509;
  tri   n510;
  tri   n511;
  tri   n1612;
  tri   n512;
  tri   n513;
  tri   n514;
  tri   n515;
  tri   n1615;
  tri   N76;
  tri   N77;
  tri   N73;
  tri   N75;
  tri   P1_N5897;
  tri   P1_N5898;
  tri   P1_N5900;
  tri   P1_N5899;
  tri   P1_N5902;
  tri   P1_N5901;
  tri   P1_N5904;
  tri   P1_N5903;
  tri   P1_N5906;
  tri   P1_N5905;
  tri   P1_N5834;
  tri   P1_N5836;
  tri   P1_N5835;
  tri   P1_N5838;
  tri   P1_N5837;
  tri   P1_N5840;
  tri   P1_N5839;
  tri   P1_N5842;
  tri   P1_N5841;
  tri   P1_N5846;
  tri   P1_N5845;
  tri   P1_N5848;
  tri   P1_N5847;
  tri   P1_N5850;
  tri   P1_N5849;
  tri   P1_N5852;
  tri   P1_N5851;
  tri   P1_N5854;
  tri   P1_N5853;
  tri   P1_N5856;
  tri   P1_N5855;
  tri   P1_N5858;
  tri   P1_N5857;
  tri   P1_N5860;
  tri   P1_N5859;
  tri   P1_N5862;
  tri   P1_N5861;
  tri   P1_N5864;
  tri   P1_N5863;
  tri   P1_N5866;
  tri   P1_N5865;
  tri   P1_N5868;
  tri   P1_N5867;
  tri   P1_N5870;
  tri   P1_N5869;
  tri   P1_N5872;
  tri   P1_N5871;
  tri   P1_N5874;
  tri   P1_N5873;
  tri   P1_N5876;
  tri   P1_N5875;
  tri   P1_N5878;
  tri   P1_N5877;
  tri   P1_N5880;
  tri   P1_N5879;
  tri   P1_N5882;
  tri   P1_N5881;
  tri   P1_N5884;
  tri   P1_N5883;
  tri   P1_N5886;
  tri   P1_N5885;
  tri   P1_N5888;
  tri   P1_N5887;
  tri   P1_N5890;
  tri   P1_N5889;
  tri   P1_N5892;
  tri   P1_N5891;
  tri   P1_N5894;
  tri   P1_N5893;
  tri   P1_N5896;
  tri   P1_N5895;
  tri   P1_N5772;
  tri   P1_N5774;
  tri   P1_N5773;
  tri   P1_N5776;
  tri   P1_N5775;
  tri   P1_N5778;
  tri   P1_N5777;
  tri   P1_N5780;
  tri   P1_N5779;
  tri   P1_N5782;
  tri   P1_N5781;
  tri   P1_N5784;
  tri   P1_N5783;
  tri   P1_N5786;
  tri   P1_N5785;
  tri   P1_N5788;
  tri   P1_N5787;
  tri   P1_N5790;
  tri   P1_N5789;
  tri   P1_N5792;
  tri   P1_N5791;
  tri   P1_N5794;
  tri   P1_N5793;
  tri   P1_N5796;
  tri   P1_N5795;
  tri   P1_N5798;
  tri   P1_N5797;
  tri   P1_N5800;
  tri   P1_N5799;
  tri   P1_N5802;
  tri   P1_N5801;
  tri   P1_N5804;
  tri   P1_N5803;
  tri   P1_N5806;
  tri   P1_N5805;
  tri   P1_N5808;
  tri   P1_N5807;
  tri   P1_N5810;
  tri   P1_N5809;
  tri   P1_N5812;
  tri   P1_N5811;
  tri   P1_N5814;
  tri   P1_N5813;
  tri   P1_N5816;
  tri   P1_N5815;
  tri   P1_N5818;
  tri   P1_N5817;
  tri   P1_N5820;
  tri   P1_N5819;
  tri   P1_N5822;
  tri   P1_N5821;
  tri   P1_N5824;
  tri   P1_N5823;
  tri   P1_N5826;
  tri   P1_N5825;
  tri   P1_N5828;
  tri   P1_N5827;
  tri   P1_N5830;
  tri   P1_N5829;
  tri   P1_N5832;
  tri   P1_N5831;
  tri   P1_N5833;
  tri   P1_N5712;
  tri   P1_N5711;
  tri   P1_N5714;
  tri   P1_N5713;
  tri   P1_N5716;
  tri   P1_N5715;
  tri   P1_N5718;
  tri   P1_N5717;
  tri   P1_N5720;
  tri   P1_N5719;
  tri   P1_N5722;
  tri   P1_N5721;
  tri   P1_N5724;
  tri   P1_N5723;
  tri   P1_N5726;
  tri   P1_N5725;
  tri   P1_N5728;
  tri   P1_N5727;
  tri   P1_N5730;
  tri   P1_N5729;
  tri   P1_N5732;
  tri   P1_N5731;
  tri   P1_N5734;
  tri   P1_N5733;
  tri   P1_N5736;
  tri   P1_N5735;
  tri   P1_N5738;
  tri   P1_N5737;
  tri   P1_N5740;
  tri   P1_N5739;
  tri   P1_N5742;
  tri   P1_N5741;
  tri   P1_N5744;
  tri   P1_N5743;
  tri   P1_N5746;
  tri   P1_N5745;
  tri   P1_N5748;
  tri   P1_N5747;
  tri   P1_N5750;
  tri   P1_N5749;
  tri   P1_N5752;
  tri   P1_N5751;
  tri   P1_N5758;
  tri   P1_N5757;
  tri   P1_N5760;
  tri   P1_N5759;
  tri   P1_N5762;
  tri   P1_N5761;
  tri   P1_N5764;
  tri   P1_N5763;
  tri   P1_N5766;
  tri   P1_N5765;
  tri   P1_N5768;
  tri   P1_N5767;
  tri   P1_N5770;
  tri   P1_N5769;
  tri   P1_N5771;
  tri   P1_N5644;
  tri   P1_N5646;
  tri   P1_N5645;
  tri   P1_N5648;
  tri   P1_N5647;
  tri   P1_N5652;
  tri   P1_N5651;
  tri   P1_N5656;
  tri   P1_N5655;
  tri   P1_N5658;
  tri   P1_N5657;
  tri   P1_N5660;
  tri   P1_N5659;
  tri   P1_N5662;
  tri   P1_N5661;
  tri   P1_N5664;
  tri   P1_N5663;
  tri   P1_N5666;
  tri   P1_N5665;
  tri   P1_N5668;
  tri   P1_N5667;
  tri   P1_N5670;
  tri   P1_N5669;
  tri   P1_N5672;
  tri   P1_N5671;
  tri   P1_N5674;
  tri   P1_N5673;
  tri   P1_N5676;
  tri   P1_N5675;
  tri   P1_N5678;
  tri   P1_N5677;
  tri   P1_N5680;
  tri   P1_N5679;
  tri   P1_N5682;
  tri   P1_N5681;
  tri   P1_N5684;
  tri   P1_N5683;
  tri   P1_N5686;
  tri   P1_N5685;
  tri   P1_N5688;
  tri   P1_N5687;
  tri   P1_N5690;
  tri   P1_N5689;
  tri   P1_N5692;
  tri   P1_N5691;
  tri   P1_N5694;
  tri   P1_N5693;
  tri   P1_N5696;
  tri   P1_N5695;
  tri   P1_N5698;
  tri   P1_N5697;
  tri   P1_N5700;
  tri   P1_N5699;
  tri   P1_N5702;
  tri   P1_N5701;
  tri   P1_N5704;
  tri   P1_N5703;
  tri   P1_N5708;
  tri   P1_N5707;
  tri   P1_N5592;
  tri   P1_N5591;
  tri   P1_N5594;
  tri   P1_N5593;
  tri   P1_N5596;
  tri   P1_N5595;
  tri   P1_N5598;
  tri   P1_N5597;
  tri   P1_N5600;
  tri   P1_N5599;
  tri   P1_N5602;
  tri   P1_N5601;
  tri   P1_N5604;
  tri   P1_N5603;
  tri   P1_N5606;
  tri   P1_N5605;
  tri   P1_N5608;
  tri   P1_N5607;
  tri   P1_N5610;
  tri   P1_N5609;
  tri   P1_N5612;
  tri   P1_N5611;
  tri   P1_N5614;
  tri   P1_N5613;
  tri   P1_N5616;
  tri   P1_N5615;
  tri   P1_N5618;
  tri   P1_N5617;
  tri   P1_N5620;
  tri   P1_N5619;
  tri   P1_N5622;
  tri   P1_N5621;
  tri   P1_N5624;
  tri   P1_N5623;
  tri   P1_N5626;
  tri   P1_N5625;
  tri   P1_N5628;
  tri   P1_N5627;
  tri   P1_N5630;
  tri   P1_N5629;
  tri   P1_N5632;
  tri   P1_N5631;
  tri   P1_N5634;
  tri   P1_N5633;
  tri   P1_N5636;
  tri   P1_N5635;
  tri   P1_N5638;
  tri   P1_N5637;
  tri   P1_N5640;
  tri   P1_N5639;
  tri   P1_N5642;
  tri   P1_N5641;
  tri   P1_N5643;
  tri   P2_N6540;
  tri   P2_N6539;
  tri   P2_N6604;
  tri   P2_N6603;
  tri   P2_N5803;
  tri   P2_N5804;
  tri   P2_N5806;
  tri   P2_N5805;
  tri   P2_N5808;
  tri   P2_N5807;
  tri   P2_N5810;
  tri   P2_N5809;
  tri   P2_N5812;
  tri   P2_N5811;
  tri   P2_N5814;
  tri   P2_N5813;
  tri   P2_N5816;
  tri   P2_N5815;
  tri   P2_N5818;
  tri   P2_N5817;
  tri   P2_N5820;
  tri   P2_N5819;
  tri   P2_N5822;
  tri   P2_N5821;
  tri   P2_N5824;
  tri   P2_N5823;
  tri   P2_N5826;
  tri   P2_N5825;
  tri   P2_N5828;
  tri   P2_N5827;
  tri   P2_N5740;
  tri   P2_N5742;
  tri   P2_N5741;
  tri   P2_N5744;
  tri   P2_N5743;
  tri   P2_N5746;
  tri   P2_N5745;
  tri   P2_N5748;
  tri   P2_N5747;
  tri   P2_N5750;
  tri   P2_N5749;
  tri   P2_N5752;
  tri   P2_N5751;
  tri   P2_N5754;
  tri   P2_N5753;
  tri   P2_N5756;
  tri   P2_N5755;
  tri   P2_N5758;
  tri   P2_N5757;
  tri   P2_N5760;
  tri   P2_N5759;
  tri   P2_N5762;
  tri   P2_N5761;
  tri   P2_N5764;
  tri   P2_N5763;
  tri   P2_N5768;
  tri   P2_N5767;
  tri   P2_N5770;
  tri   P2_N5769;
  tri   P2_N5772;
  tri   P2_N5771;
  tri   P2_N5774;
  tri   P2_N5773;
  tri   P2_N5776;
  tri   P2_N5775;
  tri   P2_N5778;
  tri   P2_N5777;
  tri   P2_N5780;
  tri   P2_N5779;
  tri   P2_N5782;
  tri   P2_N5781;
  tri   P2_N5784;
  tri   P2_N5783;
  tri   P2_N5786;
  tri   P2_N5785;
  tri   P2_N5788;
  tri   P2_N5787;
  tri   P2_N5790;
  tri   P2_N5789;
  tri   P2_N5792;
  tri   P2_N5791;
  tri   P2_N5794;
  tri   P2_N5793;
  tri   P2_N5796;
  tri   P2_N5795;
  tri   P2_N5798;
  tri   P2_N5797;
  tri   P2_N5800;
  tri   P2_N5799;
  tri   P2_N5802;
  tri   P2_N5801;
  tri   P2_N5680;
  tri   P2_N5679;
  tri   P2_N5682;
  tri   P2_N5681;
  tri   P2_N5684;
  tri   P2_N5683;
  tri   P2_N5686;
  tri   P2_N5685;
  tri   P2_N5688;
  tri   P2_N5687;
  tri   P2_N5690;
  tri   P2_N5689;
  tri   P2_N5692;
  tri   P2_N5691;
  tri   P2_N5694;
  tri   P2_N5693;
  tri   P2_N5696;
  tri   P2_N5695;
  tri   P2_N5698;
  tri   P2_N5697;
  tri   P2_N5700;
  tri   P2_N5699;
  tri   P2_N5702;
  tri   P2_N5701;
  tri   P2_N5704;
  tri   P2_N5703;
  tri   P2_N5706;
  tri   P2_N5705;
  tri   P2_N5708;
  tri   P2_N5707;
  tri   P2_N5710;
  tri   P2_N5709;
  tri   P2_N5712;
  tri   P2_N5711;
  tri   P2_N5714;
  tri   P2_N5713;
  tri   P2_N5716;
  tri   P2_N5715;
  tri   P2_N5718;
  tri   P2_N5717;
  tri   P2_N5720;
  tri   P2_N5719;
  tri   P2_N5722;
  tri   P2_N5721;
  tri   P2_N5724;
  tri   P2_N5723;
  tri   P2_N5726;
  tri   P2_N5725;
  tri   P2_N5728;
  tri   P2_N5727;
  tri   P2_N5730;
  tri   P2_N5729;
  tri   P2_N5732;
  tri   P2_N5731;
  tri   P2_N5734;
  tri   P2_N5733;
  tri   P2_N5736;
  tri   P2_N5735;
  tri   P2_N5738;
  tri   P2_N5737;
  tri   P2_N5739;
  tri   P2_N5613;
  tri   P2_N5614;
  tri   P2_N5616;
  tri   P2_N5615;
  tri   P2_N5618;
  tri   P2_N5617;
  tri   P2_N5620;
  tri   P2_N5619;
  tri   P2_N5622;
  tri   P2_N5621;
  tri   P2_N5624;
  tri   P2_N5623;
  tri   P2_N5626;
  tri   P2_N5625;
  tri   P2_N5630;
  tri   P2_N5629;
  tri   P2_N5634;
  tri   P2_N5633;
  tri   P2_N5636;
  tri   P2_N5635;
  tri   P2_N5638;
  tri   P2_N5637;
  tri   P2_N5640;
  tri   P2_N5639;
  tri   P2_N5642;
  tri   P2_N5641;
  tri   P2_N5644;
  tri   P2_N5643;
  tri   P2_N5646;
  tri   P2_N5645;
  tri   P2_N5648;
  tri   P2_N5647;
  tri   P2_N5650;
  tri   P2_N5649;
  tri   P2_N5652;
  tri   P2_N5651;
  tri   P2_N5654;
  tri   P2_N5653;
  tri   P2_N5656;
  tri   P2_N5655;
  tri   P2_N5658;
  tri   P2_N5657;
  tri   P2_N5660;
  tri   P2_N5659;
  tri   P2_N5662;
  tri   P2_N5661;
  tri   P2_N5664;
  tri   P2_N5663;
  tri   P2_N5666;
  tri   P2_N5665;
  tri   P2_N5668;
  tri   P2_N5667;
  tri   P2_N5670;
  tri   P2_N5669;
  tri   P2_N5672;
  tri   P2_N5671;
  tri   P2_N5674;
  tri   P2_N5673;
  tri   P2_N5550;
  tri   P2_N5552;
  tri   P2_N5551;
  tri   P2_N5554;
  tri   P2_N5553;
  tri   P2_N5556;
  tri   P2_N5555;
  tri   P2_N5558;
  tri   P2_N5557;
  tri   P2_N5560;
  tri   P2_N5559;
  tri   P2_N5562;
  tri   P2_N5561;
  tri   P2_N5564;
  tri   P2_N5563;
  tri   P2_N5566;
  tri   P2_N5565;
  tri   P2_N5568;
  tri   P2_N5567;
  tri   P2_N5570;
  tri   P2_N5569;
  tri   P2_N5574;
  tri   P2_N5573;
  tri   P2_N5578;
  tri   P2_N5577;
  tri   P2_N5580;
  tri   P2_N5579;
  tri   P2_N5582;
  tri   P2_N5581;
  tri   P2_N5584;
  tri   P2_N5583;
  tri   P2_N5586;
  tri   P2_N5585;
  tri   P2_N5588;
  tri   P2_N5587;
  tri   P2_N5590;
  tri   P2_N5589;
  tri   P2_N5592;
  tri   P2_N5591;
  tri   P2_N5594;
  tri   P2_N5593;
  tri   P2_N5596;
  tri   P2_N5595;
  tri   P2_N5598;
  tri   P2_N5597;
  tri   P2_N5600;
  tri   P2_N5599;
  tri   P2_N5602;
  tri   P2_N5601;
  tri   P2_N5604;
  tri   P2_N5603;
  tri   P2_N5606;
  tri   P2_N5605;
  tri   P2_N5608;
  tri   P2_N5607;
  tri   P2_N5610;
  tri   P2_N5609;
  tri   P2_N5612;
  tri   P2_N5611;
  tri   P2_N5514;
  tri   P2_N5513;
  tri   P2_N5516;
  tri   P2_N5515;
  tri   P2_N5518;
  tri   P2_N5517;
  tri   P2_N5520;
  tri   P2_N5519;
  tri   P2_N5522;
  tri   P2_N5521;
  tri   P2_N5524;
  tri   P2_N5523;
  tri   P2_N5526;
  tri   P2_N5525;
  tri   P2_N5528;
  tri   P2_N5527;
  tri   P2_N5530;
  tri   P2_N5529;
  tri   P2_N5532;
  tri   P2_N5531;
  tri   P2_N5534;
  tri   P2_N5533;
  tri   P2_N5536;
  tri   P2_N5535;
  tri   P2_N5538;
  tri   P2_N5537;
  tri   P2_N5540;
  tri   P2_N5539;
  tri   P2_N5542;
  tri   P2_N5541;
  tri   P2_N5544;
  tri   P2_N5543;
  tri   P2_N5546;
  tri   P2_N5545;
  tri   P2_N5548;
  tri   P2_N5547;
  tri   P2_N5549;
  tri   P2_lt_696_n27;
  tri   P2_lt_696_n25;
  tri   P2_lt_696_n22;
  tri   P2_lt_696_n21;
  tri   P2_lt_696_n20;
  tri   P2_lt_696_n19;
  tri   P2_lt_696_n18;
  tri   P2_lt_696_n17;
  tri   P2_lt_696_n16;
  tri   P2_lt_696_n15;
  tri   P2_lt_696_n12;
  tri   P2_lt_696_n11;
  tri   P2_lt_696_n10;
  tri   P2_lt_696_n9;
  tri   P2_lt_696_n8;
  tri   P2_lt_696_n7;
  tri   P2_lt_696_n6;
  tri   P2_lt_696_n4;
  tri   P2_lt_696_n3;
  tri   P2_lt_696_n2;
  tri   P2_lt_696_n142;
  tri   P2_lt_696_n140;
  tri   P2_lt_696_n139;
  tri   P2_lt_696_n138;
  tri   P2_lt_696_n137;
  tri   P2_lt_696_n136;
  tri   P2_lt_696_n135;
  tri   P2_lt_696_n132;
  tri   P2_lt_696_n131;
  tri   P2_lt_696_n130;
  tri   P2_lt_696_n129;
  tri   P2_lt_696_n128;
  tri   P2_lt_696_n127;
  tri   P2_lt_696_n126;
  tri   P2_lt_696_n125;
  tri   P2_lt_696_n122;
  tri   P2_lt_696_n121;
  tri   P2_lt_696_n120;
  tri   P2_lt_696_n119;
  tri   P2_lt_696_n118;
  tri   P2_lt_696_n117;
  tri   P2_lt_696_n116;
  tri   P2_lt_696_n115;
  tri   P2_lt_696_n113;
  tri   P2_lt_696_n112;
  tri   P2_lt_696_n110;
  tri   P2_lt_696_n109;
  tri   P2_lt_696_n108;
  tri   P2_lt_696_n107;
  tri   P2_lt_696_n106;
  tri   P2_lt_696_n105;
  tri   P2_lt_696_n102;
  tri   P2_lt_696_n101;
  tri   P2_lt_696_n100;
  tri   P2_lt_696_n99;
  tri   P2_lt_696_n98;
  tri   P2_lt_696_n97;
  tri   P2_lt_696_n96;
  tri   P2_lt_696_n95;
  tri   P2_lt_696_n92;
  tri   P2_lt_696_n91;
  tri   P2_lt_696_n90;
  tri   P2_lt_696_n89;
  tri   P2_lt_696_n88;
  tri   P2_lt_696_n87;
  tri   P2_lt_696_n86;
  tri   P2_lt_696_n85;
  tri   P2_lt_696_n82;
  tri   P2_lt_696_n81;
  tri   P2_lt_696_n80;
  tri   P2_lt_696_n79;
  tri   P2_lt_696_n78;
  tri   P2_lt_696_n77;
  tri   P2_lt_696_n76;
  tri   P2_lt_696_n75;
  tri   P2_lt_696_n72;
  tri   P2_lt_696_n71;
  tri   P2_lt_696_n70;
  tri   P2_lt_696_n69;
  tri   P2_lt_696_n68;
  tri   P2_lt_696_n67;
  tri   P2_lt_696_n66;
  tri   P2_lt_696_n65;
  tri   P2_lt_696_n62;
  tri   P2_lt_696_n61;
  tri   P2_lt_696_n60;
  tri   P2_lt_696_n59;
  tri   P2_lt_696_n58;
  tri   P2_lt_696_n57;
  tri   P2_lt_696_n56;
  tri   P2_lt_696_n55;
  tri   P2_lt_696_n52;
  tri   P2_lt_696_n51;
  tri   P2_lt_696_n50;
  tri   P2_lt_696_n49;
  tri   P2_lt_696_n48;
  tri   P2_lt_696_n47;
  tri   P2_lt_696_n46;
  tri   P2_lt_696_n45;
  tri   P2_lt_696_n42;
  tri   P2_lt_696_n41;
  tri   P2_lt_696_n40;
  tri   P2_lt_696_n39;
  tri   P2_lt_696_n38;
  tri   P2_lt_696_n37;
  tri   P2_lt_696_n36;
  tri   P2_lt_696_n35;
  tri   P2_lt_696_n32;
  tri   P2_lt_696_n31;
  tri   P2_lt_696_n28;
  tri   P2_lt_696_n26;
  tri   P2_lt_696_n30;
  tri   P2_lt_696_n29;
  tri   P2_lt_696_n1;
  tri   P2_lt_696_n5;
  tri   P2_lt_696_n14;
  tri   P2_lt_696_n13;
  tri   P2_lt_696_n24;
  tri   P2_lt_696_n23;
  tri   P2_lt_696_n34;
  tri   P2_lt_696_n33;
  tri   P2_lt_696_n44;
  tri   P2_lt_696_n43;
  tri   P2_lt_696_n54;
  tri   P2_lt_696_n53;
  tri   P2_lt_696_n64;
  tri   P2_lt_696_n63;
  tri   P2_lt_696_n74;
  tri   P2_lt_696_n73;
  tri   P2_lt_696_n84;
  tri   P2_lt_696_n83;
  tri   P2_lt_696_n94;
  tri   P2_lt_696_n93;
  tri   P2_lt_696_n104;
  tri   P2_lt_696_n103;
  tri   P2_lt_696_n114;
  tri   P2_lt_696_n124;
  tri   P2_lt_696_n123;
  tri   P2_lt_696_n134;
  tri   P2_lt_696_n133;
  tri   P2_lt_696_n143;
  tri   P2_lt_696_n156;
  tri   P2_lt_696_n155;
  tri   P2_lt_696_n154;
  tri   P2_lt_696_n153;
  tri   P2_lt_696_n152;
  tri   P2_lt_696_n151;
  tri   P2_lt_696_n150;
  tri   P2_lt_696_n149;
  tri   P2_lt_696_n148;
  tri   P2_lt_696_n147;
  tri   P2_lt_696_n146;
  tri   P2_lt_696_n145;
  tri   P2_lt_696_n144;
  tri   P2_lt_696_n141;
  tri   P2_lt_734_n107;
  tri   P2_lt_734_n105;
  tri   P2_lt_734_n102;
  tri   P2_lt_734_n101;
  tri   P2_lt_734_n100;
  tri   P2_lt_734_n99;
  tri   P2_lt_734_n98;
  tri   P2_lt_734_n97;
  tri   P2_lt_734_n96;
  tri   P2_lt_734_n95;
  tri   P2_lt_734_n92;
  tri   P2_lt_734_n91;
  tri   P2_lt_734_n90;
  tri   P2_lt_734_n89;
  tri   P2_lt_734_n88;
  tri   P2_lt_734_n87;
  tri   P2_lt_734_n86;
  tri   P2_lt_734_n85;
  tri   P2_lt_734_n82;
  tri   P2_lt_734_n81;
  tri   P2_lt_734_n80;
  tri   P2_lt_734_n79;
  tri   P2_lt_734_n78;
  tri   P2_lt_734_n77;
  tri   P2_lt_734_n76;
  tri   P2_lt_734_n75;
  tri   P2_lt_734_n72;
  tri   P2_lt_734_n71;
  tri   P2_lt_734_n70;
  tri   P2_lt_734_n69;
  tri   P2_lt_734_n68;
  tri   P2_lt_734_n67;
  tri   P2_lt_734_n66;
  tri   P2_lt_734_n65;
  tri   P2_lt_734_n62;
  tri   P2_lt_734_n61;
  tri   P2_lt_734_n60;
  tri   P2_lt_734_n59;
  tri   P2_lt_734_n58;
  tri   P2_lt_734_n57;
  tri   P2_lt_734_n56;
  tri   P2_lt_734_n55;
  tri   P2_lt_734_n52;
  tri   P2_lt_734_n51;
  tri   P2_lt_734_n50;
  tri   P2_lt_734_n49;
  tri   P2_lt_734_n48;
  tri   P2_lt_734_n47;
  tri   P2_lt_734_n46;
  tri   P2_lt_734_n45;
  tri   P2_lt_734_n42;
  tri   P2_lt_734_n41;
  tri   P2_lt_734_n40;
  tri   P2_lt_734_n39;
  tri   P2_lt_734_n38;
  tri   P2_lt_734_n37;
  tri   P2_lt_734_n36;
  tri   P2_lt_734_n35;
  tri   P2_lt_734_n32;
  tri   P2_lt_734_n31;
  tri   P2_lt_734_n30;
  tri   P2_lt_734_n29;
  tri   P2_lt_734_n28;
  tri   P2_lt_734_n27;
  tri   P2_lt_734_n26;
  tri   P2_lt_734_n25;
  tri   P2_lt_734_n22;
  tri   P2_lt_734_n21;
  tri   P2_lt_734_n20;
  tri   P2_lt_734_n19;
  tri   P2_lt_734_n18;
  tri   P2_lt_734_n17;
  tri   P2_lt_734_n16;
  tri   P2_lt_734_n15;
  tri   P2_lt_734_n12;
  tri   P2_lt_734_n11;
  tri   P2_lt_734_n10;
  tri   P2_lt_734_n9;
  tri   P2_lt_734_n8;
  tri   P2_lt_734_n7;
  tri   P2_lt_734_n6;
  tri   P2_lt_734_n4;
  tri   P2_lt_734_n3;
  tri   P2_lt_734_n2;
  tri   P2_lt_734_n1;
  tri   P2_lt_734_n5;
  tri   P2_lt_734_n14;
  tri   P2_lt_734_n13;
  tri   P2_lt_734_n24;
  tri   P2_lt_734_n23;
  tri   P2_lt_734_n34;
  tri   P2_lt_734_n33;
  tri   P2_lt_734_n44;
  tri   P2_lt_734_n43;
  tri   P2_lt_734_n54;
  tri   P2_lt_734_n53;
  tri   P2_lt_734_n64;
  tri   P2_lt_734_n63;
  tri   P2_lt_734_n74;
  tri   P2_lt_734_n73;
  tri   P2_lt_734_n84;
  tri   P2_lt_734_n83;
  tri   P2_lt_734_n94;
  tri   P2_lt_734_n93;
  tri   P2_lt_734_n104;
  tri   P2_lt_734_n103;
  tri   P2_lt_734_n156;
  tri   P2_lt_734_n155;
  tri   P2_lt_734_n154;
  tri   P2_lt_734_n153;
  tri   P2_lt_734_n152;
  tri   P2_lt_734_n151;
  tri   P2_lt_734_n150;
  tri   P2_lt_734_n149;
  tri   P2_lt_734_n148;
  tri   P2_lt_734_n147;
  tri   P2_lt_734_n146;
  tri   P2_lt_734_n145;
  tri   P2_lt_734_n144;
  tri   P2_lt_734_n143;
  tri   P2_lt_734_n142;
  tri   P2_lt_734_n141;
  tri   P2_lt_734_n140;
  tri   P2_lt_734_n139;
  tri   P2_lt_734_n138;
  tri   P2_lt_734_n137;
  tri   P2_lt_734_n136;
  tri   P2_lt_734_n135;
  tri   P2_lt_734_n134;
  tri   P2_lt_734_n133;
  tri   P2_lt_734_n132;
  tri   P2_lt_734_n131;
  tri   P2_lt_734_n130;
  tri   P2_lt_734_n129;
  tri   P2_lt_734_n128;
  tri   P2_lt_734_n127;
  tri   P2_lt_734_n126;
  tri   P2_lt_734_n125;
  tri   P2_lt_734_n124;
  tri   P2_lt_734_n123;
  tri   P2_lt_734_n122;
  tri   P2_lt_734_n121;
  tri   P2_lt_734_n120;
  tri   P2_lt_734_n119;
  tri   P2_lt_734_n118;
  tri   P2_lt_734_n117;
  tri   P2_lt_734_n116;
  tri   P2_lt_734_n115;
  tri   P2_lt_734_n114;
  tri   P2_lt_734_n108;
  tri   P2_lt_734_n113;
  tri   P2_lt_734_n112;
  tri   P2_lt_734_n106;
  tri   P2_lt_734_n110;
  tri   P2_lt_734_n109;
  tri   P2_lt_742_n70;
  tri   P2_lt_742_n68;
  tri   P2_lt_742_n67;
  tri   P2_lt_742_n66;
  tri   P2_lt_742_n65;
  tri   P2_lt_742_n62;
  tri   P2_lt_742_n61;
  tri   P2_lt_742_n60;
  tri   P2_lt_742_n59;
  tri   P2_lt_742_n58;
  tri   P2_lt_742_n57;
  tri   P2_lt_742_n56;
  tri   P2_lt_742_n55;
  tri   P2_lt_742_n52;
  tri   P2_lt_742_n51;
  tri   P2_lt_742_n50;
  tri   P2_lt_742_n49;
  tri   P2_lt_742_n48;
  tri   P2_lt_742_n47;
  tri   P2_lt_742_n46;
  tri   P2_lt_742_n45;
  tri   P2_lt_742_n42;
  tri   P2_lt_742_n41;
  tri   P2_lt_742_n40;
  tri   P2_lt_742_n39;
  tri   P2_lt_742_n38;
  tri   P2_lt_742_n37;
  tri   P2_lt_742_n36;
  tri   P2_lt_742_n35;
  tri   P2_lt_742_n32;
  tri   P2_lt_742_n31;
  tri   P2_lt_742_n30;
  tri   P2_lt_742_n29;
  tri   P2_lt_742_n28;
  tri   P2_lt_742_n27;
  tri   P2_lt_742_n26;
  tri   P2_lt_742_n25;
  tri   P2_lt_742_n22;
  tri   P2_lt_742_n21;
  tri   P2_lt_742_n20;
  tri   P2_lt_742_n19;
  tri   P2_lt_742_n18;
  tri   P2_lt_742_n17;
  tri   P2_lt_742_n16;
  tri   P2_lt_742_n15;
  tri   P2_lt_742_n12;
  tri   P2_lt_742_n11;
  tri   P2_lt_742_n10;
  tri   P2_lt_742_n9;
  tri   P2_lt_742_n8;
  tri   P2_lt_742_n7;
  tri   P2_lt_742_n6;
  tri   P2_lt_742_n4;
  tri   P2_lt_742_n3;
  tri   P2_lt_742_n2;
  tri   P2_lt_742_n44;
  tri   P2_lt_742_n43;
  tri   P2_lt_742_n54;
  tri   P2_lt_742_n53;
  tri   P2_lt_742_n64;
  tri   P2_lt_742_n63;
  tri   P2_lt_742_n156;
  tri   P2_lt_742_n155;
  tri   P2_lt_742_n154;
  tri   P2_lt_742_n153;
  tri   P2_lt_742_n152;
  tri   P2_lt_742_n151;
  tri   P2_lt_742_n150;
  tri   P2_lt_742_n149;
  tri   P2_lt_742_n148;
  tri   P2_lt_742_n147;
  tri   P2_lt_742_n146;
  tri   P2_lt_742_n145;
  tri   P2_lt_742_n144;
  tri   P2_lt_742_n143;
  tri   P2_lt_742_n142;
  tri   P2_lt_742_n141;
  tri   P2_lt_742_n140;
  tri   P2_lt_742_n139;
  tri   P2_lt_742_n138;
  tri   P2_lt_742_n137;
  tri   P2_lt_742_n136;
  tri   P2_lt_742_n135;
  tri   P2_lt_742_n134;
  tri   P2_lt_742_n133;
  tri   P2_lt_742_n132;
  tri   P2_lt_742_n131;
  tri   P2_lt_742_n130;
  tri   P2_lt_742_n129;
  tri   P2_lt_742_n128;
  tri   P2_lt_742_n127;
  tri   P2_lt_742_n126;
  tri   P2_lt_742_n125;
  tri   P2_lt_742_n124;
  tri   P2_lt_742_n123;
  tri   P2_lt_742_n122;
  tri   P2_lt_742_n121;
  tri   P2_lt_742_n120;
  tri   P2_lt_742_n119;
  tri   P2_lt_742_n118;
  tri   P2_lt_742_n117;
  tri   P2_lt_742_n116;
  tri   P2_lt_742_n115;
  tri   P2_lt_742_n114;
  tri   P2_lt_742_n113;
  tri   P2_lt_742_n112;
  tri   P2_lt_742_n110;
  tri   P2_lt_742_n109;
  tri   P2_lt_742_n108;
  tri   P2_lt_742_n107;
  tri   P2_lt_742_n106;
  tri   P2_lt_742_n105;
  tri   P2_lt_742_n104;
  tri   P2_lt_742_n103;
  tri   P2_lt_742_n102;
  tri   P2_lt_742_n101;
  tri   P2_lt_742_n100;
  tri   P2_lt_742_n99;
  tri   P2_lt_742_n98;
  tri   P2_lt_742_n97;
  tri   P2_lt_742_n96;
  tri   P2_lt_742_n95;
  tri   P2_lt_742_n94;
  tri   P2_lt_742_n93;
  tri   P2_lt_742_n92;
  tri   P2_lt_742_n91;
  tri   P2_lt_742_n90;
  tri   P2_lt_742_n89;
  tri   P2_lt_742_n88;
  tri   P2_lt_742_n87;
  tri   P2_lt_742_n86;
  tri   P2_lt_742_n85;
  tri   P2_lt_742_n84;
  tri   P2_lt_742_n83;
  tri   P2_lt_742_n82;
  tri   P2_lt_742_n81;
  tri   P2_lt_742_n80;
  tri   P2_lt_742_n79;
  tri   P2_lt_742_n78;
  tri   P2_lt_742_n77;
  tri   P2_lt_742_n76;
  tri   P2_lt_742_n75;
  tri   P2_lt_742_n74;
  tri   P2_lt_742_n73;
  tri   P2_lt_742_n72;
  tri   P2_lt_742_n71;
  tri   P2_lt_742_n69;
  tri   P2_lt_742_n1;
  tri   P2_lt_742_n5;
  tri   P2_lt_742_n14;
  tri   P2_lt_742_n13;
  tri   P2_lt_742_n24;
  tri   P2_lt_742_n23;
  tri   P2_lt_742_n34;
  tri   P2_lt_742_n33;
  tri   P2_add_918_n90;
  tri   P2_add_918_n89;
  tri   P2_add_918_n88;
  tri   P2_add_918_n86;
  tri   P2_add_918_n85;
  tri   P2_add_918_n84;
  tri   P2_add_918_n82;
  tri   P2_add_918_n81;
  tri   P2_add_918_n80;
  tri   P2_add_918_n79;
  tri   P2_add_918_n78;
  tri   P2_add_918_n77;
  tri   P2_add_918_n76;
  tri   P2_add_918_n75;
  tri   P2_add_918_n74;
  tri   P2_add_918_n72;
  tri   P2_add_918_n71;
  tri   P2_add_918_n70;
  tri   P2_add_918_n69;
  tri   P2_add_918_n68;
  tri   P2_add_918_n66;
  tri   P2_add_918_n65;
  tri   P2_add_918_n64;
  tri   P2_add_918_n63;
  tri   P2_add_918_n62;
  tri   P2_add_918_n61;
  tri   P2_add_918_n60;
  tri   P2_add_918_n59;
  tri   P2_add_918_n58;
  tri   P2_add_918_n57;
  tri   P2_add_918_n55;
  tri   P2_add_918_n54;
  tri   P2_add_918_n53;
  tri   P2_add_918_n51;
  tri   P2_add_918_n50;
  tri   P2_add_918_n48;
  tri   P2_add_918_n47;
  tri   P2_add_918_n46;
  tri   P2_add_918_n44;
  tri   P2_add_918_n43;
  tri   P2_add_918_n41;
  tri   P2_add_918_n40;
  tri   P2_add_918_n39;
  tri   P2_add_918_n37;
  tri   P2_add_918_n36;
  tri   P2_add_918_n34;
  tri   P2_add_918_n33;
  tri   P2_add_918_n32;
  tri   P2_add_918_n30;
  tri   P2_add_918_n29;
  tri   P2_add_918_n27;
  tri   P2_add_918_n26;
  tri   P2_add_918_n25;
  tri   P2_add_918_n23;
  tri   P2_add_918_n22;
  tri   P2_add_918_n20;
  tri   P2_add_918_n19;
  tri   P2_add_918_n18;
  tri   P2_add_918_n16;
  tri   P2_add_918_n15;
  tri   P2_add_918_n13;
  tri   P2_add_918_n12;
  tri   P2_add_918_n11;
  tri   P2_add_918_n9;
  tri   P2_add_918_n8;
  tri   P2_add_918_n6;
  tri   P2_add_918_n5;
  tri   P2_add_918_n4;
  tri   P2_add_918_n2;
  tri   P2_add_918_n1;
  tri   P2_add_918_n176;
  tri   P2_add_918_n175;
  tri   P2_add_918_n173;
  tri   P2_add_918_n172;
  tri   P2_add_918_n171;
  tri   P2_add_918_n169;
  tri   P2_add_918_n168;
  tri   P2_add_918_n167;
  tri   P2_add_918_n166;
  tri   P2_add_918_n165;
  tri   P2_add_918_n164;
  tri   P2_add_918_n163;
  tri   P2_add_918_n162;
  tri   P2_add_918_n161;
  tri   P2_add_918_n159;
  tri   P2_add_918_n158;
  tri   P2_add_918_n157;
  tri   P2_add_918_n156;
  tri   P2_add_918_n155;
  tri   P2_add_918_n153;
  tri   P2_add_918_n152;
  tri   P2_add_918_n150;
  tri   P2_add_918_n149;
  tri   P2_add_918_n148;
  tri   P2_add_918_n147;
  tri   P2_add_918_n146;
  tri   P2_add_918_n145;
  tri   P2_add_918_n144;
  tri   P2_add_918_n142;
  tri   P2_add_918_n141;
  tri   P2_add_918_n140;
  tri   P2_add_918_n139;
  tri   P2_add_918_n138;
  tri   P2_add_918_n137;
  tri   P2_add_918_n136;
  tri   P2_add_918_n135;
  tri   P2_add_918_n134;
  tri   P2_add_918_n132;
  tri   P2_add_918_n131;
  tri   P2_add_918_n130;
  tri   P2_add_918_n129;
  tri   P2_add_918_n128;
  tri   P2_add_918_n127;
  tri   P2_add_918_n126;
  tri   P2_add_918_n125;
  tri   P2_add_918_n124;
  tri   P2_add_918_n122;
  tri   P2_add_918_n121;
  tri   P2_add_918_n120;
  tri   P2_add_918_n119;
  tri   P2_add_918_n118;
  tri   P2_add_918_n117;
  tri   P2_add_918_n116;
  tri   P2_add_918_n115;
  tri   P2_add_918_n114;
  tri   P2_add_918_n112;
  tri   P2_add_918_n111;
  tri   P2_add_918_n110;
  tri   P2_add_918_n109;
  tri   P2_add_918_n108;
  tri   P2_add_918_n107;
  tri   P2_add_918_n106;
  tri   P2_add_918_n105;
  tri   P2_add_918_n104;
  tri   P2_add_918_n102;
  tri   P2_add_918_n101;
  tri   P2_add_918_n100;
  tri   P2_add_918_n99;
  tri   P2_add_918_n98;
  tri   P2_add_918_n97;
  tri   P2_add_918_n96;
  tri   P2_add_918_n87;
  tri   P2_add_918_n95;
  tri   P2_add_918_n94;
  tri   P2_add_918_n91;
  tri   P2_add_918_n92;
  tri   P2_add_918_n259;
  tri   P2_add_918_n258;
  tri   P2_add_918_n257;
  tri   P2_add_918_n10;
  tri   P2_add_918_n256;
  tri   P2_add_918_n255;
  tri   P2_add_918_n254;
  tri   P2_add_918_n3;
  tri   P2_add_918_n253;
  tri   P2_add_918_n252;
  tri   P2_add_918_n251;
  tri   P2_add_918_n249;
  tri   P2_add_918_n248;
  tri   P2_add_918_n247;
  tri   P2_add_918_n246;
  tri   P2_add_918_n245;
  tri   P2_add_918_n244;
  tri   P2_add_918_n243;
  tri   P2_add_918_n242;
  tri   P2_add_918_n241;
  tri   P2_add_918_n239;
  tri   P2_add_918_n238;
  tri   P2_add_918_n237;
  tri   P2_add_918_n236;
  tri   P2_add_918_n235;
  tri   P2_add_918_n234;
  tri   P2_add_918_n233;
  tri   P2_add_918_n232;
  tri   P2_add_918_n231;
  tri   P2_add_918_n229;
  tri   P2_add_918_n228;
  tri   P2_add_918_n227;
  tri   P2_add_918_n226;
  tri   P2_add_918_n225;
  tri   P2_add_918_n224;
  tri   P2_add_918_n223;
  tri   P2_add_918_n222;
  tri   P2_add_918_n221;
  tri   P2_add_918_n219;
  tri   P2_add_918_n218;
  tri   P2_add_918_n217;
  tri   P2_add_918_n216;
  tri   P2_add_918_n215;
  tri   P2_add_918_n214;
  tri   P2_add_918_n213;
  tri   P2_add_918_n212;
  tri   P2_add_918_n211;
  tri   P2_add_918_n209;
  tri   P2_add_918_n208;
  tri   P2_add_918_n207;
  tri   P2_add_918_n206;
  tri   P2_add_918_n205;
  tri   P2_add_918_n204;
  tri   P2_add_918_n203;
  tri   P2_add_918_n202;
  tri   P2_add_918_n201;
  tri   P2_add_918_n199;
  tri   P2_add_918_n198;
  tri   P2_add_918_n197;
  tri   P2_add_918_n196;
  tri   P2_add_918_n195;
  tri   P2_add_918_n194;
  tri   P2_add_918_n193;
  tri   P2_add_918_n192;
  tri   P2_add_918_n191;
  tri   P2_add_918_n189;
  tri   P2_add_918_n188;
  tri   P2_add_918_n187;
  tri   P2_add_918_n186;
  tri   P2_add_918_n185;
  tri   P2_add_918_n184;
  tri   P2_add_918_n183;
  tri   P2_add_918_n174;
  tri   P2_add_918_n182;
  tri   P2_add_918_n181;
  tri   P2_add_918_n177;
  tri   P2_add_918_n179;
  tri   P2_add_918_n178;
  tri   P2_add_918_n279;
  tri   P2_add_918_n278;
  tri   P2_add_918_n151;
  tri   P2_add_918_n277;
  tri   P2_add_918_n276;
  tri   P2_add_918_n275;
  tri   P2_add_918_n52;
  tri   P2_add_918_n274;
  tri   P2_add_918_n273;
  tri   P2_add_918_n272;
  tri   P2_add_918_n45;
  tri   P2_add_918_n271;
  tri   P2_add_918_n270;
  tri   P2_add_918_n269;
  tri   P2_add_918_n38;
  tri   P2_add_918_n268;
  tri   P2_add_918_n267;
  tri   P2_add_918_n266;
  tri   P2_add_918_n31;
  tri   P2_add_918_n265;
  tri   P2_add_918_n264;
  tri   P2_add_918_n263;
  tri   P2_add_918_n24;
  tri   P2_add_918_n262;
  tri   P2_add_918_n17;
  tri   P2_add_918_n261;
  tri   P2_add_918_n260;
  tri   P2_sub_938_n34;
  tri   P2_sub_938_n33;
  tri   P2_sub_938_n31;
  tri   P2_sub_938_n30;
  tri   P2_sub_938_n29;
  tri   P2_sub_938_n27;
  tri   P2_sub_938_n26;
  tri   P2_sub_938_n24;
  tri   P2_sub_938_n23;
  tri   P2_sub_938_n22;
  tri   P2_sub_938_n20;
  tri   P2_sub_938_n19;
  tri   P2_sub_938_n17;
  tri   P2_sub_938_n16;
  tri   P2_sub_938_n15;
  tri   P2_sub_938_n13;
  tri   P2_sub_938_n12;
  tri   P2_sub_938_n10;
  tri   P2_sub_938_n9;
  tri   P2_sub_938_n8;
  tri   P2_sub_938_n6;
  tri   P2_sub_938_n5;
  tri   P2_sub_938_n3;
  tri   P2_sub_938_n2;
  tri   P2_sub_938_n1;
  tri   P2_sub_938_n128;
  tri   P2_sub_938_n127;
  tri   P2_sub_938_n124;
  tri   P2_sub_938_n123;
  tri   P2_sub_938_n122;
  tri   P2_sub_938_n121;
  tri   P2_sub_938_n120;
  tri   P2_sub_938_n119;
  tri   P2_sub_938_n118;
  tri   P2_sub_938_n117;
  tri   P2_sub_938_n116;
  tri   P2_sub_938_n114;
  tri   P2_sub_938_n113;
  tri   P2_sub_938_n112;
  tri   P2_sub_938_n111;
  tri   P2_sub_938_n110;
  tri   P2_sub_938_n109;
  tri   P2_sub_938_n108;
  tri   P2_sub_938_n107;
  tri   P2_sub_938_n106;
  tri   P2_sub_938_n105;
  tri   P2_sub_938_n104;
  tri   P2_sub_938_n103;
  tri   P2_sub_938_n102;
  tri   P2_sub_938_n101;
  tri   P2_sub_938_n100;
  tri   P2_sub_938_n99;
  tri   P2_sub_938_n98;
  tri   P2_sub_938_n97;
  tri   P2_sub_938_n96;
  tri   P2_sub_938_n95;
  tri   P2_sub_938_n94;
  tri   P2_sub_938_n93;
  tri   P2_sub_938_n92;
  tri   P2_sub_938_n91;
  tri   P2_sub_938_n90;
  tri   P2_sub_938_n89;
  tri   P2_sub_938_n88;
  tri   P2_sub_938_n87;
  tri   P2_sub_938_n86;
  tri   P2_sub_938_n85;
  tri   P2_sub_938_n84;
  tri   P2_sub_938_n83;
  tri   P2_sub_938_n82;
  tri   P2_sub_938_n81;
  tri   P2_sub_938_n80;
  tri   P2_sub_938_n79;
  tri   P2_sub_938_n78;
  tri   P2_sub_938_n77;
  tri   P2_sub_938_n76;
  tri   P2_sub_938_n75;
  tri   P2_sub_938_n74;
  tri   P2_sub_938_n73;
  tri   P2_sub_938_n72;
  tri   P2_sub_938_n71;
  tri   P2_sub_938_n70;
  tri   P2_sub_938_n69;
  tri   P2_sub_938_n67;
  tri   P2_sub_938_n66;
  tri   P2_sub_938_n65;
  tri   P2_sub_938_n64;
  tri   P2_sub_938_n63;
  tri   P2_sub_938_n62;
  tri   P2_sub_938_n61;
  tri   P2_sub_938_n59;
  tri   P2_sub_938_n60;
  tri   P2_sub_938_n58;
  tri   P2_sub_938_n57;
  tri   P2_sub_938_n55;
  tri   P2_sub_938_n54;
  tri   P2_sub_938_n52;
  tri   P2_sub_938_n51;
  tri   P2_sub_938_n50;
  tri   P2_sub_938_n48;
  tri   P2_sub_938_n47;
  tri   P2_sub_938_n45;
  tri   P2_sub_938_n44;
  tri   P2_sub_938_n43;
  tri   P2_sub_938_n41;
  tri   P2_sub_938_n40;
  tri   P2_sub_938_n36;
  tri   P2_sub_938_n37;
  tri   P2_sub_938_n38;
  tri   P2_sub_938_n216;
  tri   P2_sub_938_n212;
  tri   P2_sub_938_n211;
  tri   P2_sub_938_n210;
  tri   P2_sub_938_n209;
  tri   P2_sub_938_n208;
  tri   P2_sub_938_n207;
  tri   P2_sub_938_n206;
  tri   P2_sub_938_n205;
  tri   P2_sub_938_n204;
  tri   P2_sub_938_n202;
  tri   P2_sub_938_n201;
  tri   P2_sub_938_n200;
  tri   P2_sub_938_n199;
  tri   P2_sub_938_n198;
  tri   P2_sub_938_n197;
  tri   P2_sub_938_n196;
  tri   P2_sub_938_n195;
  tri   P2_sub_938_n194;
  tri   P2_sub_938_n193;
  tri   P2_sub_938_n192;
  tri   P2_sub_938_n191;
  tri   P2_sub_938_n190;
  tri   P2_sub_938_n189;
  tri   P2_sub_938_n188;
  tri   P2_sub_938_n187;
  tri   P2_sub_938_n186;
  tri   P2_sub_938_n185;
  tri   P2_sub_938_n184;
  tri   P2_sub_938_n183;
  tri   P2_sub_938_n182;
  tri   P2_sub_938_n181;
  tri   P2_sub_938_n180;
  tri   P2_sub_938_n179;
  tri   P2_sub_938_n178;
  tri   P2_sub_938_n177;
  tri   P2_sub_938_n176;
  tri   P2_sub_938_n175;
  tri   P2_sub_938_n174;
  tri   P2_sub_938_n173;
  tri   P2_sub_938_n172;
  tri   P2_sub_938_n171;
  tri   P2_sub_938_n170;
  tri   P2_sub_938_n169;
  tri   P2_sub_938_n168;
  tri   P2_sub_938_n167;
  tri   P2_sub_938_n166;
  tri   P2_sub_938_n165;
  tri   P2_sub_938_n164;
  tri   P2_sub_938_n163;
  tri   P2_sub_938_n162;
  tri   P2_sub_938_n161;
  tri   P2_sub_938_n160;
  tri   P2_sub_938_n159;
  tri   P2_sub_938_n158;
  tri   P2_sub_938_n157;
  tri   P2_sub_938_n154;
  tri   P2_sub_938_n153;
  tri   P2_sub_938_n151;
  tri   P2_sub_938_n150;
  tri   P2_sub_938_n149;
  tri   P2_sub_938_n148;
  tri   P2_sub_938_n147;
  tri   P2_sub_938_n146;
  tri   P2_sub_938_n145;
  tri   P2_sub_938_n144;
  tri   P2_sub_938_n143;
  tri   P2_sub_938_n142;
  tri   P2_sub_938_n141;
  tri   P2_sub_938_n140;
  tri   P2_sub_938_n139;
  tri   P2_sub_938_n125;
  tri   P2_sub_938_n138;
  tri   P2_sub_938_n137;
  tri   P2_sub_938_n136;
  tri   P2_sub_938_n135;
  tri   P2_sub_938_n134;
  tri   P2_sub_938_n133;
  tri   P2_sub_938_n132;
  tri   P2_sub_938_n131;
  tri   P2_sub_938_n126;
  tri   P2_sub_938_n130;
  tri   P2_sub_938_n129;
  tri   P2_sub_938_n115;
  tri   P2_sub_938_n281;
  tri   P2_sub_938_n280;
  tri   P2_sub_938_n279;
  tri   P2_sub_938_n278;
  tri   P2_sub_938_n152;
  tri   P2_sub_938_n277;
  tri   P2_sub_938_n156;
  tri   P2_sub_938_n276;
  tri   P2_sub_938_n275;
  tri   P2_sub_938_n274;
  tri   P2_sub_938_n53;
  tri   P2_sub_938_n56;
  tri   P2_sub_938_n273;
  tri   P2_sub_938_n272;
  tri   P2_sub_938_n271;
  tri   P2_sub_938_n46;
  tri   P2_sub_938_n49;
  tri   P2_sub_938_n270;
  tri   P2_sub_938_n269;
  tri   P2_sub_938_n268;
  tri   P2_sub_938_n39;
  tri   P2_sub_938_n42;
  tri   P2_sub_938_n267;
  tri   P2_sub_938_n266;
  tri   P2_sub_938_n265;
  tri   P2_sub_938_n32;
  tri   P2_sub_938_n35;
  tri   P2_sub_938_n264;
  tri   P2_sub_938_n263;
  tri   P2_sub_938_n262;
  tri   P2_sub_938_n25;
  tri   P2_sub_938_n28;
  tri   P2_sub_938_n261;
  tri   P2_sub_938_n260;
  tri   P2_sub_938_n259;
  tri   P2_sub_938_n18;
  tri   P2_sub_938_n21;
  tri   P2_sub_938_n258;
  tri   P2_sub_938_n257;
  tri   P2_sub_938_n256;
  tri   P2_sub_938_n11;
  tri   P2_sub_938_n14;
  tri   P2_sub_938_n255;
  tri   P2_sub_938_n254;
  tri   P2_sub_938_n253;
  tri   P2_sub_938_n4;
  tri   P2_sub_938_n7;
  tri   P2_sub_938_n252;
  tri   P2_sub_938_n251;
  tri   P2_sub_938_n250;
  tri   P2_sub_938_n249;
  tri   P2_sub_938_n248;
  tri   P2_sub_938_n247;
  tri   P2_sub_938_n246;
  tri   P2_sub_938_n245;
  tri   P2_sub_938_n244;
  tri   P2_sub_938_n243;
  tri   P2_sub_938_n242;
  tri   P2_sub_938_n241;
  tri   P2_sub_938_n240;
  tri   P2_sub_938_n239;
  tri   P2_sub_938_n238;
  tri   P2_sub_938_n237;
  tri   P2_sub_938_n236;
  tri   P2_sub_938_n235;
  tri   P2_sub_938_n234;
  tri   P2_sub_938_n233;
  tri   P2_sub_938_n232;
  tri   P2_sub_938_n231;
  tri   P2_sub_938_n230;
  tri   P2_sub_938_n229;
  tri   P2_sub_938_n228;
  tri   P2_sub_938_n227;
  tri   P2_sub_938_n213;
  tri   P2_sub_938_n226;
  tri   P2_sub_938_n225;
  tri   P2_sub_938_n224;
  tri   P2_sub_938_n223;
  tri   P2_sub_938_n222;
  tri   P2_sub_938_n221;
  tri   P2_sub_938_n220;
  tri   P2_sub_938_n219;
  tri   P2_sub_938_n214;
  tri   P2_sub_938_n218;
  tri   P2_sub_938_n217;
  tri   P2_sub_938_n215;
  tri   P2_sub_938_n203;
  tri   P2_add_958_n62;
  tri   P2_add_958_n59;
  tri   P2_add_958_n58;
  tri   P2_add_958_n57;
  tri   P2_add_958_n55;
  tri   P2_add_958_n54;
  tri   P2_add_958_n53;
  tri   P2_add_958_n51;
  tri   P2_add_958_n50;
  tri   P2_add_958_n48;
  tri   P2_add_958_n47;
  tri   P2_add_958_n46;
  tri   P2_add_958_n44;
  tri   P2_add_958_n43;
  tri   P2_add_958_n41;
  tri   P2_add_958_n40;
  tri   P2_add_958_n39;
  tri   P2_add_958_n37;
  tri   P2_add_958_n36;
  tri   P2_add_958_n34;
  tri   P2_add_958_n33;
  tri   P2_add_958_n32;
  tri   P2_add_958_n30;
  tri   P2_add_958_n29;
  tri   P2_add_958_n27;
  tri   P2_add_958_n26;
  tri   P2_add_958_n25;
  tri   P2_add_958_n23;
  tri   P2_add_958_n22;
  tri   P2_add_958_n20;
  tri   P2_add_958_n19;
  tri   P2_add_958_n18;
  tri   P2_add_958_n16;
  tri   P2_add_958_n15;
  tri   P2_add_958_n13;
  tri   P2_add_958_n12;
  tri   P2_add_958_n11;
  tri   P2_add_958_n9;
  tri   P2_add_958_n8;
  tri   P2_add_958_n6;
  tri   P2_add_958_n5;
  tri   P2_add_958_n4;
  tri   P2_add_958_n2;
  tri   P2_add_958_n1;
  tri   P2_add_958_n146;
  tri   P2_add_958_n145;
  tri   P2_add_958_n142;
  tri   P2_add_958_n141;
  tri   P2_add_958_n140;
  tri   P2_add_958_n139;
  tri   P2_add_958_n138;
  tri   P2_add_958_n137;
  tri   P2_add_958_n136;
  tri   P2_add_958_n135;
  tri   P2_add_958_n134;
  tri   P2_add_958_n132;
  tri   P2_add_958_n131;
  tri   P2_add_958_n130;
  tri   P2_add_958_n129;
  tri   P2_add_958_n128;
  tri   P2_add_958_n127;
  tri   P2_add_958_n126;
  tri   P2_add_958_n125;
  tri   P2_add_958_n124;
  tri   P2_add_958_n122;
  tri   P2_add_958_n121;
  tri   P2_add_958_n120;
  tri   P2_add_958_n119;
  tri   P2_add_958_n118;
  tri   P2_add_958_n117;
  tri   P2_add_958_n116;
  tri   P2_add_958_n115;
  tri   P2_add_958_n114;
  tri   P2_add_958_n112;
  tri   P2_add_958_n111;
  tri   P2_add_958_n110;
  tri   P2_add_958_n109;
  tri   P2_add_958_n108;
  tri   P2_add_958_n107;
  tri   P2_add_958_n106;
  tri   P2_add_958_n105;
  tri   P2_add_958_n104;
  tri   P2_add_958_n102;
  tri   P2_add_958_n101;
  tri   P2_add_958_n100;
  tri   P2_add_958_n99;
  tri   P2_add_958_n98;
  tri   P2_add_958_n97;
  tri   P2_add_958_n96;
  tri   P2_add_958_n95;
  tri   P2_add_958_n94;
  tri   P2_add_958_n92;
  tri   P2_add_958_n91;
  tri   P2_add_958_n90;
  tri   P2_add_958_n89;
  tri   P2_add_958_n88;
  tri   P2_add_958_n87;
  tri   P2_add_958_n86;
  tri   P2_add_958_n85;
  tri   P2_add_958_n84;
  tri   P2_add_958_n82;
  tri   P2_add_958_n81;
  tri   P2_add_958_n80;
  tri   P2_add_958_n79;
  tri   P2_add_958_n78;
  tri   P2_add_958_n77;
  tri   P2_add_958_n76;
  tri   P2_add_958_n75;
  tri   P2_add_958_n74;
  tri   P2_add_958_n72;
  tri   P2_add_958_n71;
  tri   P2_add_958_n70;
  tri   P2_add_958_n69;
  tri   P2_add_958_n68;
  tri   P2_add_958_n60;
  tri   P2_add_958_n66;
  tri   P2_add_958_n65;
  tri   P2_add_958_n61;
  tri   P2_add_958_n63;
  tri   P2_add_958_n64;
  tri   P2_add_958_n232;
  tri   P2_add_958_n229;
  tri   P2_add_958_n228;
  tri   P2_add_958_n227;
  tri   P2_add_958_n226;
  tri   P2_add_958_n225;
  tri   P2_add_958_n224;
  tri   P2_add_958_n223;
  tri   P2_add_958_n222;
  tri   P2_add_958_n221;
  tri   P2_add_958_n219;
  tri   P2_add_958_n218;
  tri   P2_add_958_n217;
  tri   P2_add_958_n216;
  tri   P2_add_958_n215;
  tri   P2_add_958_n214;
  tri   P2_add_958_n213;
  tri   P2_add_958_n212;
  tri   P2_add_958_n211;
  tri   P2_add_958_n209;
  tri   P2_add_958_n208;
  tri   P2_add_958_n207;
  tri   P2_add_958_n206;
  tri   P2_add_958_n205;
  tri   P2_add_958_n204;
  tri   P2_add_958_n203;
  tri   P2_add_958_n202;
  tri   P2_add_958_n201;
  tri   P2_add_958_n199;
  tri   P2_add_958_n198;
  tri   P2_add_958_n197;
  tri   P2_add_958_n196;
  tri   P2_add_958_n195;
  tri   P2_add_958_n194;
  tri   P2_add_958_n193;
  tri   P2_add_958_n192;
  tri   P2_add_958_n191;
  tri   P2_add_958_n189;
  tri   P2_add_958_n188;
  tri   P2_add_958_n187;
  tri   P2_add_958_n186;
  tri   P2_add_958_n185;
  tri   P2_add_958_n184;
  tri   P2_add_958_n183;
  tri   P2_add_958_n182;
  tri   P2_add_958_n181;
  tri   P2_add_958_n179;
  tri   P2_add_958_n178;
  tri   P2_add_958_n177;
  tri   P2_add_958_n176;
  tri   P2_add_958_n175;
  tri   P2_add_958_n174;
  tri   P2_add_958_n173;
  tri   P2_add_958_n172;
  tri   P2_add_958_n171;
  tri   P2_add_958_n169;
  tri   P2_add_958_n168;
  tri   P2_add_958_n167;
  tri   P2_add_958_n166;
  tri   P2_add_958_n165;
  tri   P2_add_958_n164;
  tri   P2_add_958_n163;
  tri   P2_add_958_n162;
  tri   P2_add_958_n161;
  tri   P2_add_958_n159;
  tri   P2_add_958_n158;
  tri   P2_add_958_n157;
  tri   P2_add_958_n156;
  tri   P2_add_958_n155;
  tri   P2_add_958_n153;
  tri   P2_add_958_n152;
  tri   P2_add_958_n150;
  tri   P2_add_958_n149;
  tri   P2_add_958_n148;
  tri   P2_add_958_n144;
  tri   P2_add_958_n147;
  tri   P2_add_958_n279;
  tri   P2_add_958_n278;
  tri   P2_add_958_n151;
  tri   P2_add_958_n277;
  tri   P2_add_958_n276;
  tri   P2_add_958_n275;
  tri   P2_add_958_n52;
  tri   P2_add_958_n274;
  tri   P2_add_958_n273;
  tri   P2_add_958_n272;
  tri   P2_add_958_n45;
  tri   P2_add_958_n271;
  tri   P2_add_958_n270;
  tri   P2_add_958_n269;
  tri   P2_add_958_n38;
  tri   P2_add_958_n268;
  tri   P2_add_958_n267;
  tri   P2_add_958_n266;
  tri   P2_add_958_n31;
  tri   P2_add_958_n265;
  tri   P2_add_958_n264;
  tri   P2_add_958_n263;
  tri   P2_add_958_n24;
  tri   P2_add_958_n262;
  tri   P2_add_958_n261;
  tri   P2_add_958_n260;
  tri   P2_add_958_n17;
  tri   P2_add_958_n259;
  tri   P2_add_958_n258;
  tri   P2_add_958_n257;
  tri   P2_add_958_n10;
  tri   P2_add_958_n256;
  tri   P2_add_958_n255;
  tri   P2_add_958_n254;
  tri   P2_add_958_n3;
  tri   P2_add_958_n253;
  tri   P2_add_958_n252;
  tri   P2_add_958_n251;
  tri   P2_add_958_n249;
  tri   P2_add_958_n248;
  tri   P2_add_958_n247;
  tri   P2_add_958_n246;
  tri   P2_add_958_n245;
  tri   P2_add_958_n244;
  tri   P2_add_958_n243;
  tri   P2_add_958_n242;
  tri   P2_add_958_n241;
  tri   P2_add_958_n239;
  tri   P2_add_958_n238;
  tri   P2_add_958_n237;
  tri   P2_add_958_n236;
  tri   P2_add_958_n235;
  tri   P2_add_958_n231;
  tri   P2_add_958_n233;
  tri   P2_add_958_n234;
  tri   P2_sub_978_n98;
  tri   P2_sub_978_n97;
  tri   P2_sub_978_n94;
  tri   P2_sub_978_n93;
  tri   P2_sub_978_n92;
  tri   P2_sub_978_n91;
  tri   P2_sub_978_n90;
  tri   P2_sub_978_n89;
  tri   P2_sub_978_n88;
  tri   P2_sub_978_n87;
  tri   P2_sub_978_n86;
  tri   P2_sub_978_n85;
  tri   P2_sub_978_n84;
  tri   P2_sub_978_n83;
  tri   P2_sub_978_n82;
  tri   P2_sub_978_n81;
  tri   P2_sub_978_n80;
  tri   P2_sub_978_n79;
  tri   P2_sub_978_n78;
  tri   P2_sub_978_n77;
  tri   P2_sub_978_n76;
  tri   P2_sub_978_n75;
  tri   P2_sub_978_n74;
  tri   P2_sub_978_n73;
  tri   P2_sub_978_n72;
  tri   P2_sub_978_n71;
  tri   P2_sub_978_n70;
  tri   P2_sub_978_n69;
  tri   P2_sub_978_n67;
  tri   P2_sub_978_n66;
  tri   P2_sub_978_n65;
  tri   P2_sub_978_n64;
  tri   P2_sub_978_n63;
  tri   P2_sub_978_n62;
  tri   P2_sub_978_n61;
  tri   P2_sub_978_n59;
  tri   P2_sub_978_n60;
  tri   P2_sub_978_n58;
  tri   P2_sub_978_n57;
  tri   P2_sub_978_n55;
  tri   P2_sub_978_n54;
  tri   P2_sub_978_n52;
  tri   P2_sub_978_n51;
  tri   P2_sub_978_n50;
  tri   P2_sub_978_n48;
  tri   P2_sub_978_n47;
  tri   P2_sub_978_n45;
  tri   P2_sub_978_n44;
  tri   P2_sub_978_n43;
  tri   P2_sub_978_n41;
  tri   P2_sub_978_n40;
  tri   P2_sub_978_n38;
  tri   P2_sub_978_n37;
  tri   P2_sub_978_n36;
  tri   P2_sub_978_n34;
  tri   P2_sub_978_n33;
  tri   P2_sub_978_n31;
  tri   P2_sub_978_n30;
  tri   P2_sub_978_n29;
  tri   P2_sub_978_n27;
  tri   P2_sub_978_n26;
  tri   P2_sub_978_n24;
  tri   P2_sub_978_n23;
  tri   P2_sub_978_n22;
  tri   P2_sub_978_n20;
  tri   P2_sub_978_n19;
  tri   P2_sub_978_n17;
  tri   P2_sub_978_n16;
  tri   P2_sub_978_n15;
  tri   P2_sub_978_n13;
  tri   P2_sub_978_n12;
  tri   P2_sub_978_n10;
  tri   P2_sub_978_n9;
  tri   P2_sub_978_n8;
  tri   P2_sub_978_n6;
  tri   P2_sub_978_n5;
  tri   P2_sub_978_n3;
  tri   P2_sub_978_n2;
  tri   P2_sub_978_n1;
  tri   P2_sub_978_n186;
  tri   P2_sub_978_n185;
  tri   P2_sub_978_n182;
  tri   P2_sub_978_n181;
  tri   P2_sub_978_n180;
  tri   P2_sub_978_n179;
  tri   P2_sub_978_n178;
  tri   P2_sub_978_n177;
  tri   P2_sub_978_n176;
  tri   P2_sub_978_n175;
  tri   P2_sub_978_n174;
  tri   P2_sub_978_n172;
  tri   P2_sub_978_n171;
  tri   P2_sub_978_n170;
  tri   P2_sub_978_n169;
  tri   P2_sub_978_n168;
  tri   P2_sub_978_n167;
  tri   P2_sub_978_n166;
  tri   P2_sub_978_n165;
  tri   P2_sub_978_n164;
  tri   P2_sub_978_n163;
  tri   P2_sub_978_n162;
  tri   P2_sub_978_n161;
  tri   P2_sub_978_n160;
  tri   P2_sub_978_n159;
  tri   P2_sub_978_n158;
  tri   P2_sub_978_n157;
  tri   P2_sub_978_n154;
  tri   P2_sub_978_n153;
  tri   P2_sub_978_n151;
  tri   P2_sub_978_n150;
  tri   P2_sub_978_n149;
  tri   P2_sub_978_n148;
  tri   P2_sub_978_n147;
  tri   P2_sub_978_n146;
  tri   P2_sub_978_n145;
  tri   P2_sub_978_n144;
  tri   P2_sub_978_n143;
  tri   P2_sub_978_n142;
  tri   P2_sub_978_n141;
  tri   P2_sub_978_n140;
  tri   P2_sub_978_n139;
  tri   P2_sub_978_n138;
  tri   P2_sub_978_n137;
  tri   P2_sub_978_n136;
  tri   P2_sub_978_n135;
  tri   P2_sub_978_n134;
  tri   P2_sub_978_n133;
  tri   P2_sub_978_n132;
  tri   P2_sub_978_n131;
  tri   P2_sub_978_n130;
  tri   P2_sub_978_n129;
  tri   P2_sub_978_n128;
  tri   P2_sub_978_n127;
  tri   P2_sub_978_n126;
  tri   P2_sub_978_n125;
  tri   P2_sub_978_n124;
  tri   P2_sub_978_n123;
  tri   P2_sub_978_n122;
  tri   P2_sub_978_n121;
  tri   P2_sub_978_n120;
  tri   P2_sub_978_n119;
  tri   P2_sub_978_n118;
  tri   P2_sub_978_n117;
  tri   P2_sub_978_n116;
  tri   P2_sub_978_n115;
  tri   P2_sub_978_n114;
  tri   P2_sub_978_n113;
  tri   P2_sub_978_n112;
  tri   P2_sub_978_n111;
  tri   P2_sub_978_n110;
  tri   P2_sub_978_n109;
  tri   P2_sub_978_n95;
  tri   P2_sub_978_n108;
  tri   P2_sub_978_n107;
  tri   P2_sub_978_n106;
  tri   P2_sub_978_n105;
  tri   P2_sub_978_n104;
  tri   P2_sub_978_n103;
  tri   P2_sub_978_n102;
  tri   P2_sub_978_n101;
  tri   P2_sub_978_n96;
  tri   P2_sub_978_n100;
  tri   P2_sub_978_n99;
  tri   P2_sub_978_n35;
  tri   P2_sub_978_n263;
  tri   P2_sub_978_n25;
  tri   P2_sub_978_n28;
  tri   P2_sub_978_n261;
  tri   P2_sub_978_n260;
  tri   P2_sub_978_n259;
  tri   P2_sub_978_n18;
  tri   P2_sub_978_n21;
  tri   P2_sub_978_n258;
  tri   P2_sub_978_n257;
  tri   P2_sub_978_n256;
  tri   P2_sub_978_n11;
  tri   P2_sub_978_n14;
  tri   P2_sub_978_n255;
  tri   P2_sub_978_n254;
  tri   P2_sub_978_n253;
  tri   P2_sub_978_n4;
  tri   P2_sub_978_n7;
  tri   P2_sub_978_n252;
  tri   P2_sub_978_n251;
  tri   P2_sub_978_n250;
  tri   P2_sub_978_n248;
  tri   P2_sub_978_n247;
  tri   P2_sub_978_n246;
  tri   P2_sub_978_n245;
  tri   P2_sub_978_n244;
  tri   P2_sub_978_n242;
  tri   P2_sub_978_n241;
  tri   P2_sub_978_n240;
  tri   P2_sub_978_n239;
  tri   P2_sub_978_n238;
  tri   P2_sub_978_n237;
  tri   P2_sub_978_n236;
  tri   P2_sub_978_n235;
  tri   P2_sub_978_n234;
  tri   P2_sub_978_n233;
  tri   P2_sub_978_n232;
  tri   P2_sub_978_n231;
  tri   P2_sub_978_n230;
  tri   P2_sub_978_n229;
  tri   P2_sub_978_n228;
  tri   P2_sub_978_n227;
  tri   P2_sub_978_n226;
  tri   P2_sub_978_n225;
  tri   P2_sub_978_n224;
  tri   P2_sub_978_n223;
  tri   P2_sub_978_n222;
  tri   P2_sub_978_n221;
  tri   P2_sub_978_n220;
  tri   P2_sub_978_n219;
  tri   P2_sub_978_n218;
  tri   P2_sub_978_n217;
  tri   P2_sub_978_n216;
  tri   P2_sub_978_n215;
  tri   P2_sub_978_n214;
  tri   P2_sub_978_n213;
  tri   P2_sub_978_n212;
  tri   P2_sub_978_n211;
  tri   P2_sub_978_n210;
  tri   P2_sub_978_n209;
  tri   P2_sub_978_n208;
  tri   P2_sub_978_n207;
  tri   P2_sub_978_n206;
  tri   P2_sub_978_n205;
  tri   P2_sub_978_n204;
  tri   P2_sub_978_n203;
  tri   P2_sub_978_n202;
  tri   P2_sub_978_n201;
  tri   P2_sub_978_n200;
  tri   P2_sub_978_n199;
  tri   P2_sub_978_n198;
  tri   P2_sub_978_n197;
  tri   P2_sub_978_n183;
  tri   P2_sub_978_n196;
  tri   P2_sub_978_n195;
  tri   P2_sub_978_n194;
  tri   P2_sub_978_n193;
  tri   P2_sub_978_n192;
  tri   P2_sub_978_n191;
  tri   P2_sub_978_n190;
  tri   P2_sub_978_n189;
  tri   P2_sub_978_n184;
  tri   P2_sub_978_n188;
  tri   P2_sub_978_n187;
  tri   P2_sub_978_n173;
  tri   P2_sub_978_n281;
  tri   P2_sub_978_n280;
  tri   P2_sub_978_n243;
  tri   P2_sub_978_n249;
  tri   P2_sub_978_n279;
  tri   P2_sub_978_n278;
  tri   P2_sub_978_n152;
  tri   P2_sub_978_n277;
  tri   P2_sub_978_n156;
  tri   P2_sub_978_n276;
  tri   P2_sub_978_n275;
  tri   P2_sub_978_n274;
  tri   P2_sub_978_n53;
  tri   P2_sub_978_n56;
  tri   P2_sub_978_n273;
  tri   P2_sub_978_n272;
  tri   P2_sub_978_n271;
  tri   P2_sub_978_n46;
  tri   P2_sub_978_n49;
  tri   P2_sub_978_n270;
  tri   P2_sub_978_n269;
  tri   P2_sub_978_n268;
  tri   P2_sub_978_n39;
  tri   P2_sub_978_n42;
  tri   P2_sub_978_n267;
  tri   P2_sub_978_n266;
  tri   P2_sub_978_n265;
  tri   P2_sub_978_n262;
  tri   P2_sub_978_n264;
  tri   P2_sub_978_n32;
  tri   P2_add_998_n27;
  tri   P2_add_998_n26;
  tri   P2_add_998_n25;
  tri   P2_add_998_n23;
  tri   P2_add_998_n22;
  tri   P2_add_998_n20;
  tri   P2_add_998_n19;
  tri   P2_add_998_n18;
  tri   P2_add_998_n16;
  tri   P2_add_998_n15;
  tri   P2_add_998_n13;
  tri   P2_add_998_n12;
  tri   P2_add_998_n11;
  tri   P2_add_998_n9;
  tri   P2_add_998_n8;
  tri   P2_add_998_n6;
  tri   P2_add_998_n5;
  tri   P2_add_998_n4;
  tri   P2_add_998_n2;
  tri   P2_add_998_n1;
  tri   P2_add_998_n116;
  tri   P2_add_998_n115;
  tri   P2_add_998_n114;
  tri   P2_add_998_n112;
  tri   P2_add_998_n111;
  tri   P2_add_998_n110;
  tri   P2_add_998_n109;
  tri   P2_add_998_n108;
  tri   P2_add_998_n107;
  tri   P2_add_998_n106;
  tri   P2_add_998_n105;
  tri   P2_add_998_n104;
  tri   P2_add_998_n102;
  tri   P2_add_998_n101;
  tri   P2_add_998_n100;
  tri   P2_add_998_n99;
  tri   P2_add_998_n98;
  tri   P2_add_998_n97;
  tri   P2_add_998_n96;
  tri   P2_add_998_n95;
  tri   P2_add_998_n94;
  tri   P2_add_998_n92;
  tri   P2_add_998_n91;
  tri   P2_add_998_n90;
  tri   P2_add_998_n89;
  tri   P2_add_998_n88;
  tri   P2_add_998_n87;
  tri   P2_add_998_n86;
  tri   P2_add_998_n85;
  tri   P2_add_998_n84;
  tri   P2_add_998_n82;
  tri   P2_add_998_n81;
  tri   P2_add_998_n80;
  tri   P2_add_998_n79;
  tri   P2_add_998_n78;
  tri   P2_add_998_n77;
  tri   P2_add_998_n76;
  tri   P2_add_998_n75;
  tri   P2_add_998_n74;
  tri   P2_add_998_n72;
  tri   P2_add_998_n71;
  tri   P2_add_998_n70;
  tri   P2_add_998_n69;
  tri   P2_add_998_n68;
  tri   P2_add_998_n66;
  tri   P2_add_998_n65;
  tri   P2_add_998_n64;
  tri   P2_add_998_n63;
  tri   P2_add_998_n62;
  tri   P2_add_998_n61;
  tri   P2_add_998_n60;
  tri   P2_add_998_n59;
  tri   P2_add_998_n58;
  tri   P2_add_998_n57;
  tri   P2_add_998_n55;
  tri   P2_add_998_n54;
  tri   P2_add_998_n53;
  tri   P2_add_998_n51;
  tri   P2_add_998_n50;
  tri   P2_add_998_n48;
  tri   P2_add_998_n47;
  tri   P2_add_998_n46;
  tri   P2_add_998_n44;
  tri   P2_add_998_n43;
  tri   P2_add_998_n41;
  tri   P2_add_998_n40;
  tri   P2_add_998_n39;
  tri   P2_add_998_n37;
  tri   P2_add_998_n36;
  tri   P2_add_998_n34;
  tri   P2_add_998_n33;
  tri   P2_add_998_n29;
  tri   P2_add_998_n30;
  tri   P2_add_998_n32;
  tri   P2_add_998_n203;
  tri   P2_add_998_n202;
  tri   P2_add_998_n199;
  tri   P2_add_998_n198;
  tri   P2_add_998_n197;
  tri   P2_add_998_n196;
  tri   P2_add_998_n195;
  tri   P2_add_998_n194;
  tri   P2_add_998_n193;
  tri   P2_add_998_n192;
  tri   P2_add_998_n191;
  tri   P2_add_998_n189;
  tri   P2_add_998_n188;
  tri   P2_add_998_n187;
  tri   P2_add_998_n186;
  tri   P2_add_998_n185;
  tri   P2_add_998_n184;
  tri   P2_add_998_n183;
  tri   P2_add_998_n182;
  tri   P2_add_998_n181;
  tri   P2_add_998_n179;
  tri   P2_add_998_n178;
  tri   P2_add_998_n177;
  tri   P2_add_998_n176;
  tri   P2_add_998_n175;
  tri   P2_add_998_n174;
  tri   P2_add_998_n173;
  tri   P2_add_998_n172;
  tri   P2_add_998_n171;
  tri   P2_add_998_n169;
  tri   P2_add_998_n168;
  tri   P2_add_998_n167;
  tri   P2_add_998_n166;
  tri   P2_add_998_n165;
  tri   P2_add_998_n164;
  tri   P2_add_998_n163;
  tri   P2_add_998_n162;
  tri   P2_add_998_n161;
  tri   P2_add_998_n159;
  tri   P2_add_998_n158;
  tri   P2_add_998_n157;
  tri   P2_add_998_n156;
  tri   P2_add_998_n155;
  tri   P2_add_998_n153;
  tri   P2_add_998_n152;
  tri   P2_add_998_n150;
  tri   P2_add_998_n149;
  tri   P2_add_998_n148;
  tri   P2_add_998_n147;
  tri   P2_add_998_n146;
  tri   P2_add_998_n145;
  tri   P2_add_998_n144;
  tri   P2_add_998_n142;
  tri   P2_add_998_n141;
  tri   P2_add_998_n140;
  tri   P2_add_998_n139;
  tri   P2_add_998_n138;
  tri   P2_add_998_n137;
  tri   P2_add_998_n136;
  tri   P2_add_998_n135;
  tri   P2_add_998_n134;
  tri   P2_add_998_n132;
  tri   P2_add_998_n131;
  tri   P2_add_998_n130;
  tri   P2_add_998_n129;
  tri   P2_add_998_n128;
  tri   P2_add_998_n127;
  tri   P2_add_998_n126;
  tri   P2_add_998_n125;
  tri   P2_add_998_n124;
  tri   P2_add_998_n122;
  tri   P2_add_998_n121;
  tri   P2_add_998_n120;
  tri   P2_add_998_n117;
  tri   P2_add_998_n119;
  tri   P2_add_998_n118;
  tri   P2_add_998_n279;
  tri   P2_add_998_n278;
  tri   P2_add_998_n151;
  tri   P2_add_998_n277;
  tri   P2_add_998_n276;
  tri   P2_add_998_n275;
  tri   P2_add_998_n52;
  tri   P2_add_998_n274;
  tri   P2_add_998_n273;
  tri   P2_add_998_n272;
  tri   P2_add_998_n45;
  tri   P2_add_998_n271;
  tri   P2_add_998_n270;
  tri   P2_add_998_n269;
  tri   P2_add_998_n38;
  tri   P2_add_998_n268;
  tri   P2_add_998_n267;
  tri   P2_add_998_n266;
  tri   P2_add_998_n31;
  tri   P2_add_998_n265;
  tri   P2_add_998_n264;
  tri   P2_add_998_n263;
  tri   P2_add_998_n24;
  tri   P2_add_998_n262;
  tri   P2_add_998_n261;
  tri   P2_add_998_n260;
  tri   P2_add_998_n17;
  tri   P2_add_998_n259;
  tri   P2_add_998_n258;
  tri   P2_add_998_n257;
  tri   P2_add_998_n10;
  tri   P2_add_998_n256;
  tri   P2_add_998_n255;
  tri   P2_add_998_n254;
  tri   P2_add_998_n3;
  tri   P2_add_998_n253;
  tri   P2_add_998_n252;
  tri   P2_add_998_n251;
  tri   P2_add_998_n249;
  tri   P2_add_998_n248;
  tri   P2_add_998_n247;
  tri   P2_add_998_n246;
  tri   P2_add_998_n245;
  tri   P2_add_998_n244;
  tri   P2_add_998_n243;
  tri   P2_add_998_n242;
  tri   P2_add_998_n241;
  tri   P2_add_998_n239;
  tri   P2_add_998_n238;
  tri   P2_add_998_n237;
  tri   P2_add_998_n236;
  tri   P2_add_998_n235;
  tri   P2_add_998_n234;
  tri   P2_add_998_n233;
  tri   P2_add_998_n232;
  tri   P2_add_998_n231;
  tri   P2_add_998_n229;
  tri   P2_add_998_n228;
  tri   P2_add_998_n227;
  tri   P2_add_998_n226;
  tri   P2_add_998_n225;
  tri   P2_add_998_n224;
  tri   P2_add_998_n223;
  tri   P2_add_998_n222;
  tri   P2_add_998_n221;
  tri   P2_add_998_n219;
  tri   P2_add_998_n218;
  tri   P2_add_998_n217;
  tri   P2_add_998_n216;
  tri   P2_add_998_n215;
  tri   P2_add_998_n214;
  tri   P2_add_998_n213;
  tri   P2_add_998_n212;
  tri   P2_add_998_n211;
  tri   P2_add_998_n209;
  tri   P2_add_998_n208;
  tri   P2_add_998_n207;
  tri   P2_add_998_n206;
  tri   P2_add_998_n205;
  tri   P2_add_998_n201;
  tri   P2_add_998_n204;
  tri   P2_add_998_n49;
  tri   P2_add_998_n296;
  tri   P2_sub_1030_n62;
  tri   P2_sub_1030_n61;
  tri   P2_sub_1030_n59;
  tri   P2_sub_1030_n58;
  tri   P2_sub_1030_n57;
  tri   P2_sub_1030_n55;
  tri   P2_sub_1030_n54;
  tri   P2_sub_1030_n52;
  tri   P2_sub_1030_n51;
  tri   P2_sub_1030_n50;
  tri   P2_sub_1030_n48;
  tri   P2_sub_1030_n47;
  tri   P2_sub_1030_n45;
  tri   P2_sub_1030_n44;
  tri   P2_sub_1030_n43;
  tri   P2_sub_1030_n41;
  tri   P2_sub_1030_n40;
  tri   P2_sub_1030_n38;
  tri   P2_sub_1030_n37;
  tri   P2_sub_1030_n36;
  tri   P2_sub_1030_n34;
  tri   P2_sub_1030_n33;
  tri   P2_sub_1030_n31;
  tri   P2_sub_1030_n30;
  tri   P2_sub_1030_n29;
  tri   P2_sub_1030_n27;
  tri   P2_sub_1030_n26;
  tri   P2_sub_1030_n24;
  tri   P2_sub_1030_n23;
  tri   P2_sub_1030_n22;
  tri   P2_sub_1030_n20;
  tri   P2_sub_1030_n19;
  tri   P2_sub_1030_n17;
  tri   P2_sub_1030_n16;
  tri   P2_sub_1030_n15;
  tri   P2_sub_1030_n13;
  tri   P2_sub_1030_n12;
  tri   P2_sub_1030_n10;
  tri   P2_sub_1030_n9;
  tri   P2_sub_1030_n8;
  tri   P2_sub_1030_n6;
  tri   P2_sub_1030_n5;
  tri   P2_sub_1030_n3;
  tri   P2_sub_1030_n2;
  tri   P2_sub_1030_n1;
  tri   P2_sub_1030_n151;
  tri   P2_sub_1030_n148;
  tri   P2_sub_1030_n147;
  tri   P2_sub_1030_n146;
  tri   P2_sub_1030_n145;
  tri   P2_sub_1030_n144;
  tri   P2_sub_1030_n142;
  tri   P2_sub_1030_n141;
  tri   P2_sub_1030_n140;
  tri   P2_sub_1030_n139;
  tri   P2_sub_1030_n138;
  tri   P2_sub_1030_n137;
  tri   P2_sub_1030_n136;
  tri   P2_sub_1030_n135;
  tri   P2_sub_1030_n134;
  tri   P2_sub_1030_n132;
  tri   P2_sub_1030_n131;
  tri   P2_sub_1030_n130;
  tri   P2_sub_1030_n129;
  tri   P2_sub_1030_n128;
  tri   P2_sub_1030_n127;
  tri   P2_sub_1030_n126;
  tri   P2_sub_1030_n125;
  tri   P2_sub_1030_n124;
  tri   P2_sub_1030_n122;
  tri   P2_sub_1030_n121;
  tri   P2_sub_1030_n120;
  tri   P2_sub_1030_n119;
  tri   P2_sub_1030_n118;
  tri   P2_sub_1030_n117;
  tri   P2_sub_1030_n116;
  tri   P2_sub_1030_n115;
  tri   P2_sub_1030_n114;
  tri   P2_sub_1030_n112;
  tri   P2_sub_1030_n111;
  tri   P2_sub_1030_n110;
  tri   P2_sub_1030_n109;
  tri   P2_sub_1030_n108;
  tri   P2_sub_1030_n107;
  tri   P2_sub_1030_n106;
  tri   P2_sub_1030_n105;
  tri   P2_sub_1030_n104;
  tri   P2_sub_1030_n102;
  tri   P2_sub_1030_n101;
  tri   P2_sub_1030_n100;
  tri   P2_sub_1030_n99;
  tri   P2_sub_1030_n98;
  tri   P2_sub_1030_n97;
  tri   P2_sub_1030_n96;
  tri   P2_sub_1030_n95;
  tri   P2_sub_1030_n94;
  tri   P2_sub_1030_n92;
  tri   P2_sub_1030_n91;
  tri   P2_sub_1030_n90;
  tri   P2_sub_1030_n89;
  tri   P2_sub_1030_n88;
  tri   P2_sub_1030_n87;
  tri   P2_sub_1030_n86;
  tri   P2_sub_1030_n85;
  tri   P2_sub_1030_n84;
  tri   P2_sub_1030_n82;
  tri   P2_sub_1030_n81;
  tri   P2_sub_1030_n80;
  tri   P2_sub_1030_n79;
  tri   P2_sub_1030_n78;
  tri   P2_sub_1030_n77;
  tri   P2_sub_1030_n76;
  tri   P2_sub_1030_n75;
  tri   P2_sub_1030_n74;
  tri   P2_sub_1030_n73;
  tri   P2_sub_1030_n71;
  tri   P2_sub_1030_n70;
  tri   P2_sub_1030_n69;
  tri   P2_sub_1030_n67;
  tri   P2_sub_1030_n68;
  tri   P2_sub_1030_n66;
  tri   P2_sub_1030_n65;
  tri   P2_sub_1030_n190;
  tri   P2_sub_1030_n189;
  tri   P2_sub_1030_n188;
  tri   P2_sub_1030_n60;
  tri   P2_sub_1030_n187;
  tri   P2_sub_1030_n186;
  tri   P2_sub_1030_n185;
  tri   P2_sub_1030_n184;
  tri   P2_sub_1030_n53;
  tri   P2_sub_1030_n183;
  tri   P2_sub_1030_n182;
  tri   P2_sub_1030_n181;
  tri   P2_sub_1030_n46;
  tri   P2_sub_1030_n180;
  tri   P2_sub_1030_n179;
  tri   P2_sub_1030_n178;
  tri   P2_sub_1030_n39;
  tri   P2_sub_1030_n177;
  tri   P2_sub_1030_n176;
  tri   P2_sub_1030_n175;
  tri   P2_sub_1030_n32;
  tri   P2_sub_1030_n174;
  tri   P2_sub_1030_n173;
  tri   P2_sub_1030_n172;
  tri   P2_sub_1030_n25;
  tri   P2_sub_1030_n171;
  tri   P2_sub_1030_n170;
  tri   P2_sub_1030_n169;
  tri   P2_sub_1030_n18;
  tri   P2_sub_1030_n168;
  tri   P2_sub_1030_n167;
  tri   P2_sub_1030_n166;
  tri   P2_sub_1030_n11;
  tri   P2_sub_1030_n165;
  tri   P2_sub_1030_n164;
  tri   P2_sub_1030_n163;
  tri   P2_sub_1030_n4;
  tri   P2_sub_1030_n162;
  tri   P2_sub_1030_n161;
  tri   P2_sub_1030_n160;
  tri   P2_sub_1030_n159;
  tri   P2_sub_1030_n158;
  tri   P2_sub_1030_n157;
  tri   P2_sub_1030_n149;
  tri   P2_sub_1030_n156;
  tri   P2_sub_1030_n155;
  tri   P2_sub_1030_n150;
  tri   P2_sub_1030_n152;
  tri   P2_sub_1030_n154;
  tri   P2_sub_1031_n88;
  tri   P2_sub_1031_n87;
  tri   P2_sub_1031_n86;
  tri   P2_sub_1031_n85;
  tri   P2_sub_1031_n82;
  tri   P2_sub_1031_n81;
  tri   P2_sub_1031_n80;
  tri   P2_sub_1031_n79;
  tri   P2_sub_1031_n78;
  tri   P2_sub_1031_n77;
  tri   P2_sub_1031_n76;
  tri   P2_sub_1031_n75;
  tri   P2_sub_1031_n74;
  tri   P2_sub_1031_n73;
  tri   P2_sub_1031_n71;
  tri   P2_sub_1031_n70;
  tri   P2_sub_1031_n69;
  tri   P2_sub_1031_n67;
  tri   P2_sub_1031_n68;
  tri   P2_sub_1031_n66;
  tri   P2_sub_1031_n65;
  tri   P2_sub_1031_n62;
  tri   P2_sub_1031_n61;
  tri   P2_sub_1031_n59;
  tri   P2_sub_1031_n58;
  tri   P2_sub_1031_n57;
  tri   P2_sub_1031_n55;
  tri   P2_sub_1031_n54;
  tri   P2_sub_1031_n52;
  tri   P2_sub_1031_n51;
  tri   P2_sub_1031_n50;
  tri   P2_sub_1031_n48;
  tri   P2_sub_1031_n47;
  tri   P2_sub_1031_n45;
  tri   P2_sub_1031_n44;
  tri   P2_sub_1031_n43;
  tri   P2_sub_1031_n41;
  tri   P2_sub_1031_n40;
  tri   P2_sub_1031_n38;
  tri   P2_sub_1031_n37;
  tri   P2_sub_1031_n36;
  tri   P2_sub_1031_n34;
  tri   P2_sub_1031_n33;
  tri   P2_sub_1031_n31;
  tri   P2_sub_1031_n30;
  tri   P2_sub_1031_n29;
  tri   P2_sub_1031_n27;
  tri   P2_sub_1031_n26;
  tri   P2_sub_1031_n24;
  tri   P2_sub_1031_n23;
  tri   P2_sub_1031_n22;
  tri   P2_sub_1031_n20;
  tri   P2_sub_1031_n19;
  tri   P2_sub_1031_n17;
  tri   P2_sub_1031_n16;
  tri   P2_sub_1031_n15;
  tri   P2_sub_1031_n13;
  tri   P2_sub_1031_n12;
  tri   P2_sub_1031_n10;
  tri   P2_sub_1031_n9;
  tri   P2_sub_1031_n8;
  tri   P2_sub_1031_n6;
  tri   P2_sub_1031_n5;
  tri   P2_sub_1031_n3;
  tri   P2_sub_1031_n2;
  tri   P2_sub_1031_n1;
  tri   P2_sub_1031_n18;
  tri   P2_sub_1031_n168;
  tri   P2_sub_1031_n167;
  tri   P2_sub_1031_n166;
  tri   P2_sub_1031_n11;
  tri   P2_sub_1031_n165;
  tri   P2_sub_1031_n164;
  tri   P2_sub_1031_n163;
  tri   P2_sub_1031_n4;
  tri   P2_sub_1031_n162;
  tri   P2_sub_1031_n161;
  tri   P2_sub_1031_n160;
  tri   P2_sub_1031_n158;
  tri   P2_sub_1031_n157;
  tri   P2_sub_1031_n156;
  tri   P2_sub_1031_n155;
  tri   P2_sub_1031_n154;
  tri   P2_sub_1031_n152;
  tri   P2_sub_1031_n151;
  tri   P2_sub_1031_n150;
  tri   P2_sub_1031_n149;
  tri   P2_sub_1031_n148;
  tri   P2_sub_1031_n147;
  tri   P2_sub_1031_n146;
  tri   P2_sub_1031_n145;
  tri   P2_sub_1031_n144;
  tri   P2_sub_1031_n142;
  tri   P2_sub_1031_n141;
  tri   P2_sub_1031_n140;
  tri   P2_sub_1031_n139;
  tri   P2_sub_1031_n138;
  tri   P2_sub_1031_n137;
  tri   P2_sub_1031_n136;
  tri   P2_sub_1031_n135;
  tri   P2_sub_1031_n134;
  tri   P2_sub_1031_n132;
  tri   P2_sub_1031_n131;
  tri   P2_sub_1031_n130;
  tri   P2_sub_1031_n129;
  tri   P2_sub_1031_n128;
  tri   P2_sub_1031_n127;
  tri   P2_sub_1031_n126;
  tri   P2_sub_1031_n125;
  tri   P2_sub_1031_n124;
  tri   P2_sub_1031_n122;
  tri   P2_sub_1031_n121;
  tri   P2_sub_1031_n120;
  tri   P2_sub_1031_n119;
  tri   P2_sub_1031_n118;
  tri   P2_sub_1031_n117;
  tri   P2_sub_1031_n116;
  tri   P2_sub_1031_n115;
  tri   P2_sub_1031_n114;
  tri   P2_sub_1031_n112;
  tri   P2_sub_1031_n111;
  tri   P2_sub_1031_n110;
  tri   P2_sub_1031_n109;
  tri   P2_sub_1031_n108;
  tri   P2_sub_1031_n107;
  tri   P2_sub_1031_n106;
  tri   P2_sub_1031_n105;
  tri   P2_sub_1031_n104;
  tri   P2_sub_1031_n102;
  tri   P2_sub_1031_n101;
  tri   P2_sub_1031_n100;
  tri   P2_sub_1031_n99;
  tri   P2_sub_1031_n98;
  tri   P2_sub_1031_n97;
  tri   P2_sub_1031_n89;
  tri   P2_sub_1031_n96;
  tri   P2_sub_1031_n95;
  tri   P2_sub_1031_n94;
  tri   P2_sub_1031_n92;
  tri   P2_sub_1031_n84;
  tri   P2_sub_1031_n91;
  tri   P2_sub_1031_n90;
  tri   P2_sub_1031_n190;
  tri   P2_sub_1031_n159;
  tri   P2_sub_1031_n189;
  tri   P2_sub_1031_n188;
  tri   P2_sub_1031_n60;
  tri   P2_sub_1031_n187;
  tri   P2_sub_1031_n186;
  tri   P2_sub_1031_n185;
  tri   P2_sub_1031_n184;
  tri   P2_sub_1031_n53;
  tri   P2_sub_1031_n183;
  tri   P2_sub_1031_n182;
  tri   P2_sub_1031_n181;
  tri   P2_sub_1031_n46;
  tri   P2_sub_1031_n180;
  tri   P2_sub_1031_n179;
  tri   P2_sub_1031_n178;
  tri   P2_sub_1031_n39;
  tri   P2_sub_1031_n177;
  tri   P2_sub_1031_n176;
  tri   P2_sub_1031_n175;
  tri   P2_sub_1031_n32;
  tri   P2_sub_1031_n174;
  tri   P2_sub_1031_n173;
  tri   P2_sub_1031_n172;
  tri   P2_sub_1031_n169;
  tri   P2_sub_1031_n25;
  tri   P2_sub_1031_n170;
  tri   P2_sub_1031_n171;
  tri   P2_lt_688_n62;
  tri   P2_lt_688_n60;
  tri   P2_lt_688_n59;
  tri   P2_lt_688_n58;
  tri   P2_lt_688_n57;
  tri   P2_lt_688_n56;
  tri   P2_lt_688_n55;
  tri   P2_lt_688_n52;
  tri   P2_lt_688_n51;
  tri   P2_lt_688_n50;
  tri   P2_lt_688_n49;
  tri   P2_lt_688_n48;
  tri   P2_lt_688_n47;
  tri   P2_lt_688_n46;
  tri   P2_lt_688_n45;
  tri   P2_lt_688_n42;
  tri   P2_lt_688_n41;
  tri   P2_lt_688_n40;
  tri   P2_lt_688_n39;
  tri   P2_lt_688_n38;
  tri   P2_lt_688_n37;
  tri   P2_lt_688_n36;
  tri   P2_lt_688_n35;
  tri   P2_lt_688_n32;
  tri   P2_lt_688_n31;
  tri   P2_lt_688_n30;
  tri   P2_lt_688_n29;
  tri   P2_lt_688_n28;
  tri   P2_lt_688_n27;
  tri   P2_lt_688_n26;
  tri   P2_lt_688_n25;
  tri   P2_lt_688_n22;
  tri   P2_lt_688_n21;
  tri   P2_lt_688_n20;
  tri   P2_lt_688_n19;
  tri   P2_lt_688_n18;
  tri   P2_lt_688_n17;
  tri   P2_lt_688_n16;
  tri   P2_lt_688_n15;
  tri   P2_lt_688_n12;
  tri   P2_lt_688_n11;
  tri   P2_lt_688_n10;
  tri   P2_lt_688_n9;
  tri   P2_lt_688_n8;
  tri   P2_lt_688_n7;
  tri   P2_lt_688_n6;
  tri   P2_lt_688_n4;
  tri   P2_lt_688_n3;
  tri   P2_lt_688_n2;
  tri   P2_lt_688_n156;
  tri   P2_lt_688_n155;
  tri   P2_lt_688_n154;
  tri   P2_lt_688_n153;
  tri   P2_lt_688_n152;
  tri   P2_lt_688_n151;
  tri   P2_lt_688_n150;
  tri   P2_lt_688_n149;
  tri   P2_lt_688_n148;
  tri   P2_lt_688_n147;
  tri   P2_lt_688_n146;
  tri   P2_lt_688_n145;
  tri   P2_lt_688_n144;
  tri   P2_lt_688_n143;
  tri   P2_lt_688_n142;
  tri   P2_lt_688_n141;
  tri   P2_lt_688_n140;
  tri   P2_lt_688_n139;
  tri   P2_lt_688_n138;
  tri   P2_lt_688_n137;
  tri   P2_lt_688_n136;
  tri   P2_lt_688_n135;
  tri   P2_lt_688_n134;
  tri   P2_lt_688_n133;
  tri   P2_lt_688_n132;
  tri   P2_lt_688_n131;
  tri   P2_lt_688_n130;
  tri   P2_lt_688_n129;
  tri   P2_lt_688_n128;
  tri   P2_lt_688_n127;
  tri   P2_lt_688_n126;
  tri   P2_lt_688_n125;
  tri   P2_lt_688_n124;
  tri   P2_lt_688_n123;
  tri   P2_lt_688_n122;
  tri   P2_lt_688_n121;
  tri   P2_lt_688_n120;
  tri   P2_lt_688_n119;
  tri   P2_lt_688_n118;
  tri   P2_lt_688_n117;
  tri   P2_lt_688_n116;
  tri   P2_lt_688_n115;
  tri   P2_lt_688_n114;
  tri   P2_lt_688_n113;
  tri   P2_lt_688_n112;
  tri   P2_lt_688_n110;
  tri   P2_lt_688_n109;
  tri   P2_lt_688_n108;
  tri   P2_lt_688_n107;
  tri   P2_lt_688_n106;
  tri   P2_lt_688_n105;
  tri   P2_lt_688_n104;
  tri   P2_lt_688_n103;
  tri   P2_lt_688_n102;
  tri   P2_lt_688_n101;
  tri   P2_lt_688_n100;
  tri   P2_lt_688_n99;
  tri   P2_lt_688_n98;
  tri   P2_lt_688_n97;
  tri   P2_lt_688_n96;
  tri   P2_lt_688_n95;
  tri   P2_lt_688_n94;
  tri   P2_lt_688_n93;
  tri   P2_lt_688_n92;
  tri   P2_lt_688_n91;
  tri   P2_lt_688_n90;
  tri   P2_lt_688_n89;
  tri   P2_lt_688_n88;
  tri   P2_lt_688_n87;
  tri   P2_lt_688_n86;
  tri   P2_lt_688_n85;
  tri   P2_lt_688_n84;
  tri   P2_lt_688_n83;
  tri   P2_lt_688_n82;
  tri   P2_lt_688_n81;
  tri   P2_lt_688_n80;
  tri   P2_lt_688_n79;
  tri   P2_lt_688_n78;
  tri   P2_lt_688_n77;
  tri   P2_lt_688_n76;
  tri   P2_lt_688_n75;
  tri   P2_lt_688_n74;
  tri   P2_lt_688_n73;
  tri   P2_lt_688_n72;
  tri   P2_lt_688_n71;
  tri   P2_lt_688_n70;
  tri   P2_lt_688_n69;
  tri   P2_lt_688_n68;
  tri   P2_lt_688_n67;
  tri   P2_lt_688_n66;
  tri   P2_lt_688_n65;
  tri   P2_lt_688_n61;
  tri   P2_lt_688_n1;
  tri   P2_lt_688_n5;
  tri   P2_lt_688_n14;
  tri   P2_lt_688_n13;
  tri   P2_lt_688_n24;
  tri   P2_lt_688_n23;
  tri   P2_lt_688_n34;
  tri   P2_lt_688_n33;
  tri   P2_lt_688_n44;
  tri   P2_lt_688_n43;
  tri   P2_lt_688_n54;
  tri   P2_lt_688_n53;
  tri   P2_lt_688_n64;
  tri   P2_lt_688_n63;
  tri   P1_sub_488_n94;
  tri   P1_sub_488_n93;
  tri   P1_sub_488_n90;
  tri   P1_sub_488_n89;
  tri   P1_sub_488_n88;
  tri   P1_sub_488_n87;
  tri   P1_sub_488_n86;
  tri   P1_sub_488_n84;
  tri   P1_sub_488_n83;
  tri   P1_sub_488_n82;
  tri   P1_sub_488_n81;
  tri   P1_sub_488_n80;
  tri   P1_sub_488_n79;
  tri   P1_sub_488_n78;
  tri   P1_sub_488_n77;
  tri   P1_sub_488_n76;
  tri   P1_sub_488_n75;
  tri   P1_sub_488_n74;
  tri   P1_sub_488_n73;
  tri   P1_sub_488_n72;
  tri   P1_sub_488_n71;
  tri   P1_sub_488_n70;
  tri   P1_sub_488_n69;
  tri   P1_sub_488_n67;
  tri   P1_sub_488_n66;
  tri   P1_sub_488_n65;
  tri   P1_sub_488_n64;
  tri   P1_sub_488_n63;
  tri   P1_sub_488_n62;
  tri   P1_sub_488_n61;
  tri   P1_sub_488_n59;
  tri   P1_sub_488_n60;
  tri   P1_sub_488_n58;
  tri   P1_sub_488_n57;
  tri   P1_sub_488_n55;
  tri   P1_sub_488_n54;
  tri   P1_sub_488_n52;
  tri   P1_sub_488_n51;
  tri   P1_sub_488_n50;
  tri   P1_sub_488_n48;
  tri   P1_sub_488_n47;
  tri   P1_sub_488_n45;
  tri   P1_sub_488_n44;
  tri   P1_sub_488_n43;
  tri   P1_sub_488_n41;
  tri   P1_sub_488_n40;
  tri   P1_sub_488_n38;
  tri   P1_sub_488_n37;
  tri   P1_sub_488_n36;
  tri   P1_sub_488_n34;
  tri   P1_sub_488_n33;
  tri   P1_sub_488_n31;
  tri   P1_sub_488_n30;
  tri   P1_sub_488_n29;
  tri   P1_sub_488_n27;
  tri   P1_sub_488_n26;
  tri   P1_sub_488_n24;
  tri   P1_sub_488_n23;
  tri   P1_sub_488_n22;
  tri   P1_sub_488_n20;
  tri   P1_sub_488_n19;
  tri   P1_sub_488_n17;
  tri   P1_sub_488_n16;
  tri   P1_sub_488_n15;
  tri   P1_sub_488_n13;
  tri   P1_sub_488_n12;
  tri   P1_sub_488_n10;
  tri   P1_sub_488_n9;
  tri   P1_sub_488_n8;
  tri   P1_sub_488_n6;
  tri   P1_sub_488_n5;
  tri   P1_sub_488_n3;
  tri   P1_sub_488_n2;
  tri   P1_sub_488_n1;
  tri   P1_sub_488_n181;
  tri   P1_sub_488_n178;
  tri   P1_sub_488_n177;
  tri   P1_sub_488_n176;
  tri   P1_sub_488_n175;
  tri   P1_sub_488_n174;
  tri   P1_sub_488_n172;
  tri   P1_sub_488_n171;
  tri   P1_sub_488_n170;
  tri   P1_sub_488_n169;
  tri   P1_sub_488_n168;
  tri   P1_sub_488_n167;
  tri   P1_sub_488_n166;
  tri   P1_sub_488_n165;
  tri   P1_sub_488_n164;
  tri   P1_sub_488_n163;
  tri   P1_sub_488_n162;
  tri   P1_sub_488_n161;
  tri   P1_sub_488_n160;
  tri   P1_sub_488_n159;
  tri   P1_sub_488_n158;
  tri   P1_sub_488_n157;
  tri   P1_sub_488_n154;
  tri   P1_sub_488_n153;
  tri   P1_sub_488_n151;
  tri   P1_sub_488_n150;
  tri   P1_sub_488_n149;
  tri   P1_sub_488_n148;
  tri   P1_sub_488_n147;
  tri   P1_sub_488_n146;
  tri   P1_sub_488_n145;
  tri   P1_sub_488_n144;
  tri   P1_sub_488_n143;
  tri   P1_sub_488_n142;
  tri   P1_sub_488_n141;
  tri   P1_sub_488_n140;
  tri   P1_sub_488_n139;
  tri   P1_sub_488_n138;
  tri   P1_sub_488_n137;
  tri   P1_sub_488_n136;
  tri   P1_sub_488_n135;
  tri   P1_sub_488_n134;
  tri   P1_sub_488_n133;
  tri   P1_sub_488_n132;
  tri   P1_sub_488_n131;
  tri   P1_sub_488_n130;
  tri   P1_sub_488_n129;
  tri   P1_sub_488_n128;
  tri   P1_sub_488_n127;
  tri   P1_sub_488_n126;
  tri   P1_sub_488_n125;
  tri   P1_sub_488_n124;
  tri   P1_sub_488_n123;
  tri   P1_sub_488_n122;
  tri   P1_sub_488_n121;
  tri   P1_sub_488_n120;
  tri   P1_sub_488_n119;
  tri   P1_sub_488_n118;
  tri   P1_sub_488_n117;
  tri   P1_sub_488_n116;
  tri   P1_sub_488_n115;
  tri   P1_sub_488_n114;
  tri   P1_sub_488_n113;
  tri   P1_sub_488_n112;
  tri   P1_sub_488_n111;
  tri   P1_sub_488_n110;
  tri   P1_sub_488_n109;
  tri   P1_sub_488_n95;
  tri   P1_sub_488_n108;
  tri   P1_sub_488_n107;
  tri   P1_sub_488_n106;
  tri   P1_sub_488_n105;
  tri   P1_sub_488_n104;
  tri   P1_sub_488_n103;
  tri   P1_sub_488_n102;
  tri   P1_sub_488_n101;
  tri   P1_sub_488_n100;
  tri   P1_sub_488_n99;
  tri   P1_sub_488_n85;
  tri   P1_sub_488_n91;
  tri   P1_sub_488_n98;
  tri   P1_sub_488_n97;
  tri   P1_sub_488_n92;
  tri   P1_sub_488_n96;
  tri   P1_sub_488_n28;
  tri   P1_sub_488_n260;
  tri   P1_sub_488_n18;
  tri   P1_sub_488_n21;
  tri   P1_sub_488_n258;
  tri   P1_sub_488_n257;
  tri   P1_sub_488_n256;
  tri   P1_sub_488_n11;
  tri   P1_sub_488_n14;
  tri   P1_sub_488_n255;
  tri   P1_sub_488_n254;
  tri   P1_sub_488_n253;
  tri   P1_sub_488_n4;
  tri   P1_sub_488_n7;
  tri   P1_sub_488_n252;
  tri   P1_sub_488_n251;
  tri   P1_sub_488_n250;
  tri   P1_sub_488_n248;
  tri   P1_sub_488_n247;
  tri   P1_sub_488_n246;
  tri   P1_sub_488_n245;
  tri   P1_sub_488_n244;
  tri   P1_sub_488_n242;
  tri   P1_sub_488_n241;
  tri   P1_sub_488_n240;
  tri   P1_sub_488_n239;
  tri   P1_sub_488_n238;
  tri   P1_sub_488_n237;
  tri   P1_sub_488_n236;
  tri   P1_sub_488_n235;
  tri   P1_sub_488_n234;
  tri   P1_sub_488_n233;
  tri   P1_sub_488_n232;
  tri   P1_sub_488_n231;
  tri   P1_sub_488_n230;
  tri   P1_sub_488_n229;
  tri   P1_sub_488_n228;
  tri   P1_sub_488_n227;
  tri   P1_sub_488_n226;
  tri   P1_sub_488_n225;
  tri   P1_sub_488_n224;
  tri   P1_sub_488_n223;
  tri   P1_sub_488_n222;
  tri   P1_sub_488_n221;
  tri   P1_sub_488_n220;
  tri   P1_sub_488_n219;
  tri   P1_sub_488_n218;
  tri   P1_sub_488_n217;
  tri   P1_sub_488_n216;
  tri   P1_sub_488_n215;
  tri   P1_sub_488_n214;
  tri   P1_sub_488_n213;
  tri   P1_sub_488_n212;
  tri   P1_sub_488_n211;
  tri   P1_sub_488_n210;
  tri   P1_sub_488_n209;
  tri   P1_sub_488_n208;
  tri   P1_sub_488_n207;
  tri   P1_sub_488_n206;
  tri   P1_sub_488_n205;
  tri   P1_sub_488_n204;
  tri   P1_sub_488_n203;
  tri   P1_sub_488_n202;
  tri   P1_sub_488_n201;
  tri   P1_sub_488_n200;
  tri   P1_sub_488_n199;
  tri   P1_sub_488_n198;
  tri   P1_sub_488_n197;
  tri   P1_sub_488_n183;
  tri   P1_sub_488_n196;
  tri   P1_sub_488_n195;
  tri   P1_sub_488_n194;
  tri   P1_sub_488_n193;
  tri   P1_sub_488_n192;
  tri   P1_sub_488_n191;
  tri   P1_sub_488_n190;
  tri   P1_sub_488_n189;
  tri   P1_sub_488_n188;
  tri   P1_sub_488_n187;
  tri   P1_sub_488_n173;
  tri   P1_sub_488_n179;
  tri   P1_sub_488_n186;
  tri   P1_sub_488_n185;
  tri   P1_sub_488_n180;
  tri   P1_sub_488_n182;
  tri   P1_sub_488_n184;
  tri   P1_sub_488_n281;
  tri   P1_sub_488_n280;
  tri   P1_sub_488_n243;
  tri   P1_sub_488_n249;
  tri   P1_sub_488_n279;
  tri   P1_sub_488_n278;
  tri   P1_sub_488_n152;
  tri   P1_sub_488_n277;
  tri   P1_sub_488_n156;
  tri   P1_sub_488_n276;
  tri   P1_sub_488_n275;
  tri   P1_sub_488_n274;
  tri   P1_sub_488_n53;
  tri   P1_sub_488_n56;
  tri   P1_sub_488_n273;
  tri   P1_sub_488_n272;
  tri   P1_sub_488_n271;
  tri   P1_sub_488_n46;
  tri   P1_sub_488_n49;
  tri   P1_sub_488_n270;
  tri   P1_sub_488_n269;
  tri   P1_sub_488_n268;
  tri   P1_sub_488_n39;
  tri   P1_sub_488_n42;
  tri   P1_sub_488_n267;
  tri   P1_sub_488_n266;
  tri   P1_sub_488_n265;
  tri   P1_sub_488_n32;
  tri   P1_sub_488_n35;
  tri   P1_sub_488_n264;
  tri   P1_sub_488_n263;
  tri   P1_sub_488_n262;
  tri   P1_sub_488_n259;
  tri   P1_sub_488_n261;
  tri   P1_sub_488_n25;
  tri   P1_lt_178_n72;
  tri   P1_lt_178_n70;
  tri   P1_lt_178_n69;
  tri   P1_lt_178_n68;
  tri   P1_lt_178_n67;
  tri   P1_lt_178_n66;
  tri   P1_lt_178_n65;
  tri   P1_lt_178_n62;
  tri   P1_lt_178_n61;
  tri   P1_lt_178_n60;
  tri   P1_lt_178_n59;
  tri   P1_lt_178_n58;
  tri   P1_lt_178_n57;
  tri   P1_lt_178_n56;
  tri   P1_lt_178_n55;
  tri   P1_lt_178_n52;
  tri   P1_lt_178_n51;
  tri   P1_lt_178_n50;
  tri   P1_lt_178_n49;
  tri   P1_lt_178_n48;
  tri   P1_lt_178_n47;
  tri   P1_lt_178_n46;
  tri   P1_lt_178_n45;
  tri   P1_lt_178_n42;
  tri   P1_lt_178_n41;
  tri   P1_lt_178_n40;
  tri   P1_lt_178_n39;
  tri   P1_lt_178_n38;
  tri   P1_lt_178_n37;
  tri   P1_lt_178_n36;
  tri   P1_lt_178_n35;
  tri   P1_lt_178_n32;
  tri   P1_lt_178_n31;
  tri   P1_lt_178_n30;
  tri   P1_lt_178_n29;
  tri   P1_lt_178_n28;
  tri   P1_lt_178_n27;
  tri   P1_lt_178_n26;
  tri   P1_lt_178_n25;
  tri   P1_lt_178_n22;
  tri   P1_lt_178_n21;
  tri   P1_lt_178_n20;
  tri   P1_lt_178_n19;
  tri   P1_lt_178_n18;
  tri   P1_lt_178_n17;
  tri   P1_lt_178_n16;
  tri   P1_lt_178_n15;
  tri   P1_lt_178_n12;
  tri   P1_lt_178_n11;
  tri   P1_lt_178_n10;
  tri   P1_lt_178_n9;
  tri   P1_lt_178_n8;
  tri   P1_lt_178_n7;
  tri   P1_lt_178_n6;
  tri   P1_lt_178_n4;
  tri   P1_lt_178_n3;
  tri   P1_lt_178_n2;
  tri   P1_lt_178_n34;
  tri   P1_lt_178_n33;
  tri   P1_lt_178_n44;
  tri   P1_lt_178_n43;
  tri   P1_lt_178_n54;
  tri   P1_lt_178_n53;
  tri   P1_lt_178_n64;
  tri   P1_lt_178_n63;
  tri   P1_lt_178_n73;
  tri   P1_lt_178_n156;
  tri   P1_lt_178_n155;
  tri   P1_lt_178_n154;
  tri   P1_lt_178_n153;
  tri   P1_lt_178_n152;
  tri   P1_lt_178_n151;
  tri   P1_lt_178_n150;
  tri   P1_lt_178_n149;
  tri   P1_lt_178_n148;
  tri   P1_lt_178_n147;
  tri   P1_lt_178_n146;
  tri   P1_lt_178_n145;
  tri   P1_lt_178_n144;
  tri   P1_lt_178_n143;
  tri   P1_lt_178_n142;
  tri   P1_lt_178_n141;
  tri   P1_lt_178_n140;
  tri   P1_lt_178_n139;
  tri   P1_lt_178_n138;
  tri   P1_lt_178_n137;
  tri   P1_lt_178_n136;
  tri   P1_lt_178_n135;
  tri   P1_lt_178_n134;
  tri   P1_lt_178_n133;
  tri   P1_lt_178_n132;
  tri   P1_lt_178_n131;
  tri   P1_lt_178_n130;
  tri   P1_lt_178_n129;
  tri   P1_lt_178_n128;
  tri   P1_lt_178_n127;
  tri   P1_lt_178_n126;
  tri   P1_lt_178_n125;
  tri   P1_lt_178_n124;
  tri   P1_lt_178_n123;
  tri   P1_lt_178_n122;
  tri   P1_lt_178_n121;
  tri   P1_lt_178_n120;
  tri   P1_lt_178_n119;
  tri   P1_lt_178_n118;
  tri   P1_lt_178_n117;
  tri   P1_lt_178_n116;
  tri   P1_lt_178_n115;
  tri   P1_lt_178_n114;
  tri   P1_lt_178_n113;
  tri   P1_lt_178_n112;
  tri   P1_lt_178_n110;
  tri   P1_lt_178_n109;
  tri   P1_lt_178_n108;
  tri   P1_lt_178_n107;
  tri   P1_lt_178_n106;
  tri   P1_lt_178_n105;
  tri   P1_lt_178_n104;
  tri   P1_lt_178_n103;
  tri   P1_lt_178_n102;
  tri   P1_lt_178_n101;
  tri   P1_lt_178_n100;
  tri   P1_lt_178_n99;
  tri   P1_lt_178_n98;
  tri   P1_lt_178_n97;
  tri   P1_lt_178_n96;
  tri   P1_lt_178_n95;
  tri   P1_lt_178_n94;
  tri   P1_lt_178_n93;
  tri   P1_lt_178_n92;
  tri   P1_lt_178_n91;
  tri   P1_lt_178_n90;
  tri   P1_lt_178_n89;
  tri   P1_lt_178_n88;
  tri   P1_lt_178_n87;
  tri   P1_lt_178_n86;
  tri   P1_lt_178_n85;
  tri   P1_lt_178_n84;
  tri   P1_lt_178_n83;
  tri   P1_lt_178_n82;
  tri   P1_lt_178_n81;
  tri   P1_lt_178_n80;
  tri   P1_lt_178_n79;
  tri   P1_lt_178_n78;
  tri   P1_lt_178_n77;
  tri   P1_lt_178_n76;
  tri   P1_lt_178_n75;
  tri   P1_lt_178_n74;
  tri   P1_lt_178_n71;
  tri   P1_lt_178_n1;
  tri   P1_lt_178_n5;
  tri   P1_lt_178_n14;
  tri   P1_lt_178_n13;
  tri   P1_lt_178_n24;
  tri   P1_lt_178_n23;
  tri   P1_lt_186_n37;
  tri   P1_lt_186_n35;
  tri   P1_lt_186_n32;
  tri   P1_lt_186_n31;
  tri   P1_lt_186_n30;
  tri   P1_lt_186_n29;
  tri   P1_lt_186_n28;
  tri   P1_lt_186_n27;
  tri   P1_lt_186_n26;
  tri   P1_lt_186_n25;
  tri   P1_lt_186_n22;
  tri   P1_lt_186_n21;
  tri   P1_lt_186_n20;
  tri   P1_lt_186_n19;
  tri   P1_lt_186_n18;
  tri   P1_lt_186_n17;
  tri   P1_lt_186_n16;
  tri   P1_lt_186_n15;
  tri   P1_lt_186_n12;
  tri   P1_lt_186_n11;
  tri   P1_lt_186_n10;
  tri   P1_lt_186_n9;
  tri   P1_lt_186_n8;
  tri   P1_lt_186_n7;
  tri   P1_lt_186_n6;
  tri   P1_lt_186_n4;
  tri   P1_lt_186_n3;
  tri   P1_lt_186_n2;
  tri   P1_lt_186_n152;
  tri   P1_lt_186_n150;
  tri   P1_lt_186_n149;
  tri   P1_lt_186_n148;
  tri   P1_lt_186_n147;
  tri   P1_lt_186_n146;
  tri   P1_lt_186_n145;
  tri   P1_lt_186_n142;
  tri   P1_lt_186_n141;
  tri   P1_lt_186_n140;
  tri   P1_lt_186_n139;
  tri   P1_lt_186_n138;
  tri   P1_lt_186_n137;
  tri   P1_lt_186_n136;
  tri   P1_lt_186_n135;
  tri   P1_lt_186_n132;
  tri   P1_lt_186_n131;
  tri   P1_lt_186_n130;
  tri   P1_lt_186_n129;
  tri   P1_lt_186_n128;
  tri   P1_lt_186_n127;
  tri   P1_lt_186_n126;
  tri   P1_lt_186_n125;
  tri   P1_lt_186_n122;
  tri   P1_lt_186_n121;
  tri   P1_lt_186_n120;
  tri   P1_lt_186_n119;
  tri   P1_lt_186_n118;
  tri   P1_lt_186_n117;
  tri   P1_lt_186_n116;
  tri   P1_lt_186_n115;
  tri   P1_lt_186_n113;
  tri   P1_lt_186_n112;
  tri   P1_lt_186_n110;
  tri   P1_lt_186_n109;
  tri   P1_lt_186_n108;
  tri   P1_lt_186_n107;
  tri   P1_lt_186_n106;
  tri   P1_lt_186_n105;
  tri   P1_lt_186_n102;
  tri   P1_lt_186_n101;
  tri   P1_lt_186_n100;
  tri   P1_lt_186_n99;
  tri   P1_lt_186_n98;
  tri   P1_lt_186_n97;
  tri   P1_lt_186_n96;
  tri   P1_lt_186_n95;
  tri   P1_lt_186_n92;
  tri   P1_lt_186_n91;
  tri   P1_lt_186_n90;
  tri   P1_lt_186_n89;
  tri   P1_lt_186_n88;
  tri   P1_lt_186_n87;
  tri   P1_lt_186_n86;
  tri   P1_lt_186_n85;
  tri   P1_lt_186_n82;
  tri   P1_lt_186_n81;
  tri   P1_lt_186_n80;
  tri   P1_lt_186_n79;
  tri   P1_lt_186_n78;
  tri   P1_lt_186_n77;
  tri   P1_lt_186_n76;
  tri   P1_lt_186_n75;
  tri   P1_lt_186_n72;
  tri   P1_lt_186_n71;
  tri   P1_lt_186_n70;
  tri   P1_lt_186_n69;
  tri   P1_lt_186_n68;
  tri   P1_lt_186_n67;
  tri   P1_lt_186_n66;
  tri   P1_lt_186_n65;
  tri   P1_lt_186_n62;
  tri   P1_lt_186_n61;
  tri   P1_lt_186_n60;
  tri   P1_lt_186_n59;
  tri   P1_lt_186_n58;
  tri   P1_lt_186_n57;
  tri   P1_lt_186_n56;
  tri   P1_lt_186_n55;
  tri   P1_lt_186_n52;
  tri   P1_lt_186_n51;
  tri   P1_lt_186_n50;
  tri   P1_lt_186_n49;
  tri   P1_lt_186_n48;
  tri   P1_lt_186_n47;
  tri   P1_lt_186_n46;
  tri   P1_lt_186_n45;
  tri   P1_lt_186_n42;
  tri   P1_lt_186_n41;
  tri   P1_lt_186_n38;
  tri   P1_lt_186_n36;
  tri   P1_lt_186_n40;
  tri   P1_lt_186_n39;
  tri   P1_lt_186_n1;
  tri   P1_lt_186_n5;
  tri   P1_lt_186_n14;
  tri   P1_lt_186_n13;
  tri   P1_lt_186_n24;
  tri   P1_lt_186_n23;
  tri   P1_lt_186_n34;
  tri   P1_lt_186_n33;
  tri   P1_lt_186_n44;
  tri   P1_lt_186_n43;
  tri   P1_lt_186_n54;
  tri   P1_lt_186_n53;
  tri   P1_lt_186_n64;
  tri   P1_lt_186_n63;
  tri   P1_lt_186_n74;
  tri   P1_lt_186_n73;
  tri   P1_lt_186_n84;
  tri   P1_lt_186_n83;
  tri   P1_lt_186_n94;
  tri   P1_lt_186_n93;
  tri   P1_lt_186_n104;
  tri   P1_lt_186_n103;
  tri   P1_lt_186_n114;
  tri   P1_lt_186_n124;
  tri   P1_lt_186_n123;
  tri   P1_lt_186_n134;
  tri   P1_lt_186_n133;
  tri   P1_lt_186_n144;
  tri   P1_lt_186_n143;
  tri   P1_lt_186_n156;
  tri   P1_lt_186_n153;
  tri   P1_lt_186_n154;
  tri   P1_lt_186_n155;
  tri   P1_lt_186_n151;
  tri   P1_lt_224_n117;
  tri   P1_lt_224_n115;
  tri   P1_lt_224_n113;
  tri   P1_lt_224_n112;
  tri   P1_lt_224_n110;
  tri   P1_lt_224_n109;
  tri   P1_lt_224_n108;
  tri   P1_lt_224_n107;
  tri   P1_lt_224_n106;
  tri   P1_lt_224_n105;
  tri   P1_lt_224_n102;
  tri   P1_lt_224_n101;
  tri   P1_lt_224_n100;
  tri   P1_lt_224_n99;
  tri   P1_lt_224_n98;
  tri   P1_lt_224_n97;
  tri   P1_lt_224_n96;
  tri   P1_lt_224_n95;
  tri   P1_lt_224_n92;
  tri   P1_lt_224_n91;
  tri   P1_lt_224_n90;
  tri   P1_lt_224_n89;
  tri   P1_lt_224_n88;
  tri   P1_lt_224_n87;
  tri   P1_lt_224_n86;
  tri   P1_lt_224_n85;
  tri   P1_lt_224_n82;
  tri   P1_lt_224_n81;
  tri   P1_lt_224_n80;
  tri   P1_lt_224_n79;
  tri   P1_lt_224_n78;
  tri   P1_lt_224_n77;
  tri   P1_lt_224_n76;
  tri   P1_lt_224_n75;
  tri   P1_lt_224_n72;
  tri   P1_lt_224_n71;
  tri   P1_lt_224_n70;
  tri   P1_lt_224_n69;
  tri   P1_lt_224_n68;
  tri   P1_lt_224_n67;
  tri   P1_lt_224_n66;
  tri   P1_lt_224_n65;
  tri   P1_lt_224_n62;
  tri   P1_lt_224_n61;
  tri   P1_lt_224_n60;
  tri   P1_lt_224_n59;
  tri   P1_lt_224_n58;
  tri   P1_lt_224_n57;
  tri   P1_lt_224_n56;
  tri   P1_lt_224_n55;
  tri   P1_lt_224_n52;
  tri   P1_lt_224_n51;
  tri   P1_lt_224_n50;
  tri   P1_lt_224_n49;
  tri   P1_lt_224_n48;
  tri   P1_lt_224_n47;
  tri   P1_lt_224_n46;
  tri   P1_lt_224_n45;
  tri   P1_lt_224_n42;
  tri   P1_lt_224_n41;
  tri   P1_lt_224_n40;
  tri   P1_lt_224_n39;
  tri   P1_lt_224_n38;
  tri   P1_lt_224_n37;
  tri   P1_lt_224_n36;
  tri   P1_lt_224_n35;
  tri   P1_lt_224_n32;
  tri   P1_lt_224_n31;
  tri   P1_lt_224_n30;
  tri   P1_lt_224_n29;
  tri   P1_lt_224_n28;
  tri   P1_lt_224_n27;
  tri   P1_lt_224_n26;
  tri   P1_lt_224_n25;
  tri   P1_lt_224_n22;
  tri   P1_lt_224_n21;
  tri   P1_lt_224_n20;
  tri   P1_lt_224_n19;
  tri   P1_lt_224_n18;
  tri   P1_lt_224_n17;
  tri   P1_lt_224_n16;
  tri   P1_lt_224_n15;
  tri   P1_lt_224_n12;
  tri   P1_lt_224_n11;
  tri   P1_lt_224_n10;
  tri   P1_lt_224_n9;
  tri   P1_lt_224_n8;
  tri   P1_lt_224_n7;
  tri   P1_lt_224_n6;
  tri   P1_lt_224_n4;
  tri   P1_lt_224_n3;
  tri   P1_lt_224_n2;
  tri   P1_lt_224_n1;
  tri   P1_lt_224_n5;
  tri   P1_lt_224_n14;
  tri   P1_lt_224_n13;
  tri   P1_lt_224_n24;
  tri   P1_lt_224_n23;
  tri   P1_lt_224_n34;
  tri   P1_lt_224_n33;
  tri   P1_lt_224_n44;
  tri   P1_lt_224_n43;
  tri   P1_lt_224_n54;
  tri   P1_lt_224_n53;
  tri   P1_lt_224_n64;
  tri   P1_lt_224_n63;
  tri   P1_lt_224_n74;
  tri   P1_lt_224_n73;
  tri   P1_lt_224_n84;
  tri   P1_lt_224_n83;
  tri   P1_lt_224_n94;
  tri   P1_lt_224_n93;
  tri   P1_lt_224_n104;
  tri   P1_lt_224_n103;
  tri   P1_lt_224_n114;
  tri   P1_lt_224_n156;
  tri   P1_lt_224_n155;
  tri   P1_lt_224_n154;
  tri   P1_lt_224_n153;
  tri   P1_lt_224_n152;
  tri   P1_lt_224_n151;
  tri   P1_lt_224_n150;
  tri   P1_lt_224_n149;
  tri   P1_lt_224_n148;
  tri   P1_lt_224_n147;
  tri   P1_lt_224_n146;
  tri   P1_lt_224_n145;
  tri   P1_lt_224_n144;
  tri   P1_lt_224_n143;
  tri   P1_lt_224_n142;
  tri   P1_lt_224_n141;
  tri   P1_lt_224_n140;
  tri   P1_lt_224_n139;
  tri   P1_lt_224_n138;
  tri   P1_lt_224_n137;
  tri   P1_lt_224_n136;
  tri   P1_lt_224_n135;
  tri   P1_lt_224_n134;
  tri   P1_lt_224_n133;
  tri   P1_lt_224_n132;
  tri   P1_lt_224_n131;
  tri   P1_lt_224_n130;
  tri   P1_lt_224_n129;
  tri   P1_lt_224_n128;
  tri   P1_lt_224_n127;
  tri   P1_lt_224_n126;
  tri   P1_lt_224_n125;
  tri   P1_lt_224_n124;
  tri   P1_lt_224_n123;
  tri   P1_lt_224_n122;
  tri   P1_lt_224_n121;
  tri   P1_lt_224_n118;
  tri   P1_lt_224_n116;
  tri   P1_lt_224_n120;
  tri   P1_lt_224_n119;
  tri   P1_lt_232_n80;
  tri   P1_lt_232_n78;
  tri   P1_lt_232_n77;
  tri   P1_lt_232_n76;
  tri   P1_lt_232_n75;
  tri   P1_lt_232_n72;
  tri   P1_lt_232_n71;
  tri   P1_lt_232_n70;
  tri   P1_lt_232_n69;
  tri   P1_lt_232_n68;
  tri   P1_lt_232_n67;
  tri   P1_lt_232_n66;
  tri   P1_lt_232_n65;
  tri   P1_lt_232_n62;
  tri   P1_lt_232_n61;
  tri   P1_lt_232_n60;
  tri   P1_lt_232_n59;
  tri   P1_lt_232_n58;
  tri   P1_lt_232_n57;
  tri   P1_lt_232_n56;
  tri   P1_lt_232_n55;
  tri   P1_lt_232_n52;
  tri   P1_lt_232_n51;
  tri   P1_lt_232_n50;
  tri   P1_lt_232_n49;
  tri   P1_lt_232_n48;
  tri   P1_lt_232_n47;
  tri   P1_lt_232_n46;
  tri   P1_lt_232_n45;
  tri   P1_lt_232_n42;
  tri   P1_lt_232_n41;
  tri   P1_lt_232_n40;
  tri   P1_lt_232_n39;
  tri   P1_lt_232_n38;
  tri   P1_lt_232_n37;
  tri   P1_lt_232_n36;
  tri   P1_lt_232_n35;
  tri   P1_lt_232_n32;
  tri   P1_lt_232_n31;
  tri   P1_lt_232_n30;
  tri   P1_lt_232_n29;
  tri   P1_lt_232_n28;
  tri   P1_lt_232_n27;
  tri   P1_lt_232_n26;
  tri   P1_lt_232_n25;
  tri   P1_lt_232_n22;
  tri   P1_lt_232_n21;
  tri   P1_lt_232_n20;
  tri   P1_lt_232_n19;
  tri   P1_lt_232_n18;
  tri   P1_lt_232_n17;
  tri   P1_lt_232_n16;
  tri   P1_lt_232_n15;
  tri   P1_lt_232_n12;
  tri   P1_lt_232_n11;
  tri   P1_lt_232_n10;
  tri   P1_lt_232_n9;
  tri   P1_lt_232_n8;
  tri   P1_lt_232_n7;
  tri   P1_lt_232_n6;
  tri   P1_lt_232_n4;
  tri   P1_lt_232_n3;
  tri   P1_lt_232_n2;
  tri   P1_lt_232_n1;
  tri   P1_lt_232_n5;
  tri   P1_lt_232_n14;
  tri   P1_lt_232_n13;
  tri   P1_lt_232_n24;
  tri   P1_lt_232_n23;
  tri   P1_lt_232_n34;
  tri   P1_lt_232_n33;
  tri   P1_lt_232_n44;
  tri   P1_lt_232_n43;
  tri   P1_lt_232_n54;
  tri   P1_lt_232_n53;
  tri   P1_lt_232_n64;
  tri   P1_lt_232_n63;
  tri   P1_lt_232_n74;
  tri   P1_lt_232_n73;
  tri   P1_lt_232_n156;
  tri   P1_lt_232_n155;
  tri   P1_lt_232_n154;
  tri   P1_lt_232_n153;
  tri   P1_lt_232_n152;
  tri   P1_lt_232_n151;
  tri   P1_lt_232_n150;
  tri   P1_lt_232_n149;
  tri   P1_lt_232_n148;
  tri   P1_lt_232_n147;
  tri   P1_lt_232_n146;
  tri   P1_lt_232_n145;
  tri   P1_lt_232_n144;
  tri   P1_lt_232_n143;
  tri   P1_lt_232_n142;
  tri   P1_lt_232_n141;
  tri   P1_lt_232_n140;
  tri   P1_lt_232_n139;
  tri   P1_lt_232_n138;
  tri   P1_lt_232_n137;
  tri   P1_lt_232_n136;
  tri   P1_lt_232_n135;
  tri   P1_lt_232_n134;
  tri   P1_lt_232_n133;
  tri   P1_lt_232_n132;
  tri   P1_lt_232_n131;
  tri   P1_lt_232_n130;
  tri   P1_lt_232_n129;
  tri   P1_lt_232_n128;
  tri   P1_lt_232_n127;
  tri   P1_lt_232_n126;
  tri   P1_lt_232_n125;
  tri   P1_lt_232_n124;
  tri   P1_lt_232_n123;
  tri   P1_lt_232_n122;
  tri   P1_lt_232_n121;
  tri   P1_lt_232_n120;
  tri   P1_lt_232_n119;
  tri   P1_lt_232_n118;
  tri   P1_lt_232_n117;
  tri   P1_lt_232_n116;
  tri   P1_lt_232_n115;
  tri   P1_lt_232_n114;
  tri   P1_lt_232_n113;
  tri   P1_lt_232_n112;
  tri   P1_lt_232_n110;
  tri   P1_lt_232_n109;
  tri   P1_lt_232_n108;
  tri   P1_lt_232_n107;
  tri   P1_lt_232_n106;
  tri   P1_lt_232_n105;
  tri   P1_lt_232_n104;
  tri   P1_lt_232_n103;
  tri   P1_lt_232_n102;
  tri   P1_lt_232_n101;
  tri   P1_lt_232_n100;
  tri   P1_lt_232_n99;
  tri   P1_lt_232_n98;
  tri   P1_lt_232_n97;
  tri   P1_lt_232_n96;
  tri   P1_lt_232_n95;
  tri   P1_lt_232_n94;
  tri   P1_lt_232_n93;
  tri   P1_lt_232_n92;
  tri   P1_lt_232_n91;
  tri   P1_lt_232_n90;
  tri   P1_lt_232_n89;
  tri   P1_lt_232_n88;
  tri   P1_lt_232_n87;
  tri   P1_lt_232_n86;
  tri   P1_lt_232_n85;
  tri   P1_lt_232_n84;
  tri   P1_lt_232_n83;
  tri   P1_lt_232_n82;
  tri   P1_lt_232_n81;
  tri   P1_lt_232_n79;
  tri   P2_sub_858_n2;
  tri   P2_sub_858_n100;
  tri   P2_sub_858_n99;
  tri   P2_sub_858_n98;
  tri   P2_sub_858_n97;
  tri   P2_sub_858_n94;
  tri   P2_sub_858_n93;
  tri   P2_sub_858_n92;
  tri   P2_sub_858_n91;
  tri   P2_sub_858_n90;
  tri   P2_sub_858_n89;
  tri   P2_sub_858_n88;
  tri   P2_sub_858_n87;
  tri   P2_sub_858_n86;
  tri   P2_sub_858_n85;
  tri   P2_sub_858_n84;
  tri   P2_sub_858_n83;
  tri   P2_sub_858_n82;
  tri   P2_sub_858_n81;
  tri   P2_sub_858_n80;
  tri   P2_sub_858_n79;
  tri   P2_sub_858_n78;
  tri   P2_sub_858_n77;
  tri   P2_sub_858_n76;
  tri   P2_sub_858_n75;
  tri   P2_sub_858_n74;
  tri   P2_sub_858_n73;
  tri   P2_sub_858_n72;
  tri   P2_sub_858_n71;
  tri   P2_sub_858_n70;
  tri   P2_sub_858_n69;
  tri   P2_sub_858_n67;
  tri   P2_sub_858_n66;
  tri   P2_sub_858_n65;
  tri   P2_sub_858_n64;
  tri   P2_sub_858_n63;
  tri   P2_sub_858_n62;
  tri   P2_sub_858_n61;
  tri   P2_sub_858_n59;
  tri   P2_sub_858_n60;
  tri   P2_sub_858_n58;
  tri   P2_sub_858_n57;
  tri   P2_sub_858_n55;
  tri   P2_sub_858_n54;
  tri   P2_sub_858_n52;
  tri   P2_sub_858_n51;
  tri   P2_sub_858_n50;
  tri   P2_sub_858_n48;
  tri   P2_sub_858_n47;
  tri   P2_sub_858_n45;
  tri   P2_sub_858_n44;
  tri   P2_sub_858_n43;
  tri   P2_sub_858_n41;
  tri   P2_sub_858_n40;
  tri   P2_sub_858_n38;
  tri   P2_sub_858_n37;
  tri   P2_sub_858_n36;
  tri   P2_sub_858_n34;
  tri   P2_sub_858_n33;
  tri   P2_sub_858_n31;
  tri   P2_sub_858_n30;
  tri   P2_sub_858_n29;
  tri   P2_sub_858_n27;
  tri   P2_sub_858_n26;
  tri   P2_sub_858_n24;
  tri   P2_sub_858_n23;
  tri   P2_sub_858_n22;
  tri   P2_sub_858_n20;
  tri   P2_sub_858_n19;
  tri   P2_sub_858_n17;
  tri   P2_sub_858_n16;
  tri   P2_sub_858_n15;
  tri   P2_sub_858_n13;
  tri   P2_sub_858_n12;
  tri   P2_sub_858_n10;
  tri   P2_sub_858_n9;
  tri   P2_sub_858_n8;
  tri   P2_sub_858_n6;
  tri   P2_sub_858_n5;
  tri   P2_sub_858_n1;
  tri   P2_sub_858_n3;
  tri   P2_sub_858_n188;
  tri   P2_sub_858_n186;
  tri   P2_sub_858_n185;
  tri   P2_sub_858_n182;
  tri   P2_sub_858_n181;
  tri   P2_sub_858_n180;
  tri   P2_sub_858_n179;
  tri   P2_sub_858_n178;
  tri   P2_sub_858_n177;
  tri   P2_sub_858_n176;
  tri   P2_sub_858_n175;
  tri   P2_sub_858_n174;
  tri   P2_sub_858_n173;
  tri   P2_sub_858_n172;
  tri   P2_sub_858_n171;
  tri   P2_sub_858_n170;
  tri   P2_sub_858_n169;
  tri   P2_sub_858_n168;
  tri   P2_sub_858_n167;
  tri   P2_sub_858_n166;
  tri   P2_sub_858_n165;
  tri   P2_sub_858_n164;
  tri   P2_sub_858_n163;
  tri   P2_sub_858_n162;
  tri   P2_sub_858_n161;
  tri   P2_sub_858_n160;
  tri   P2_sub_858_n159;
  tri   P2_sub_858_n158;
  tri   P2_sub_858_n157;
  tri   P2_sub_858_n154;
  tri   P2_sub_858_n153;
  tri   P2_sub_858_n151;
  tri   P2_sub_858_n150;
  tri   P2_sub_858_n149;
  tri   P2_sub_858_n148;
  tri   P2_sub_858_n147;
  tri   P2_sub_858_n146;
  tri   P2_sub_858_n145;
  tri   P2_sub_858_n144;
  tri   P2_sub_858_n143;
  tri   P2_sub_858_n142;
  tri   P2_sub_858_n141;
  tri   P2_sub_858_n140;
  tri   P2_sub_858_n139;
  tri   P2_sub_858_n138;
  tri   P2_sub_858_n137;
  tri   P2_sub_858_n136;
  tri   P2_sub_858_n135;
  tri   P2_sub_858_n134;
  tri   P2_sub_858_n133;
  tri   P2_sub_858_n132;
  tri   P2_sub_858_n131;
  tri   P2_sub_858_n130;
  tri   P2_sub_858_n129;
  tri   P2_sub_858_n128;
  tri   P2_sub_858_n127;
  tri   P2_sub_858_n126;
  tri   P2_sub_858_n125;
  tri   P2_sub_858_n124;
  tri   P2_sub_858_n123;
  tri   P2_sub_858_n122;
  tri   P2_sub_858_n121;
  tri   P2_sub_858_n120;
  tri   P2_sub_858_n119;
  tri   P2_sub_858_n118;
  tri   P2_sub_858_n117;
  tri   P2_sub_858_n116;
  tri   P2_sub_858_n115;
  tri   P2_sub_858_n114;
  tri   P2_sub_858_n113;
  tri   P2_sub_858_n112;
  tri   P2_sub_858_n111;
  tri   P2_sub_858_n110;
  tri   P2_sub_858_n109;
  tri   P2_sub_858_n95;
  tri   P2_sub_858_n101;
  tri   P2_sub_858_n108;
  tri   P2_sub_858_n107;
  tri   P2_sub_858_n106;
  tri   P2_sub_858_n105;
  tri   P2_sub_858_n104;
  tri   P2_sub_858_n96;
  tri   P2_sub_858_n103;
  tri   P2_sub_858_n102;
  tri   P2_sub_858_n32;
  tri   P2_sub_858_n35;
  tri   P2_sub_858_n264;
  tri   P2_sub_858_n263;
  tri   P2_sub_858_n262;
  tri   P2_sub_858_n25;
  tri   P2_sub_858_n28;
  tri   P2_sub_858_n261;
  tri   P2_sub_858_n260;
  tri   P2_sub_858_n259;
  tri   P2_sub_858_n18;
  tri   P2_sub_858_n21;
  tri   P2_sub_858_n258;
  tri   P2_sub_858_n257;
  tri   P2_sub_858_n256;
  tri   P2_sub_858_n11;
  tri   P2_sub_858_n14;
  tri   P2_sub_858_n255;
  tri   P2_sub_858_n254;
  tri   P2_sub_858_n253;
  tri   P2_sub_858_n4;
  tri   P2_sub_858_n7;
  tri   P2_sub_858_n252;
  tri   P2_sub_858_n251;
  tri   P2_sub_858_n250;
  tri   P2_sub_858_n248;
  tri   P2_sub_858_n247;
  tri   P2_sub_858_n246;
  tri   P2_sub_858_n245;
  tri   P2_sub_858_n244;
  tri   P2_sub_858_n242;
  tri   P2_sub_858_n241;
  tri   P2_sub_858_n240;
  tri   P2_sub_858_n239;
  tri   P2_sub_858_n238;
  tri   P2_sub_858_n237;
  tri   P2_sub_858_n236;
  tri   P2_sub_858_n235;
  tri   P2_sub_858_n234;
  tri   P2_sub_858_n233;
  tri   P2_sub_858_n232;
  tri   P2_sub_858_n231;
  tri   P2_sub_858_n230;
  tri   P2_sub_858_n229;
  tri   P2_sub_858_n228;
  tri   P2_sub_858_n227;
  tri   P2_sub_858_n226;
  tri   P2_sub_858_n225;
  tri   P2_sub_858_n224;
  tri   P2_sub_858_n223;
  tri   P2_sub_858_n222;
  tri   P2_sub_858_n221;
  tri   P2_sub_858_n220;
  tri   P2_sub_858_n219;
  tri   P2_sub_858_n218;
  tri   P2_sub_858_n217;
  tri   P2_sub_858_n216;
  tri   P2_sub_858_n215;
  tri   P2_sub_858_n214;
  tri   P2_sub_858_n213;
  tri   P2_sub_858_n212;
  tri   P2_sub_858_n211;
  tri   P2_sub_858_n210;
  tri   P2_sub_858_n209;
  tri   P2_sub_858_n208;
  tri   P2_sub_858_n207;
  tri   P2_sub_858_n206;
  tri   P2_sub_858_n205;
  tri   P2_sub_858_n204;
  tri   P2_sub_858_n203;
  tri   P2_sub_858_n202;
  tri   P2_sub_858_n201;
  tri   P2_sub_858_n200;
  tri   P2_sub_858_n199;
  tri   P2_sub_858_n198;
  tri   P2_sub_858_n197;
  tri   P2_sub_858_n183;
  tri   P2_sub_858_n196;
  tri   P2_sub_858_n195;
  tri   P2_sub_858_n194;
  tri   P2_sub_858_n193;
  tri   P2_sub_858_n192;
  tri   P2_sub_858_n191;
  tri   P2_sub_858_n190;
  tri   P2_sub_858_n187;
  tri   P2_sub_858_n184;
  tri   P2_sub_858_n189;
  tri   P2_sub_858_n281;
  tri   P2_sub_858_n280;
  tri   P2_sub_858_n243;
  tri   P2_sub_858_n249;
  tri   P2_sub_858_n279;
  tri   P2_sub_858_n278;
  tri   P2_sub_858_n152;
  tri   P2_sub_858_n277;
  tri   P2_sub_858_n156;
  tri   P2_sub_858_n276;
  tri   P2_sub_858_n275;
  tri   P2_sub_858_n274;
  tri   P2_sub_858_n53;
  tri   P2_sub_858_n56;
  tri   P2_sub_858_n273;
  tri   P2_sub_858_n272;
  tri   P2_sub_858_n271;
  tri   P2_sub_858_n46;
  tri   P2_sub_858_n49;
  tri   P2_sub_858_n270;
  tri   P2_sub_858_n269;
  tri   P2_sub_858_n268;
  tri   P2_sub_858_n265;
  tri   P2_sub_858_n39;
  tri   P2_sub_858_n266;
  tri   P2_sub_858_n42;
  tri   P2_sub_858_n267;
  tri   P2_sub_878_n37;
  tri   P2_sub_878_n36;
  tri   P2_sub_878_n34;
  tri   P2_sub_878_n33;
  tri   P2_sub_878_n31;
  tri   P2_sub_878_n30;
  tri   P2_sub_878_n29;
  tri   P2_sub_878_n27;
  tri   P2_sub_878_n26;
  tri   P2_sub_878_n24;
  tri   P2_sub_878_n23;
  tri   P2_sub_878_n22;
  tri   P2_sub_878_n20;
  tri   P2_sub_878_n19;
  tri   P2_sub_878_n17;
  tri   P2_sub_878_n16;
  tri   P2_sub_878_n15;
  tri   P2_sub_878_n13;
  tri   P2_sub_878_n12;
  tri   P2_sub_878_n10;
  tri   P2_sub_878_n9;
  tri   P2_sub_878_n8;
  tri   P2_sub_878_n6;
  tri   P2_sub_878_n5;
  tri   P2_sub_878_n3;
  tri   P2_sub_878_n2;
  tri   P2_sub_878_n1;
  tri   P2_sub_878_n128;
  tri   P2_sub_878_n127;
  tri   P2_sub_878_n124;
  tri   P2_sub_878_n123;
  tri   P2_sub_878_n122;
  tri   P2_sub_878_n121;
  tri   P2_sub_878_n120;
  tri   P2_sub_878_n119;
  tri   P2_sub_878_n118;
  tri   P2_sub_878_n117;
  tri   P2_sub_878_n116;
  tri   P2_sub_878_n115;
  tri   P2_sub_878_n114;
  tri   P2_sub_878_n113;
  tri   P2_sub_878_n112;
  tri   P2_sub_878_n111;
  tri   P2_sub_878_n110;
  tri   P2_sub_878_n109;
  tri   P2_sub_878_n108;
  tri   P2_sub_878_n107;
  tri   P2_sub_878_n106;
  tri   P2_sub_878_n105;
  tri   P2_sub_878_n104;
  tri   P2_sub_878_n103;
  tri   P2_sub_878_n102;
  tri   P2_sub_878_n101;
  tri   P2_sub_878_n100;
  tri   P2_sub_878_n99;
  tri   P2_sub_878_n98;
  tri   P2_sub_878_n97;
  tri   P2_sub_878_n96;
  tri   P2_sub_878_n95;
  tri   P2_sub_878_n94;
  tri   P2_sub_878_n93;
  tri   P2_sub_878_n92;
  tri   P2_sub_878_n91;
  tri   P2_sub_878_n90;
  tri   P2_sub_878_n89;
  tri   P2_sub_878_n88;
  tri   P2_sub_878_n87;
  tri   P2_sub_878_n86;
  tri   P2_sub_878_n85;
  tri   P2_sub_878_n84;
  tri   P2_sub_878_n83;
  tri   P2_sub_878_n82;
  tri   P2_sub_878_n81;
  tri   P2_sub_878_n80;
  tri   P2_sub_878_n79;
  tri   P2_sub_878_n78;
  tri   P2_sub_878_n77;
  tri   P2_sub_878_n76;
  tri   P2_sub_878_n75;
  tri   P2_sub_878_n74;
  tri   P2_sub_878_n73;
  tri   P2_sub_878_n72;
  tri   P2_sub_878_n71;
  tri   P2_sub_878_n70;
  tri   P2_sub_878_n69;
  tri   P2_sub_878_n67;
  tri   P2_sub_878_n66;
  tri   P2_sub_878_n65;
  tri   P2_sub_878_n64;
  tri   P2_sub_878_n63;
  tri   P2_sub_878_n62;
  tri   P2_sub_878_n61;
  tri   P2_sub_878_n59;
  tri   P2_sub_878_n60;
  tri   P2_sub_878_n58;
  tri   P2_sub_878_n57;
  tri   P2_sub_878_n55;
  tri   P2_sub_878_n54;
  tri   P2_sub_878_n52;
  tri   P2_sub_878_n51;
  tri   P2_sub_878_n50;
  tri   P2_sub_878_n48;
  tri   P2_sub_878_n47;
  tri   P2_sub_878_n45;
  tri   P2_sub_878_n44;
  tri   P2_sub_878_n43;
  tri   P2_sub_878_n38;
  tri   P2_sub_878_n41;
  tri   P2_sub_878_n40;
  tri   P2_sub_878_n216;
  tri   P2_sub_878_n215;
  tri   P2_sub_878_n212;
  tri   P2_sub_878_n211;
  tri   P2_sub_878_n210;
  tri   P2_sub_878_n209;
  tri   P2_sub_878_n208;
  tri   P2_sub_878_n207;
  tri   P2_sub_878_n206;
  tri   P2_sub_878_n205;
  tri   P2_sub_878_n204;
  tri   P2_sub_878_n203;
  tri   P2_sub_878_n202;
  tri   P2_sub_878_n201;
  tri   P2_sub_878_n200;
  tri   P2_sub_878_n199;
  tri   P2_sub_878_n198;
  tri   P2_sub_878_n197;
  tri   P2_sub_878_n196;
  tri   P2_sub_878_n195;
  tri   P2_sub_878_n194;
  tri   P2_sub_878_n193;
  tri   P2_sub_878_n192;
  tri   P2_sub_878_n191;
  tri   P2_sub_878_n190;
  tri   P2_sub_878_n189;
  tri   P2_sub_878_n188;
  tri   P2_sub_878_n187;
  tri   P2_sub_878_n186;
  tri   P2_sub_878_n185;
  tri   P2_sub_878_n184;
  tri   P2_sub_878_n183;
  tri   P2_sub_878_n182;
  tri   P2_sub_878_n181;
  tri   P2_sub_878_n180;
  tri   P2_sub_878_n179;
  tri   P2_sub_878_n178;
  tri   P2_sub_878_n177;
  tri   P2_sub_878_n176;
  tri   P2_sub_878_n175;
  tri   P2_sub_878_n174;
  tri   P2_sub_878_n173;
  tri   P2_sub_878_n172;
  tri   P2_sub_878_n171;
  tri   P2_sub_878_n170;
  tri   P2_sub_878_n169;
  tri   P2_sub_878_n168;
  tri   P2_sub_878_n167;
  tri   P2_sub_878_n166;
  tri   P2_sub_878_n165;
  tri   P2_sub_878_n164;
  tri   P2_sub_878_n163;
  tri   P2_sub_878_n162;
  tri   P2_sub_878_n161;
  tri   P2_sub_878_n160;
  tri   P2_sub_878_n159;
  tri   P2_sub_878_n158;
  tri   P2_sub_878_n157;
  tri   P2_sub_878_n154;
  tri   P2_sub_878_n153;
  tri   P2_sub_878_n151;
  tri   P2_sub_878_n150;
  tri   P2_sub_878_n149;
  tri   P2_sub_878_n148;
  tri   P2_sub_878_n147;
  tri   P2_sub_878_n146;
  tri   P2_sub_878_n145;
  tri   P2_sub_878_n144;
  tri   P2_sub_878_n143;
  tri   P2_sub_878_n142;
  tri   P2_sub_878_n141;
  tri   P2_sub_878_n140;
  tri   P2_sub_878_n139;
  tri   P2_sub_878_n125;
  tri   P2_sub_878_n138;
  tri   P2_sub_878_n137;
  tri   P2_sub_878_n136;
  tri   P2_sub_878_n135;
  tri   P2_sub_878_n134;
  tri   P2_sub_878_n133;
  tri   P2_sub_878_n132;
  tri   P2_sub_878_n129;
  tri   P2_sub_878_n130;
  tri   P2_sub_878_n131;
  tri   P2_sub_878_n126;
  tri   P2_sub_878_n281;
  tri   P2_sub_878_n280;
  tri   P2_sub_878_n279;
  tri   P2_sub_878_n278;
  tri   P2_sub_878_n152;
  tri   P2_sub_878_n277;
  tri   P2_sub_878_n156;
  tri   P2_sub_878_n276;
  tri   P2_sub_878_n275;
  tri   P2_sub_878_n274;
  tri   P2_sub_878_n53;
  tri   P2_sub_878_n56;
  tri   P2_sub_878_n273;
  tri   P2_sub_878_n272;
  tri   P2_sub_878_n271;
  tri   P2_sub_878_n46;
  tri   P2_sub_878_n49;
  tri   P2_sub_878_n270;
  tri   P2_sub_878_n269;
  tri   P2_sub_878_n268;
  tri   P2_sub_878_n39;
  tri   P2_sub_878_n42;
  tri   P2_sub_878_n267;
  tri   P2_sub_878_n266;
  tri   P2_sub_878_n265;
  tri   P2_sub_878_n32;
  tri   P2_sub_878_n35;
  tri   P2_sub_878_n264;
  tri   P2_sub_878_n263;
  tri   P2_sub_878_n262;
  tri   P2_sub_878_n25;
  tri   P2_sub_878_n28;
  tri   P2_sub_878_n261;
  tri   P2_sub_878_n260;
  tri   P2_sub_878_n259;
  tri   P2_sub_878_n18;
  tri   P2_sub_878_n21;
  tri   P2_sub_878_n258;
  tri   P2_sub_878_n257;
  tri   P2_sub_878_n256;
  tri   P2_sub_878_n11;
  tri   P2_sub_878_n14;
  tri   P2_sub_878_n255;
  tri   P2_sub_878_n254;
  tri   P2_sub_878_n253;
  tri   P2_sub_878_n4;
  tri   P2_sub_878_n7;
  tri   P2_sub_878_n252;
  tri   P2_sub_878_n251;
  tri   P2_sub_878_n250;
  tri   P2_sub_878_n249;
  tri   P2_sub_878_n248;
  tri   P2_sub_878_n247;
  tri   P2_sub_878_n246;
  tri   P2_sub_878_n245;
  tri   P2_sub_878_n244;
  tri   P2_sub_878_n243;
  tri   P2_sub_878_n242;
  tri   P2_sub_878_n241;
  tri   P2_sub_878_n240;
  tri   P2_sub_878_n239;
  tri   P2_sub_878_n238;
  tri   P2_sub_878_n237;
  tri   P2_sub_878_n236;
  tri   P2_sub_878_n235;
  tri   P2_sub_878_n234;
  tri   P2_sub_878_n233;
  tri   P2_sub_878_n232;
  tri   P2_sub_878_n231;
  tri   P2_sub_878_n230;
  tri   P2_sub_878_n229;
  tri   P2_sub_878_n228;
  tri   P2_sub_878_n227;
  tri   P2_sub_878_n213;
  tri   P2_sub_878_n226;
  tri   P2_sub_878_n225;
  tri   P2_sub_878_n224;
  tri   P2_sub_878_n223;
  tri   P2_sub_878_n222;
  tri   P2_sub_878_n221;
  tri   P2_sub_878_n220;
  tri   P2_sub_878_n219;
  tri   P2_sub_878_n214;
  tri   P2_sub_878_n218;
  tri   P2_sub_878_n217;
  tri   P2_add_898_n63;
  tri   P2_add_898_n62;
  tri   P2_add_898_n61;
  tri   P2_add_898_n59;
  tri   P2_add_898_n58;
  tri   P2_add_898_n57;
  tri   P2_add_898_n55;
  tri   P2_add_898_n54;
  tri   P2_add_898_n53;
  tri   P2_add_898_n51;
  tri   P2_add_898_n50;
  tri   P2_add_898_n48;
  tri   P2_add_898_n47;
  tri   P2_add_898_n46;
  tri   P2_add_898_n44;
  tri   P2_add_898_n43;
  tri   P2_add_898_n41;
  tri   P2_add_898_n40;
  tri   P2_add_898_n39;
  tri   P2_add_898_n37;
  tri   P2_add_898_n36;
  tri   P2_add_898_n34;
  tri   P2_add_898_n33;
  tri   P2_add_898_n32;
  tri   P2_add_898_n30;
  tri   P2_add_898_n29;
  tri   P2_add_898_n27;
  tri   P2_add_898_n26;
  tri   P2_add_898_n25;
  tri   P2_add_898_n23;
  tri   P2_add_898_n22;
  tri   P2_add_898_n20;
  tri   P2_add_898_n19;
  tri   P2_add_898_n18;
  tri   P2_add_898_n16;
  tri   P2_add_898_n15;
  tri   P2_add_898_n13;
  tri   P2_add_898_n12;
  tri   P2_add_898_n11;
  tri   P2_add_898_n9;
  tri   P2_add_898_n8;
  tri   P2_add_898_n6;
  tri   P2_add_898_n5;
  tri   P2_add_898_n4;
  tri   P2_add_898_n2;
  tri   P2_add_898_n1;
  tri   P2_add_898_n146;
  tri   P2_add_898_n145;
  tri   P2_add_898_n144;
  tri   P2_add_898_n142;
  tri   P2_add_898_n141;
  tri   P2_add_898_n140;
  tri   P2_add_898_n139;
  tri   P2_add_898_n138;
  tri   P2_add_898_n137;
  tri   P2_add_898_n136;
  tri   P2_add_898_n135;
  tri   P2_add_898_n134;
  tri   P2_add_898_n132;
  tri   P2_add_898_n131;
  tri   P2_add_898_n130;
  tri   P2_add_898_n129;
  tri   P2_add_898_n128;
  tri   P2_add_898_n127;
  tri   P2_add_898_n126;
  tri   P2_add_898_n125;
  tri   P2_add_898_n124;
  tri   P2_add_898_n122;
  tri   P2_add_898_n121;
  tri   P2_add_898_n120;
  tri   P2_add_898_n119;
  tri   P2_add_898_n118;
  tri   P2_add_898_n117;
  tri   P2_add_898_n116;
  tri   P2_add_898_n115;
  tri   P2_add_898_n114;
  tri   P2_add_898_n112;
  tri   P2_add_898_n111;
  tri   P2_add_898_n110;
  tri   P2_add_898_n109;
  tri   P2_add_898_n108;
  tri   P2_add_898_n107;
  tri   P2_add_898_n106;
  tri   P2_add_898_n105;
  tri   P2_add_898_n104;
  tri   P2_add_898_n102;
  tri   P2_add_898_n101;
  tri   P2_add_898_n100;
  tri   P2_add_898_n99;
  tri   P2_add_898_n98;
  tri   P2_add_898_n97;
  tri   P2_add_898_n96;
  tri   P2_add_898_n95;
  tri   P2_add_898_n94;
  tri   P2_add_898_n92;
  tri   P2_add_898_n91;
  tri   P2_add_898_n90;
  tri   P2_add_898_n89;
  tri   P2_add_898_n88;
  tri   P2_add_898_n87;
  tri   P2_add_898_n86;
  tri   P2_add_898_n85;
  tri   P2_add_898_n84;
  tri   P2_add_898_n82;
  tri   P2_add_898_n81;
  tri   P2_add_898_n80;
  tri   P2_add_898_n79;
  tri   P2_add_898_n78;
  tri   P2_add_898_n77;
  tri   P2_add_898_n76;
  tri   P2_add_898_n75;
  tri   P2_add_898_n74;
  tri   P2_add_898_n72;
  tri   P2_add_898_n71;
  tri   P2_add_898_n70;
  tri   P2_add_898_n64;
  tri   P2_add_898_n69;
  tri   P2_add_898_n68;
  tri   P2_add_898_n60;
  tri   P2_add_898_n66;
  tri   P2_add_898_n65;
  tri   P2_add_898_n233;
  tri   P2_add_898_n232;
  tri   P2_add_898_n231;
  tri   P2_add_898_n229;
  tri   P2_add_898_n228;
  tri   P2_add_898_n227;
  tri   P2_add_898_n226;
  tri   P2_add_898_n225;
  tri   P2_add_898_n224;
  tri   P2_add_898_n223;
  tri   P2_add_898_n222;
  tri   P2_add_898_n221;
  tri   P2_add_898_n219;
  tri   P2_add_898_n218;
  tri   P2_add_898_n217;
  tri   P2_add_898_n216;
  tri   P2_add_898_n215;
  tri   P2_add_898_n214;
  tri   P2_add_898_n213;
  tri   P2_add_898_n212;
  tri   P2_add_898_n211;
  tri   P2_add_898_n209;
  tri   P2_add_898_n208;
  tri   P2_add_898_n207;
  tri   P2_add_898_n206;
  tri   P2_add_898_n205;
  tri   P2_add_898_n204;
  tri   P2_add_898_n203;
  tri   P2_add_898_n202;
  tri   P2_add_898_n201;
  tri   P2_add_898_n199;
  tri   P2_add_898_n198;
  tri   P2_add_898_n197;
  tri   P2_add_898_n196;
  tri   P2_add_898_n195;
  tri   P2_add_898_n194;
  tri   P2_add_898_n193;
  tri   P2_add_898_n192;
  tri   P2_add_898_n191;
  tri   P2_add_898_n189;
  tri   P2_add_898_n188;
  tri   P2_add_898_n187;
  tri   P2_add_898_n186;
  tri   P2_add_898_n185;
  tri   P2_add_898_n184;
  tri   P2_add_898_n183;
  tri   P2_add_898_n182;
  tri   P2_add_898_n181;
  tri   P2_add_898_n179;
  tri   P2_add_898_n178;
  tri   P2_add_898_n177;
  tri   P2_add_898_n176;
  tri   P2_add_898_n175;
  tri   P2_add_898_n174;
  tri   P2_add_898_n173;
  tri   P2_add_898_n172;
  tri   P2_add_898_n171;
  tri   P2_add_898_n169;
  tri   P2_add_898_n168;
  tri   P2_add_898_n167;
  tri   P2_add_898_n166;
  tri   P2_add_898_n165;
  tri   P2_add_898_n164;
  tri   P2_add_898_n163;
  tri   P2_add_898_n162;
  tri   P2_add_898_n161;
  tri   P2_add_898_n159;
  tri   P2_add_898_n158;
  tri   P2_add_898_n157;
  tri   P2_add_898_n147;
  tri   P2_add_898_n156;
  tri   P2_add_898_n155;
  tri   P2_add_898_n153;
  tri   P2_add_898_n152;
  tri   P2_add_898_n148;
  tri   P2_add_898_n149;
  tri   P2_add_898_n150;
  tri   P2_add_898_n279;
  tri   P2_add_898_n278;
  tri   P2_add_898_n151;
  tri   P2_add_898_n277;
  tri   P2_add_898_n276;
  tri   P2_add_898_n275;
  tri   P2_add_898_n52;
  tri   P2_add_898_n274;
  tri   P2_add_898_n273;
  tri   P2_add_898_n272;
  tri   P2_add_898_n45;
  tri   P2_add_898_n271;
  tri   P2_add_898_n270;
  tri   P2_add_898_n269;
  tri   P2_add_898_n38;
  tri   P2_add_898_n268;
  tri   P2_add_898_n267;
  tri   P2_add_898_n266;
  tri   P2_add_898_n31;
  tri   P2_add_898_n265;
  tri   P2_add_898_n264;
  tri   P2_add_898_n263;
  tri   P2_add_898_n24;
  tri   P2_add_898_n262;
  tri   P2_add_898_n261;
  tri   P2_add_898_n260;
  tri   P2_add_898_n17;
  tri   P2_add_898_n259;
  tri   P2_add_898_n258;
  tri   P2_add_898_n257;
  tri   P2_add_898_n10;
  tri   P2_add_898_n256;
  tri   P2_add_898_n255;
  tri   P2_add_898_n254;
  tri   P2_add_898_n3;
  tri   P2_add_898_n253;
  tri   P2_add_898_n252;
  tri   P2_add_898_n251;
  tri   P2_add_898_n249;
  tri   P2_add_898_n248;
  tri   P2_add_898_n247;
  tri   P2_add_898_n246;
  tri   P2_add_898_n245;
  tri   P2_add_898_n244;
  tri   P2_add_898_n243;
  tri   P2_add_898_n242;
  tri   P2_add_898_n241;
  tri   P2_add_898_n239;
  tri   P2_add_898_n238;
  tri   P2_add_898_n237;
  tri   P2_add_898_n234;
  tri   P2_add_898_n236;
  tri   P2_add_898_n235;
  tri   P2_add_898_n299;
  tri   P1_sub_273_n25;
  tri   P1_sub_273_n24;
  tri   P1_sub_273_n23;
  tri   P1_sub_273_n22;
  tri   P1_sub_273_n20;
  tri   P1_sub_273_n19;
  tri   P1_sub_273_n18;
  tri   P1_sub_273_n16;
  tri   P1_sub_273_n15;
  tri   P1_sub_273_n14;
  tri   P1_sub_273_n13;
  tri   P1_sub_273_n12;
  tri   P1_sub_273_n11;
  tri   P1_sub_273_n10;
  tri   P1_sub_273_n9;
  tri   P1_sub_273_n7;
  tri   P1_sub_273_n6;
  tri   P1_sub_273_n5;
  tri   P1_sub_273_n3;
  tri   P1_sub_273_n2;
  tri   P1_sub_273_n100;
  tri   P1_sub_273_n99;
  tri   P1_sub_273_n98;
  tri   P1_sub_273_n96;
  tri   P1_sub_273_n95;
  tri   P1_sub_273_n94;
  tri   P1_sub_273_n93;
  tri   P1_sub_273_n92;
  tri   P1_sub_273_n91;
  tri   P1_sub_273_n90;
  tri   P1_sub_273_n89;
  tri   P1_sub_273_n88;
  tri   P1_sub_273_n87;
  tri   P1_sub_273_n86;
  tri   P1_sub_273_n85;
  tri   P1_sub_273_n84;
  tri   P1_sub_273_n83;
  tri   P1_sub_273_n82;
  tri   P1_sub_273_n81;
  tri   P1_sub_273_n80;
  tri   P1_sub_273_n79;
  tri   P1_sub_273_n78;
  tri   P1_sub_273_n77;
  tri   P1_sub_273_n76;
  tri   P1_sub_273_n75;
  tri   P1_sub_273_n74;
  tri   P1_sub_273_n73;
  tri   P1_sub_273_n72;
  tri   P1_sub_273_n71;
  tri   P1_sub_273_n70;
  tri   P1_sub_273_n69;
  tri   P1_sub_273_n68;
  tri   P1_sub_273_n67;
  tri   P1_sub_273_n66;
  tri   P1_sub_273_n65;
  tri   P1_sub_273_n64;
  tri   P1_sub_273_n62;
  tri   P1_sub_273_n61;
  tri   P1_sub_273_n60;
  tri   P1_sub_273_n59;
  tri   P1_sub_273_n58;
  tri   P1_sub_273_n57;
  tri   P1_sub_273_n56;
  tri   P1_sub_273_n55;
  tri   P1_sub_273_n54;
  tri   P1_sub_273_n53;
  tri   P1_sub_273_n52;
  tri   P1_sub_273_n51;
  tri   P1_sub_273_n50;
  tri   P1_sub_273_n49;
  tri   P1_sub_273_n48;
  tri   P1_sub_273_n47;
  tri   P1_sub_273_n46;
  tri   P1_sub_273_n45;
  tri   P1_sub_273_n44;
  tri   P1_sub_273_n43;
  tri   P1_sub_273_n42;
  tri   P1_sub_273_n41;
  tri   P1_sub_273_n40;
  tri   P1_sub_273_n39;
  tri   P1_sub_273_n38;
  tri   P1_sub_273_n37;
  tri   P1_sub_273_n36;
  tri   P1_sub_273_n35;
  tri   P1_sub_273_n34;
  tri   P1_sub_273_n33;
  tri   P1_sub_273_n32;
  tri   P1_sub_273_n31;
  tri   P1_sub_273_n30;
  tri   P1_sub_273_n29;
  tri   P1_sub_273_n28;
  tri   P1_sub_273_n27;
  tri   P1_sub_273_n26;
  tri   P1_sub_273_n104;
  tri   P1_sub_273_n21;
  tri   P1_sub_273_n103;
  tri   P1_sub_273_n17;
  tri   P1_sub_273_n102;
  tri   P1_sub_273_n8;
  tri   P1_sub_273_n101;
  tri   P1_sub_273_n97;
  tri   P1_sub_273_n4;
  tri   P1_add_348_n58;
  tri   P1_add_348_n57;
  tri   P1_add_348_n55;
  tri   P1_add_348_n54;
  tri   P1_add_348_n53;
  tri   P1_add_348_n51;
  tri   P1_add_348_n50;
  tri   P1_add_348_n48;
  tri   P1_add_348_n47;
  tri   P1_add_348_n46;
  tri   P1_add_348_n44;
  tri   P1_add_348_n43;
  tri   P1_add_348_n41;
  tri   P1_add_348_n40;
  tri   P1_add_348_n39;
  tri   P1_add_348_n37;
  tri   P1_add_348_n36;
  tri   P1_add_348_n34;
  tri   P1_add_348_n33;
  tri   P1_add_348_n32;
  tri   P1_add_348_n30;
  tri   P1_add_348_n29;
  tri   P1_add_348_n27;
  tri   P1_add_348_n26;
  tri   P1_add_348_n25;
  tri   P1_add_348_n23;
  tri   P1_add_348_n22;
  tri   P1_add_348_n20;
  tri   P1_add_348_n19;
  tri   P1_add_348_n18;
  tri   P1_add_348_n16;
  tri   P1_add_348_n15;
  tri   P1_add_348_n13;
  tri   P1_add_348_n12;
  tri   P1_add_348_n11;
  tri   P1_add_348_n9;
  tri   P1_add_348_n8;
  tri   P1_add_348_n6;
  tri   P1_add_348_n5;
  tri   P1_add_348_n4;
  tri   P1_add_348_n2;
  tri   P1_add_348_n1;
  tri   P1_add_348_n142;
  tri   P1_add_348_n141;
  tri   P1_add_348_n140;
  tri   P1_add_348_n139;
  tri   P1_add_348_n138;
  tri   P1_add_348_n137;
  tri   P1_add_348_n136;
  tri   P1_add_348_n135;
  tri   P1_add_348_n134;
  tri   P1_add_348_n132;
  tri   P1_add_348_n131;
  tri   P1_add_348_n130;
  tri   P1_add_348_n129;
  tri   P1_add_348_n128;
  tri   P1_add_348_n127;
  tri   P1_add_348_n126;
  tri   P1_add_348_n125;
  tri   P1_add_348_n124;
  tri   P1_add_348_n122;
  tri   P1_add_348_n121;
  tri   P1_add_348_n120;
  tri   P1_add_348_n119;
  tri   P1_add_348_n118;
  tri   P1_add_348_n117;
  tri   P1_add_348_n116;
  tri   P1_add_348_n115;
  tri   P1_add_348_n114;
  tri   P1_add_348_n112;
  tri   P1_add_348_n111;
  tri   P1_add_348_n110;
  tri   P1_add_348_n109;
  tri   P1_add_348_n108;
  tri   P1_add_348_n107;
  tri   P1_add_348_n106;
  tri   P1_add_348_n105;
  tri   P1_add_348_n104;
  tri   P1_add_348_n102;
  tri   P1_add_348_n101;
  tri   P1_add_348_n100;
  tri   P1_add_348_n99;
  tri   P1_add_348_n98;
  tri   P1_add_348_n97;
  tri   P1_add_348_n96;
  tri   P1_add_348_n95;
  tri   P1_add_348_n94;
  tri   P1_add_348_n92;
  tri   P1_add_348_n91;
  tri   P1_add_348_n90;
  tri   P1_add_348_n89;
  tri   P1_add_348_n88;
  tri   P1_add_348_n87;
  tri   P1_add_348_n86;
  tri   P1_add_348_n85;
  tri   P1_add_348_n84;
  tri   P1_add_348_n82;
  tri   P1_add_348_n81;
  tri   P1_add_348_n80;
  tri   P1_add_348_n79;
  tri   P1_add_348_n78;
  tri   P1_add_348_n77;
  tri   P1_add_348_n76;
  tri   P1_add_348_n75;
  tri   P1_add_348_n74;
  tri   P1_add_348_n72;
  tri   P1_add_348_n71;
  tri   P1_add_348_n70;
  tri   P1_add_348_n69;
  tri   P1_add_348_n68;
  tri   P1_add_348_n60;
  tri   P1_add_348_n66;
  tri   P1_add_348_n65;
  tri   P1_add_348_n64;
  tri   P1_add_348_n63;
  tri   P1_add_348_n59;
  tri   P1_add_348_n62;
  tri   P1_add_348_n61;
  tri   P1_add_348_n229;
  tri   P1_add_348_n228;
  tri   P1_add_348_n227;
  tri   P1_add_348_n226;
  tri   P1_add_348_n225;
  tri   P1_add_348_n223;
  tri   P1_add_348_n222;
  tri   P1_add_348_n221;
  tri   P1_add_348_n219;
  tri   P1_add_348_n218;
  tri   P1_add_348_n217;
  tri   P1_add_348_n216;
  tri   P1_add_348_n215;
  tri   P1_add_348_n214;
  tri   P1_add_348_n213;
  tri   P1_add_348_n212;
  tri   P1_add_348_n211;
  tri   P1_add_348_n209;
  tri   P1_add_348_n208;
  tri   P1_add_348_n207;
  tri   P1_add_348_n206;
  tri   P1_add_348_n205;
  tri   P1_add_348_n204;
  tri   P1_add_348_n203;
  tri   P1_add_348_n202;
  tri   P1_add_348_n201;
  tri   P1_add_348_n199;
  tri   P1_add_348_n198;
  tri   P1_add_348_n197;
  tri   P1_add_348_n196;
  tri   P1_add_348_n195;
  tri   P1_add_348_n194;
  tri   P1_add_348_n193;
  tri   P1_add_348_n192;
  tri   P1_add_348_n191;
  tri   P1_add_348_n189;
  tri   P1_add_348_n188;
  tri   P1_add_348_n187;
  tri   P1_add_348_n186;
  tri   P1_add_348_n185;
  tri   P1_add_348_n184;
  tri   P1_add_348_n183;
  tri   P1_add_348_n182;
  tri   P1_add_348_n181;
  tri   P1_add_348_n179;
  tri   P1_add_348_n178;
  tri   P1_add_348_n177;
  tri   P1_add_348_n176;
  tri   P1_add_348_n175;
  tri   P1_add_348_n174;
  tri   P1_add_348_n173;
  tri   P1_add_348_n172;
  tri   P1_add_348_n171;
  tri   P1_add_348_n169;
  tri   P1_add_348_n168;
  tri   P1_add_348_n167;
  tri   P1_add_348_n166;
  tri   P1_add_348_n165;
  tri   P1_add_348_n164;
  tri   P1_add_348_n163;
  tri   P1_add_348_n162;
  tri   P1_add_348_n161;
  tri   P1_add_348_n159;
  tri   P1_add_348_n158;
  tri   P1_add_348_n157;
  tri   P1_add_348_n156;
  tri   P1_add_348_n155;
  tri   P1_add_348_n153;
  tri   P1_add_348_n152;
  tri   P1_add_348_n150;
  tri   P1_add_348_n149;
  tri   P1_add_348_n148;
  tri   P1_add_348_n144;
  tri   P1_add_348_n147;
  tri   P1_add_348_n145;
  tri   P1_add_348_n146;
  tri   P1_add_348_n279;
  tri   P1_add_348_n278;
  tri   P1_add_348_n151;
  tri   P1_add_348_n277;
  tri   P1_add_348_n276;
  tri   P1_add_348_n275;
  tri   P1_add_348_n52;
  tri   P1_add_348_n274;
  tri   P1_add_348_n273;
  tri   P1_add_348_n272;
  tri   P1_add_348_n45;
  tri   P1_add_348_n271;
  tri   P1_add_348_n270;
  tri   P1_add_348_n269;
  tri   P1_add_348_n38;
  tri   P1_add_348_n268;
  tri   P1_add_348_n267;
  tri   P1_add_348_n266;
  tri   P1_add_348_n31;
  tri   P1_add_348_n265;
  tri   P1_add_348_n264;
  tri   P1_add_348_n263;
  tri   P1_add_348_n24;
  tri   P1_add_348_n262;
  tri   P1_add_348_n261;
  tri   P1_add_348_n260;
  tri   P1_add_348_n17;
  tri   P1_add_348_n259;
  tri   P1_add_348_n258;
  tri   P1_add_348_n257;
  tri   P1_add_348_n10;
  tri   P1_add_348_n256;
  tri   P1_add_348_n255;
  tri   P1_add_348_n254;
  tri   P1_add_348_n3;
  tri   P1_add_348_n253;
  tri   P1_add_348_n252;
  tri   P1_add_348_n251;
  tri   P1_add_348_n249;
  tri   P1_add_348_n248;
  tri   P1_add_348_n247;
  tri   P1_add_348_n246;
  tri   P1_add_348_n245;
  tri   P1_add_348_n244;
  tri   P1_add_348_n243;
  tri   P1_add_348_n242;
  tri   P1_add_348_n241;
  tri   P1_add_348_n239;
  tri   P1_add_348_n238;
  tri   P1_add_348_n237;
  tri   P1_add_348_n236;
  tri   P1_add_348_n235;
  tri   P1_add_348_n234;
  tri   P1_add_348_n233;
  tri   P1_add_348_n224;
  tri   P1_add_348_n232;
  tri   P1_add_348_n231;
  tri   P1_add_348_n93;
  tri   P1_add_348_n180;
  tri   P1_add_368_n86;
  tri   P1_add_368_n85;
  tri   P1_add_368_n84;
  tri   P1_add_368_n82;
  tri   P1_add_368_n81;
  tri   P1_add_368_n80;
  tri   P1_add_368_n79;
  tri   P1_add_368_n78;
  tri   P1_add_368_n77;
  tri   P1_add_368_n76;
  tri   P1_add_368_n75;
  tri   P1_add_368_n74;
  tri   P1_add_368_n72;
  tri   P1_add_368_n71;
  tri   P1_add_368_n70;
  tri   P1_add_368_n69;
  tri   P1_add_368_n68;
  tri   P1_add_368_n66;
  tri   P1_add_368_n65;
  tri   P1_add_368_n64;
  tri   P1_add_368_n63;
  tri   P1_add_368_n62;
  tri   P1_add_368_n61;
  tri   P1_add_368_n60;
  tri   P1_add_368_n59;
  tri   P1_add_368_n58;
  tri   P1_add_368_n57;
  tri   P1_add_368_n55;
  tri   P1_add_368_n54;
  tri   P1_add_368_n53;
  tri   P1_add_368_n51;
  tri   P1_add_368_n50;
  tri   P1_add_368_n48;
  tri   P1_add_368_n47;
  tri   P1_add_368_n46;
  tri   P1_add_368_n44;
  tri   P1_add_368_n43;
  tri   P1_add_368_n41;
  tri   P1_add_368_n40;
  tri   P1_add_368_n39;
  tri   P1_add_368_n37;
  tri   P1_add_368_n36;
  tri   P1_add_368_n34;
  tri   P1_add_368_n33;
  tri   P1_add_368_n32;
  tri   P1_add_368_n30;
  tri   P1_add_368_n29;
  tri   P1_add_368_n27;
  tri   P1_add_368_n26;
  tri   P1_add_368_n25;
  tri   P1_add_368_n23;
  tri   P1_add_368_n22;
  tri   P1_add_368_n20;
  tri   P1_add_368_n19;
  tri   P1_add_368_n18;
  tri   P1_add_368_n16;
  tri   P1_add_368_n15;
  tri   P1_add_368_n13;
  tri   P1_add_368_n12;
  tri   P1_add_368_n11;
  tri   P1_add_368_n9;
  tri   P1_add_368_n8;
  tri   P1_add_368_n6;
  tri   P1_add_368_n5;
  tri   P1_add_368_n4;
  tri   P1_add_368_n2;
  tri   P1_add_368_n1;
  tri   P1_add_368_n173;
  tri   P1_add_368_n172;
  tri   P1_add_368_n169;
  tri   P1_add_368_n168;
  tri   P1_add_368_n167;
  tri   P1_add_368_n166;
  tri   P1_add_368_n165;
  tri   P1_add_368_n164;
  tri   P1_add_368_n163;
  tri   P1_add_368_n162;
  tri   P1_add_368_n161;
  tri   P1_add_368_n159;
  tri   P1_add_368_n158;
  tri   P1_add_368_n157;
  tri   P1_add_368_n156;
  tri   P1_add_368_n155;
  tri   P1_add_368_n153;
  tri   P1_add_368_n152;
  tri   P1_add_368_n150;
  tri   P1_add_368_n149;
  tri   P1_add_368_n148;
  tri   P1_add_368_n147;
  tri   P1_add_368_n146;
  tri   P1_add_368_n145;
  tri   P1_add_368_n144;
  tri   P1_add_368_n142;
  tri   P1_add_368_n141;
  tri   P1_add_368_n140;
  tri   P1_add_368_n139;
  tri   P1_add_368_n138;
  tri   P1_add_368_n137;
  tri   P1_add_368_n136;
  tri   P1_add_368_n135;
  tri   P1_add_368_n134;
  tri   P1_add_368_n132;
  tri   P1_add_368_n131;
  tri   P1_add_368_n130;
  tri   P1_add_368_n129;
  tri   P1_add_368_n128;
  tri   P1_add_368_n127;
  tri   P1_add_368_n126;
  tri   P1_add_368_n125;
  tri   P1_add_368_n124;
  tri   P1_add_368_n122;
  tri   P1_add_368_n121;
  tri   P1_add_368_n120;
  tri   P1_add_368_n119;
  tri   P1_add_368_n118;
  tri   P1_add_368_n117;
  tri   P1_add_368_n116;
  tri   P1_add_368_n115;
  tri   P1_add_368_n114;
  tri   P1_add_368_n112;
  tri   P1_add_368_n111;
  tri   P1_add_368_n110;
  tri   P1_add_368_n109;
  tri   P1_add_368_n108;
  tri   P1_add_368_n107;
  tri   P1_add_368_n106;
  tri   P1_add_368_n105;
  tri   P1_add_368_n104;
  tri   P1_add_368_n102;
  tri   P1_add_368_n101;
  tri   P1_add_368_n100;
  tri   P1_add_368_n99;
  tri   P1_add_368_n98;
  tri   P1_add_368_n97;
  tri   P1_add_368_n96;
  tri   P1_add_368_n95;
  tri   P1_add_368_n94;
  tri   P1_add_368_n92;
  tri   P1_add_368_n91;
  tri   P1_add_368_n90;
  tri   P1_add_368_n87;
  tri   P1_add_368_n89;
  tri   P1_add_368_n88;
  tri   P1_add_368_n256;
  tri   P1_add_368_n255;
  tri   P1_add_368_n254;
  tri   P1_add_368_n3;
  tri   P1_add_368_n253;
  tri   P1_add_368_n252;
  tri   P1_add_368_n251;
  tri   P1_add_368_n249;
  tri   P1_add_368_n248;
  tri   P1_add_368_n247;
  tri   P1_add_368_n246;
  tri   P1_add_368_n245;
  tri   P1_add_368_n244;
  tri   P1_add_368_n243;
  tri   P1_add_368_n242;
  tri   P1_add_368_n241;
  tri   P1_add_368_n239;
  tri   P1_add_368_n238;
  tri   P1_add_368_n237;
  tri   P1_add_368_n236;
  tri   P1_add_368_n235;
  tri   P1_add_368_n234;
  tri   P1_add_368_n233;
  tri   P1_add_368_n232;
  tri   P1_add_368_n231;
  tri   P1_add_368_n229;
  tri   P1_add_368_n228;
  tri   P1_add_368_n227;
  tri   P1_add_368_n226;
  tri   P1_add_368_n225;
  tri   P1_add_368_n224;
  tri   P1_add_368_n223;
  tri   P1_add_368_n222;
  tri   P1_add_368_n221;
  tri   P1_add_368_n219;
  tri   P1_add_368_n218;
  tri   P1_add_368_n217;
  tri   P1_add_368_n216;
  tri   P1_add_368_n215;
  tri   P1_add_368_n214;
  tri   P1_add_368_n213;
  tri   P1_add_368_n212;
  tri   P1_add_368_n211;
  tri   P1_add_368_n209;
  tri   P1_add_368_n208;
  tri   P1_add_368_n207;
  tri   P1_add_368_n206;
  tri   P1_add_368_n205;
  tri   P1_add_368_n204;
  tri   P1_add_368_n203;
  tri   P1_add_368_n202;
  tri   P1_add_368_n201;
  tri   P1_add_368_n199;
  tri   P1_add_368_n198;
  tri   P1_add_368_n197;
  tri   P1_add_368_n196;
  tri   P1_add_368_n195;
  tri   P1_add_368_n194;
  tri   P1_add_368_n193;
  tri   P1_add_368_n192;
  tri   P1_add_368_n191;
  tri   P1_add_368_n189;
  tri   P1_add_368_n188;
  tri   P1_add_368_n187;
  tri   P1_add_368_n186;
  tri   P1_add_368_n185;
  tri   P1_add_368_n184;
  tri   P1_add_368_n183;
  tri   P1_add_368_n182;
  tri   P1_add_368_n181;
  tri   P1_add_368_n179;
  tri   P1_add_368_n178;
  tri   P1_add_368_n177;
  tri   P1_add_368_n176;
  tri   P1_add_368_n175;
  tri   P1_add_368_n171;
  tri   P1_add_368_n174;
  tri   P1_add_368_n279;
  tri   P1_add_368_n278;
  tri   P1_add_368_n151;
  tri   P1_add_368_n277;
  tri   P1_add_368_n276;
  tri   P1_add_368_n275;
  tri   P1_add_368_n52;
  tri   P1_add_368_n274;
  tri   P1_add_368_n273;
  tri   P1_add_368_n272;
  tri   P1_add_368_n45;
  tri   P1_add_368_n271;
  tri   P1_add_368_n270;
  tri   P1_add_368_n269;
  tri   P1_add_368_n38;
  tri   P1_add_368_n268;
  tri   P1_add_368_n267;
  tri   P1_add_368_n266;
  tri   P1_add_368_n31;
  tri   P1_add_368_n265;
  tri   P1_add_368_n264;
  tri   P1_add_368_n263;
  tri   P1_add_368_n24;
  tri   P1_add_368_n262;
  tri   P1_add_368_n261;
  tri   P1_add_368_n260;
  tri   P1_add_368_n17;
  tri   P1_add_368_n259;
  tri   P1_add_368_n10;
  tri   P1_add_368_n258;
  tri   P1_add_368_n257;
  tri   P1_sub_388_n30;
  tri   P1_sub_388_n29;
  tri   P1_sub_388_n27;
  tri   P1_sub_388_n26;
  tri   P1_sub_388_n24;
  tri   P1_sub_388_n23;
  tri   P1_sub_388_n22;
  tri   P1_sub_388_n20;
  tri   P1_sub_388_n19;
  tri   P1_sub_388_n17;
  tri   P1_sub_388_n16;
  tri   P1_sub_388_n15;
  tri   P1_sub_388_n13;
  tri   P1_sub_388_n12;
  tri   P1_sub_388_n10;
  tri   P1_sub_388_n9;
  tri   P1_sub_388_n8;
  tri   P1_sub_388_n6;
  tri   P1_sub_388_n5;
  tri   P1_sub_388_n3;
  tri   P1_sub_388_n2;
  tri   P1_sub_388_n1;
  tri   P1_sub_388_n124;
  tri   P1_sub_388_n123;
  tri   P1_sub_388_n120;
  tri   P1_sub_388_n119;
  tri   P1_sub_388_n118;
  tri   P1_sub_388_n117;
  tri   P1_sub_388_n116;
  tri   P1_sub_388_n114;
  tri   P1_sub_388_n113;
  tri   P1_sub_388_n112;
  tri   P1_sub_388_n111;
  tri   P1_sub_388_n110;
  tri   P1_sub_388_n109;
  tri   P1_sub_388_n108;
  tri   P1_sub_388_n107;
  tri   P1_sub_388_n106;
  tri   P1_sub_388_n105;
  tri   P1_sub_388_n104;
  tri   P1_sub_388_n103;
  tri   P1_sub_388_n102;
  tri   P1_sub_388_n101;
  tri   P1_sub_388_n100;
  tri   P1_sub_388_n99;
  tri   P1_sub_388_n98;
  tri   P1_sub_388_n97;
  tri   P1_sub_388_n96;
  tri   P1_sub_388_n95;
  tri   P1_sub_388_n94;
  tri   P1_sub_388_n93;
  tri   P1_sub_388_n92;
  tri   P1_sub_388_n91;
  tri   P1_sub_388_n90;
  tri   P1_sub_388_n89;
  tri   P1_sub_388_n88;
  tri   P1_sub_388_n87;
  tri   P1_sub_388_n86;
  tri   P1_sub_388_n85;
  tri   P1_sub_388_n84;
  tri   P1_sub_388_n83;
  tri   P1_sub_388_n82;
  tri   P1_sub_388_n81;
  tri   P1_sub_388_n80;
  tri   P1_sub_388_n79;
  tri   P1_sub_388_n78;
  tri   P1_sub_388_n77;
  tri   P1_sub_388_n76;
  tri   P1_sub_388_n75;
  tri   P1_sub_388_n74;
  tri   P1_sub_388_n73;
  tri   P1_sub_388_n72;
  tri   P1_sub_388_n71;
  tri   P1_sub_388_n70;
  tri   P1_sub_388_n69;
  tri   P1_sub_388_n67;
  tri   P1_sub_388_n66;
  tri   P1_sub_388_n65;
  tri   P1_sub_388_n64;
  tri   P1_sub_388_n63;
  tri   P1_sub_388_n62;
  tri   P1_sub_388_n61;
  tri   P1_sub_388_n59;
  tri   P1_sub_388_n60;
  tri   P1_sub_388_n58;
  tri   P1_sub_388_n57;
  tri   P1_sub_388_n55;
  tri   P1_sub_388_n54;
  tri   P1_sub_388_n52;
  tri   P1_sub_388_n51;
  tri   P1_sub_388_n50;
  tri   P1_sub_388_n48;
  tri   P1_sub_388_n47;
  tri   P1_sub_388_n45;
  tri   P1_sub_388_n44;
  tri   P1_sub_388_n43;
  tri   P1_sub_388_n41;
  tri   P1_sub_388_n40;
  tri   P1_sub_388_n38;
  tri   P1_sub_388_n37;
  tri   P1_sub_388_n36;
  tri   P1_sub_388_n31;
  tri   P1_sub_388_n34;
  tri   P1_sub_388_n33;
  tri   P1_sub_388_n211;
  tri   P1_sub_388_n208;
  tri   P1_sub_388_n207;
  tri   P1_sub_388_n206;
  tri   P1_sub_388_n205;
  tri   P1_sub_388_n204;
  tri   P1_sub_388_n202;
  tri   P1_sub_388_n201;
  tri   P1_sub_388_n200;
  tri   P1_sub_388_n199;
  tri   P1_sub_388_n198;
  tri   P1_sub_388_n197;
  tri   P1_sub_388_n196;
  tri   P1_sub_388_n195;
  tri   P1_sub_388_n194;
  tri   P1_sub_388_n193;
  tri   P1_sub_388_n192;
  tri   P1_sub_388_n191;
  tri   P1_sub_388_n190;
  tri   P1_sub_388_n189;
  tri   P1_sub_388_n188;
  tri   P1_sub_388_n187;
  tri   P1_sub_388_n186;
  tri   P1_sub_388_n185;
  tri   P1_sub_388_n184;
  tri   P1_sub_388_n183;
  tri   P1_sub_388_n182;
  tri   P1_sub_388_n181;
  tri   P1_sub_388_n180;
  tri   P1_sub_388_n179;
  tri   P1_sub_388_n178;
  tri   P1_sub_388_n177;
  tri   P1_sub_388_n176;
  tri   P1_sub_388_n175;
  tri   P1_sub_388_n174;
  tri   P1_sub_388_n173;
  tri   P1_sub_388_n172;
  tri   P1_sub_388_n171;
  tri   P1_sub_388_n170;
  tri   P1_sub_388_n169;
  tri   P1_sub_388_n168;
  tri   P1_sub_388_n167;
  tri   P1_sub_388_n166;
  tri   P1_sub_388_n165;
  tri   P1_sub_388_n164;
  tri   P1_sub_388_n163;
  tri   P1_sub_388_n162;
  tri   P1_sub_388_n161;
  tri   P1_sub_388_n160;
  tri   P1_sub_388_n159;
  tri   P1_sub_388_n158;
  tri   P1_sub_388_n157;
  tri   P1_sub_388_n154;
  tri   P1_sub_388_n153;
  tri   P1_sub_388_n151;
  tri   P1_sub_388_n150;
  tri   P1_sub_388_n149;
  tri   P1_sub_388_n148;
  tri   P1_sub_388_n147;
  tri   P1_sub_388_n146;
  tri   P1_sub_388_n145;
  tri   P1_sub_388_n144;
  tri   P1_sub_388_n143;
  tri   P1_sub_388_n142;
  tri   P1_sub_388_n141;
  tri   P1_sub_388_n140;
  tri   P1_sub_388_n139;
  tri   P1_sub_388_n125;
  tri   P1_sub_388_n138;
  tri   P1_sub_388_n137;
  tri   P1_sub_388_n136;
  tri   P1_sub_388_n135;
  tri   P1_sub_388_n134;
  tri   P1_sub_388_n133;
  tri   P1_sub_388_n132;
  tri   P1_sub_388_n131;
  tri   P1_sub_388_n130;
  tri   P1_sub_388_n129;
  tri   P1_sub_388_n115;
  tri   P1_sub_388_n121;
  tri   P1_sub_388_n128;
  tri   P1_sub_388_n127;
  tri   P1_sub_388_n122;
  tri   P1_sub_388_n126;
  tri   P1_sub_388_n279;
  tri   P1_sub_388_n278;
  tri   P1_sub_388_n156;
  tri   P1_sub_388_n276;
  tri   P1_sub_388_n275;
  tri   P1_sub_388_n274;
  tri   P1_sub_388_n53;
  tri   P1_sub_388_n56;
  tri   P1_sub_388_n273;
  tri   P1_sub_388_n272;
  tri   P1_sub_388_n271;
  tri   P1_sub_388_n46;
  tri   P1_sub_388_n49;
  tri   P1_sub_388_n270;
  tri   P1_sub_388_n269;
  tri   P1_sub_388_n268;
  tri   P1_sub_388_n39;
  tri   P1_sub_388_n42;
  tri   P1_sub_388_n267;
  tri   P1_sub_388_n266;
  tri   P1_sub_388_n265;
  tri   P1_sub_388_n32;
  tri   P1_sub_388_n35;
  tri   P1_sub_388_n264;
  tri   P1_sub_388_n263;
  tri   P1_sub_388_n262;
  tri   P1_sub_388_n25;
  tri   P1_sub_388_n28;
  tri   P1_sub_388_n261;
  tri   P1_sub_388_n260;
  tri   P1_sub_388_n259;
  tri   P1_sub_388_n18;
  tri   P1_sub_388_n21;
  tri   P1_sub_388_n258;
  tri   P1_sub_388_n257;
  tri   P1_sub_388_n256;
  tri   P1_sub_388_n11;
  tri   P1_sub_388_n14;
  tri   P1_sub_388_n255;
  tri   P1_sub_388_n254;
  tri   P1_sub_388_n253;
  tri   P1_sub_388_n4;
  tri   P1_sub_388_n7;
  tri   P1_sub_388_n252;
  tri   P1_sub_388_n251;
  tri   P1_sub_388_n250;
  tri   P1_sub_388_n249;
  tri   P1_sub_388_n248;
  tri   P1_sub_388_n247;
  tri   P1_sub_388_n246;
  tri   P1_sub_388_n245;
  tri   P1_sub_388_n244;
  tri   P1_sub_388_n243;
  tri   P1_sub_388_n242;
  tri   P1_sub_388_n241;
  tri   P1_sub_388_n240;
  tri   P1_sub_388_n239;
  tri   P1_sub_388_n238;
  tri   P1_sub_388_n237;
  tri   P1_sub_388_n236;
  tri   P1_sub_388_n235;
  tri   P1_sub_388_n234;
  tri   P1_sub_388_n233;
  tri   P1_sub_388_n232;
  tri   P1_sub_388_n231;
  tri   P1_sub_388_n230;
  tri   P1_sub_388_n229;
  tri   P1_sub_388_n228;
  tri   P1_sub_388_n227;
  tri   P1_sub_388_n213;
  tri   P1_sub_388_n226;
  tri   P1_sub_388_n225;
  tri   P1_sub_388_n224;
  tri   P1_sub_388_n223;
  tri   P1_sub_388_n222;
  tri   P1_sub_388_n221;
  tri   P1_sub_388_n220;
  tri   P1_sub_388_n219;
  tri   P1_sub_388_n218;
  tri   P1_sub_388_n217;
  tri   P1_sub_388_n203;
  tri   P1_sub_388_n209;
  tri   P1_sub_388_n216;
  tri   P1_sub_388_n215;
  tri   P1_sub_388_n210;
  tri   P1_sub_388_n212;
  tri   P1_sub_388_n214;
  tri   P1_sub_388_n277;
  tri   P1_sub_388_n152;
  tri   P1_sub_388_n280;
  tri   P1_sub_388_n281;
  tri   P1_sub_408_n67;
  tri   P1_sub_408_n66;
  tri   P1_sub_408_n63;
  tri   P1_sub_408_n62;
  tri   P1_sub_408_n61;
  tri   P1_sub_408_n59;
  tri   P1_sub_408_n60;
  tri   P1_sub_408_n58;
  tri   P1_sub_408_n57;
  tri   P1_sub_408_n55;
  tri   P1_sub_408_n54;
  tri   P1_sub_408_n52;
  tri   P1_sub_408_n51;
  tri   P1_sub_408_n50;
  tri   P1_sub_408_n48;
  tri   P1_sub_408_n47;
  tri   P1_sub_408_n45;
  tri   P1_sub_408_n44;
  tri   P1_sub_408_n43;
  tri   P1_sub_408_n41;
  tri   P1_sub_408_n40;
  tri   P1_sub_408_n38;
  tri   P1_sub_408_n37;
  tri   P1_sub_408_n36;
  tri   P1_sub_408_n34;
  tri   P1_sub_408_n33;
  tri   P1_sub_408_n31;
  tri   P1_sub_408_n30;
  tri   P1_sub_408_n29;
  tri   P1_sub_408_n27;
  tri   P1_sub_408_n26;
  tri   P1_sub_408_n24;
  tri   P1_sub_408_n23;
  tri   P1_sub_408_n22;
  tri   P1_sub_408_n20;
  tri   P1_sub_408_n19;
  tri   P1_sub_408_n17;
  tri   P1_sub_408_n16;
  tri   P1_sub_408_n15;
  tri   P1_sub_408_n13;
  tri   P1_sub_408_n12;
  tri   P1_sub_408_n10;
  tri   P1_sub_408_n9;
  tri   P1_sub_408_n8;
  tri   P1_sub_408_n6;
  tri   P1_sub_408_n5;
  tri   P1_sub_408_n3;
  tri   P1_sub_408_n2;
  tri   P1_sub_408_n1;
  tri   P1_sub_408_n151;
  tri   P1_sub_408_n150;
  tri   P1_sub_408_n149;
  tri   P1_sub_408_n148;
  tri   P1_sub_408_n147;
  tri   P1_sub_408_n144;
  tri   P1_sub_408_n143;
  tri   P1_sub_408_n142;
  tri   P1_sub_408_n141;
  tri   P1_sub_408_n140;
  tri   P1_sub_408_n139;
  tri   P1_sub_408_n138;
  tri   P1_sub_408_n137;
  tri   P1_sub_408_n136;
  tri   P1_sub_408_n135;
  tri   P1_sub_408_n134;
  tri   P1_sub_408_n133;
  tri   P1_sub_408_n132;
  tri   P1_sub_408_n131;
  tri   P1_sub_408_n130;
  tri   P1_sub_408_n129;
  tri   P1_sub_408_n128;
  tri   P1_sub_408_n127;
  tri   P1_sub_408_n126;
  tri   P1_sub_408_n125;
  tri   P1_sub_408_n124;
  tri   P1_sub_408_n123;
  tri   P1_sub_408_n122;
  tri   P1_sub_408_n121;
  tri   P1_sub_408_n120;
  tri   P1_sub_408_n119;
  tri   P1_sub_408_n118;
  tri   P1_sub_408_n117;
  tri   P1_sub_408_n116;
  tri   P1_sub_408_n115;
  tri   P1_sub_408_n114;
  tri   P1_sub_408_n113;
  tri   P1_sub_408_n112;
  tri   P1_sub_408_n111;
  tri   P1_sub_408_n110;
  tri   P1_sub_408_n109;
  tri   P1_sub_408_n108;
  tri   P1_sub_408_n107;
  tri   P1_sub_408_n106;
  tri   P1_sub_408_n105;
  tri   P1_sub_408_n104;
  tri   P1_sub_408_n103;
  tri   P1_sub_408_n102;
  tri   P1_sub_408_n101;
  tri   P1_sub_408_n100;
  tri   P1_sub_408_n99;
  tri   P1_sub_408_n98;
  tri   P1_sub_408_n97;
  tri   P1_sub_408_n96;
  tri   P1_sub_408_n95;
  tri   P1_sub_408_n94;
  tri   P1_sub_408_n93;
  tri   P1_sub_408_n92;
  tri   P1_sub_408_n91;
  tri   P1_sub_408_n90;
  tri   P1_sub_408_n89;
  tri   P1_sub_408_n88;
  tri   P1_sub_408_n87;
  tri   P1_sub_408_n86;
  tri   P1_sub_408_n85;
  tri   P1_sub_408_n84;
  tri   P1_sub_408_n83;
  tri   P1_sub_408_n82;
  tri   P1_sub_408_n81;
  tri   P1_sub_408_n80;
  tri   P1_sub_408_n79;
  tri   P1_sub_408_n64;
  tri   P1_sub_408_n78;
  tri   P1_sub_408_n77;
  tri   P1_sub_408_n76;
  tri   P1_sub_408_n75;
  tri   P1_sub_408_n74;
  tri   P1_sub_408_n73;
  tri   P1_sub_408_n72;
  tri   P1_sub_408_n71;
  tri   P1_sub_408_n65;
  tri   P1_sub_408_n70;
  tri   P1_sub_408_n69;
  tri   P1_sub_408_n238;
  tri   P1_sub_408_n237;
  tri   P1_sub_408_n236;
  tri   P1_sub_408_n235;
  tri   P1_sub_408_n232;
  tri   P1_sub_408_n231;
  tri   P1_sub_408_n230;
  tri   P1_sub_408_n229;
  tri   P1_sub_408_n228;
  tri   P1_sub_408_n227;
  tri   P1_sub_408_n226;
  tri   P1_sub_408_n225;
  tri   P1_sub_408_n224;
  tri   P1_sub_408_n223;
  tri   P1_sub_408_n222;
  tri   P1_sub_408_n221;
  tri   P1_sub_408_n220;
  tri   P1_sub_408_n219;
  tri   P1_sub_408_n218;
  tri   P1_sub_408_n217;
  tri   P1_sub_408_n216;
  tri   P1_sub_408_n215;
  tri   P1_sub_408_n214;
  tri   P1_sub_408_n213;
  tri   P1_sub_408_n212;
  tri   P1_sub_408_n211;
  tri   P1_sub_408_n210;
  tri   P1_sub_408_n209;
  tri   P1_sub_408_n208;
  tri   P1_sub_408_n207;
  tri   P1_sub_408_n206;
  tri   P1_sub_408_n205;
  tri   P1_sub_408_n204;
  tri   P1_sub_408_n203;
  tri   P1_sub_408_n202;
  tri   P1_sub_408_n201;
  tri   P1_sub_408_n200;
  tri   P1_sub_408_n199;
  tri   P1_sub_408_n198;
  tri   P1_sub_408_n197;
  tri   P1_sub_408_n196;
  tri   P1_sub_408_n195;
  tri   P1_sub_408_n194;
  tri   P1_sub_408_n193;
  tri   P1_sub_408_n192;
  tri   P1_sub_408_n191;
  tri   P1_sub_408_n190;
  tri   P1_sub_408_n189;
  tri   P1_sub_408_n188;
  tri   P1_sub_408_n187;
  tri   P1_sub_408_n186;
  tri   P1_sub_408_n185;
  tri   P1_sub_408_n184;
  tri   P1_sub_408_n183;
  tri   P1_sub_408_n182;
  tri   P1_sub_408_n181;
  tri   P1_sub_408_n180;
  tri   P1_sub_408_n179;
  tri   P1_sub_408_n178;
  tri   P1_sub_408_n177;
  tri   P1_sub_408_n176;
  tri   P1_sub_408_n175;
  tri   P1_sub_408_n174;
  tri   P1_sub_408_n173;
  tri   P1_sub_408_n172;
  tri   P1_sub_408_n171;
  tri   P1_sub_408_n170;
  tri   P1_sub_408_n169;
  tri   P1_sub_408_n168;
  tri   P1_sub_408_n167;
  tri   P1_sub_408_n145;
  tri   P1_sub_408_n166;
  tri   P1_sub_408_n165;
  tri   P1_sub_408_n164;
  tri   P1_sub_408_n163;
  tri   P1_sub_408_n162;
  tri   P1_sub_408_n161;
  tri   P1_sub_408_n160;
  tri   P1_sub_408_n159;
  tri   P1_sub_408_n146;
  tri   P1_sub_408_n158;
  tri   P1_sub_408_n157;
  tri   P1_sub_408_n153;
  tri   P1_sub_408_n154;
  tri   P1_sub_408_n281;
  tri   P1_sub_408_n280;
  tri   P1_sub_408_n279;
  tri   P1_sub_408_n278;
  tri   P1_sub_408_n152;
  tri   P1_sub_408_n277;
  tri   P1_sub_408_n156;
  tri   P1_sub_408_n276;
  tri   P1_sub_408_n275;
  tri   P1_sub_408_n274;
  tri   P1_sub_408_n53;
  tri   P1_sub_408_n56;
  tri   P1_sub_408_n273;
  tri   P1_sub_408_n272;
  tri   P1_sub_408_n271;
  tri   P1_sub_408_n46;
  tri   P1_sub_408_n49;
  tri   P1_sub_408_n270;
  tri   P1_sub_408_n269;
  tri   P1_sub_408_n268;
  tri   P1_sub_408_n39;
  tri   P1_sub_408_n42;
  tri   P1_sub_408_n267;
  tri   P1_sub_408_n266;
  tri   P1_sub_408_n265;
  tri   P1_sub_408_n32;
  tri   P1_sub_408_n35;
  tri   P1_sub_408_n264;
  tri   P1_sub_408_n263;
  tri   P1_sub_408_n262;
  tri   P1_sub_408_n25;
  tri   P1_sub_408_n28;
  tri   P1_sub_408_n261;
  tri   P1_sub_408_n260;
  tri   P1_sub_408_n259;
  tri   P1_sub_408_n18;
  tri   P1_sub_408_n21;
  tri   P1_sub_408_n258;
  tri   P1_sub_408_n257;
  tri   P1_sub_408_n256;
  tri   P1_sub_408_n11;
  tri   P1_sub_408_n14;
  tri   P1_sub_408_n255;
  tri   P1_sub_408_n254;
  tri   P1_sub_408_n253;
  tri   P1_sub_408_n4;
  tri   P1_sub_408_n7;
  tri   P1_sub_408_n252;
  tri   P1_sub_408_n251;
  tri   P1_sub_408_n250;
  tri   P1_sub_408_n249;
  tri   P1_sub_408_n248;
  tri   P1_sub_408_n247;
  tri   P1_sub_408_n233;
  tri   P1_sub_408_n239;
  tri   P1_sub_408_n246;
  tri   P1_sub_408_n245;
  tri   P1_sub_408_n244;
  tri   P1_sub_408_n243;
  tri   P1_sub_408_n242;
  tri   P1_sub_408_n234;
  tri   P1_sub_408_n241;
  tri   P1_sub_408_n240;
  tri   P1_add_428_n86;
  tri   P1_add_428_n85;
  tri   P1_add_428_n82;
  tri   P1_add_428_n81;
  tri   P1_add_428_n80;
  tri   P1_add_428_n79;
  tri   P1_add_428_n78;
  tri   P1_add_428_n77;
  tri   P1_add_428_n76;
  tri   P1_add_428_n75;
  tri   P1_add_428_n74;
  tri   P1_add_428_n72;
  tri   P1_add_428_n71;
  tri   P1_add_428_n70;
  tri   P1_add_428_n69;
  tri   P1_add_428_n68;
  tri   P1_add_428_n66;
  tri   P1_add_428_n65;
  tri   P1_add_428_n64;
  tri   P1_add_428_n63;
  tri   P1_add_428_n62;
  tri   P1_add_428_n61;
  tri   P1_add_428_n60;
  tri   P1_add_428_n59;
  tri   P1_add_428_n58;
  tri   P1_add_428_n57;
  tri   P1_add_428_n55;
  tri   P1_add_428_n54;
  tri   P1_add_428_n53;
  tri   P1_add_428_n51;
  tri   P1_add_428_n50;
  tri   P1_add_428_n48;
  tri   P1_add_428_n47;
  tri   P1_add_428_n46;
  tri   P1_add_428_n44;
  tri   P1_add_428_n43;
  tri   P1_add_428_n41;
  tri   P1_add_428_n40;
  tri   P1_add_428_n39;
  tri   P1_add_428_n37;
  tri   P1_add_428_n36;
  tri   P1_add_428_n34;
  tri   P1_add_428_n33;
  tri   P1_add_428_n32;
  tri   P1_add_428_n30;
  tri   P1_add_428_n29;
  tri   P1_add_428_n27;
  tri   P1_add_428_n26;
  tri   P1_add_428_n25;
  tri   P1_add_428_n23;
  tri   P1_add_428_n22;
  tri   P1_add_428_n20;
  tri   P1_add_428_n19;
  tri   P1_add_428_n18;
  tri   P1_add_428_n16;
  tri   P1_add_428_n15;
  tri   P1_add_428_n13;
  tri   P1_add_428_n12;
  tri   P1_add_428_n11;
  tri   P1_add_428_n9;
  tri   P1_add_428_n8;
  tri   P1_add_428_n6;
  tri   P1_add_428_n5;
  tri   P1_add_428_n4;
  tri   P1_add_428_n2;
  tri   P1_add_428_n1;
  tri   P1_add_428_n172;
  tri   P1_add_428_n169;
  tri   P1_add_428_n168;
  tri   P1_add_428_n167;
  tri   P1_add_428_n166;
  tri   P1_add_428_n165;
  tri   P1_add_428_n164;
  tri   P1_add_428_n163;
  tri   P1_add_428_n162;
  tri   P1_add_428_n161;
  tri   P1_add_428_n159;
  tri   P1_add_428_n158;
  tri   P1_add_428_n157;
  tri   P1_add_428_n156;
  tri   P1_add_428_n155;
  tri   P1_add_428_n153;
  tri   P1_add_428_n152;
  tri   P1_add_428_n150;
  tri   P1_add_428_n149;
  tri   P1_add_428_n148;
  tri   P1_add_428_n147;
  tri   P1_add_428_n146;
  tri   P1_add_428_n145;
  tri   P1_add_428_n144;
  tri   P1_add_428_n142;
  tri   P1_add_428_n141;
  tri   P1_add_428_n140;
  tri   P1_add_428_n139;
  tri   P1_add_428_n138;
  tri   P1_add_428_n137;
  tri   P1_add_428_n136;
  tri   P1_add_428_n135;
  tri   P1_add_428_n134;
  tri   P1_add_428_n132;
  tri   P1_add_428_n131;
  tri   P1_add_428_n130;
  tri   P1_add_428_n129;
  tri   P1_add_428_n128;
  tri   P1_add_428_n127;
  tri   P1_add_428_n126;
  tri   P1_add_428_n125;
  tri   P1_add_428_n124;
  tri   P1_add_428_n122;
  tri   P1_add_428_n121;
  tri   P1_add_428_n120;
  tri   P1_add_428_n119;
  tri   P1_add_428_n118;
  tri   P1_add_428_n117;
  tri   P1_add_428_n116;
  tri   P1_add_428_n115;
  tri   P1_add_428_n114;
  tri   P1_add_428_n112;
  tri   P1_add_428_n111;
  tri   P1_add_428_n110;
  tri   P1_add_428_n109;
  tri   P1_add_428_n108;
  tri   P1_add_428_n107;
  tri   P1_add_428_n106;
  tri   P1_add_428_n105;
  tri   P1_add_428_n104;
  tri   P1_add_428_n102;
  tri   P1_add_428_n101;
  tri   P1_add_428_n100;
  tri   P1_add_428_n99;
  tri   P1_add_428_n98;
  tri   P1_add_428_n97;
  tri   P1_add_428_n96;
  tri   P1_add_428_n95;
  tri   P1_add_428_n94;
  tri   P1_add_428_n92;
  tri   P1_add_428_n91;
  tri   P1_add_428_n90;
  tri   P1_add_428_n89;
  tri   P1_add_428_n88;
  tri   P1_add_428_n84;
  tri   P1_add_428_n87;
  tri   P1_add_428_n256;
  tri   P1_add_428_n255;
  tri   P1_add_428_n3;
  tri   P1_add_428_n253;
  tri   P1_add_428_n252;
  tri   P1_add_428_n251;
  tri   P1_add_428_n249;
  tri   P1_add_428_n248;
  tri   P1_add_428_n247;
  tri   P1_add_428_n246;
  tri   P1_add_428_n245;
  tri   P1_add_428_n244;
  tri   P1_add_428_n243;
  tri   P1_add_428_n242;
  tri   P1_add_428_n241;
  tri   P1_add_428_n239;
  tri   P1_add_428_n238;
  tri   P1_add_428_n237;
  tri   P1_add_428_n236;
  tri   P1_add_428_n235;
  tri   P1_add_428_n234;
  tri   P1_add_428_n233;
  tri   P1_add_428_n232;
  tri   P1_add_428_n231;
  tri   P1_add_428_n229;
  tri   P1_add_428_n228;
  tri   P1_add_428_n227;
  tri   P1_add_428_n226;
  tri   P1_add_428_n225;
  tri   P1_add_428_n224;
  tri   P1_add_428_n223;
  tri   P1_add_428_n222;
  tri   P1_add_428_n221;
  tri   P1_add_428_n219;
  tri   P1_add_428_n218;
  tri   P1_add_428_n217;
  tri   P1_add_428_n216;
  tri   P1_add_428_n215;
  tri   P1_add_428_n214;
  tri   P1_add_428_n213;
  tri   P1_add_428_n212;
  tri   P1_add_428_n211;
  tri   P1_add_428_n209;
  tri   P1_add_428_n208;
  tri   P1_add_428_n207;
  tri   P1_add_428_n206;
  tri   P1_add_428_n205;
  tri   P1_add_428_n204;
  tri   P1_add_428_n203;
  tri   P1_add_428_n202;
  tri   P1_add_428_n201;
  tri   P1_add_428_n199;
  tri   P1_add_428_n198;
  tri   P1_add_428_n197;
  tri   P1_add_428_n196;
  tri   P1_add_428_n195;
  tri   P1_add_428_n194;
  tri   P1_add_428_n193;
  tri   P1_add_428_n192;
  tri   P1_add_428_n191;
  tri   P1_add_428_n189;
  tri   P1_add_428_n188;
  tri   P1_add_428_n187;
  tri   P1_add_428_n186;
  tri   P1_add_428_n185;
  tri   P1_add_428_n184;
  tri   P1_add_428_n183;
  tri   P1_add_428_n182;
  tri   P1_add_428_n181;
  tri   P1_add_428_n179;
  tri   P1_add_428_n178;
  tri   P1_add_428_n177;
  tri   P1_add_428_n176;
  tri   P1_add_428_n175;
  tri   P1_add_428_n171;
  tri   P1_add_428_n173;
  tri   P1_add_428_n174;
  tri   P1_add_428_n279;
  tri   P1_add_428_n278;
  tri   P1_add_428_n151;
  tri   P1_add_428_n277;
  tri   P1_add_428_n276;
  tri   P1_add_428_n275;
  tri   P1_add_428_n52;
  tri   P1_add_428_n274;
  tri   P1_add_428_n273;
  tri   P1_add_428_n272;
  tri   P1_add_428_n45;
  tri   P1_add_428_n271;
  tri   P1_add_428_n270;
  tri   P1_add_428_n269;
  tri   P1_add_428_n38;
  tri   P1_add_428_n268;
  tri   P1_add_428_n267;
  tri   P1_add_428_n266;
  tri   P1_add_428_n31;
  tri   P1_add_428_n265;
  tri   P1_add_428_n264;
  tri   P1_add_428_n263;
  tri   P1_add_428_n24;
  tri   P1_add_428_n262;
  tri   P1_add_428_n261;
  tri   P1_add_428_n260;
  tri   P1_add_428_n17;
  tri   P1_add_428_n259;
  tri   P1_add_428_n258;
  tri   P1_add_428_n257;
  tri   P1_add_428_n254;
  tri   P1_add_428_n10;
  tri   P1_sub_448_n30;
  tri   P1_sub_448_n27;
  tri   P1_sub_448_n26;
  tri   P1_sub_448_n24;
  tri   P1_sub_448_n23;
  tri   P1_sub_448_n22;
  tri   P1_sub_448_n20;
  tri   P1_sub_448_n19;
  tri   P1_sub_448_n17;
  tri   P1_sub_448_n16;
  tri   P1_sub_448_n15;
  tri   P1_sub_448_n13;
  tri   P1_sub_448_n12;
  tri   P1_sub_448_n10;
  tri   P1_sub_448_n9;
  tri   P1_sub_448_n8;
  tri   P1_sub_448_n6;
  tri   P1_sub_448_n5;
  tri   P1_sub_448_n3;
  tri   P1_sub_448_n2;
  tri   P1_sub_448_n1;
  tri   P1_sub_448_n123;
  tri   P1_sub_448_n120;
  tri   P1_sub_448_n119;
  tri   P1_sub_448_n118;
  tri   P1_sub_448_n117;
  tri   P1_sub_448_n116;
  tri   P1_sub_448_n114;
  tri   P1_sub_448_n113;
  tri   P1_sub_448_n112;
  tri   P1_sub_448_n111;
  tri   P1_sub_448_n110;
  tri   P1_sub_448_n109;
  tri   P1_sub_448_n108;
  tri   P1_sub_448_n107;
  tri   P1_sub_448_n106;
  tri   P1_sub_448_n105;
  tri   P1_sub_448_n104;
  tri   P1_sub_448_n103;
  tri   P1_sub_448_n102;
  tri   P1_sub_448_n101;
  tri   P1_sub_448_n100;
  tri   P1_sub_448_n99;
  tri   P1_sub_448_n98;
  tri   P1_sub_448_n97;
  tri   P1_sub_448_n96;
  tri   P1_sub_448_n95;
  tri   P1_sub_448_n94;
  tri   P1_sub_448_n93;
  tri   P1_sub_448_n92;
  tri   P1_sub_448_n91;
  tri   P1_sub_448_n90;
  tri   P1_sub_448_n89;
  tri   P1_sub_448_n88;
  tri   P1_sub_448_n87;
  tri   P1_sub_448_n86;
  tri   P1_sub_448_n85;
  tri   P1_sub_448_n84;
  tri   P1_sub_448_n83;
  tri   P1_sub_448_n82;
  tri   P1_sub_448_n81;
  tri   P1_sub_448_n80;
  tri   P1_sub_448_n79;
  tri   P1_sub_448_n78;
  tri   P1_sub_448_n77;
  tri   P1_sub_448_n76;
  tri   P1_sub_448_n75;
  tri   P1_sub_448_n74;
  tri   P1_sub_448_n73;
  tri   P1_sub_448_n72;
  tri   P1_sub_448_n71;
  tri   P1_sub_448_n70;
  tri   P1_sub_448_n69;
  tri   P1_sub_448_n67;
  tri   P1_sub_448_n66;
  tri   P1_sub_448_n65;
  tri   P1_sub_448_n64;
  tri   P1_sub_448_n63;
  tri   P1_sub_448_n62;
  tri   P1_sub_448_n61;
  tri   P1_sub_448_n59;
  tri   P1_sub_448_n60;
  tri   P1_sub_448_n58;
  tri   P1_sub_448_n57;
  tri   P1_sub_448_n55;
  tri   P1_sub_448_n54;
  tri   P1_sub_448_n52;
  tri   P1_sub_448_n51;
  tri   P1_sub_448_n50;
  tri   P1_sub_448_n48;
  tri   P1_sub_448_n47;
  tri   P1_sub_448_n45;
  tri   P1_sub_448_n44;
  tri   P1_sub_448_n43;
  tri   P1_sub_448_n41;
  tri   P1_sub_448_n40;
  tri   P1_sub_448_n38;
  tri   P1_sub_448_n37;
  tri   P1_sub_448_n36;
  tri   P1_sub_448_n34;
  tri   P1_sub_448_n33;
  tri   P1_sub_448_n29;
  tri   P1_sub_448_n31;
  tri   P1_sub_448_n208;
  tri   P1_sub_448_n207;
  tri   P1_sub_448_n206;
  tri   P1_sub_448_n205;
  tri   P1_sub_448_n204;
  tri   P1_sub_448_n202;
  tri   P1_sub_448_n201;
  tri   P1_sub_448_n200;
  tri   P1_sub_448_n199;
  tri   P1_sub_448_n198;
  tri   P1_sub_448_n197;
  tri   P1_sub_448_n196;
  tri   P1_sub_448_n195;
  tri   P1_sub_448_n194;
  tri   P1_sub_448_n193;
  tri   P1_sub_448_n192;
  tri   P1_sub_448_n191;
  tri   P1_sub_448_n190;
  tri   P1_sub_448_n189;
  tri   P1_sub_448_n188;
  tri   P1_sub_448_n187;
  tri   P1_sub_448_n186;
  tri   P1_sub_448_n185;
  tri   P1_sub_448_n184;
  tri   P1_sub_448_n183;
  tri   P1_sub_448_n182;
  tri   P1_sub_448_n181;
  tri   P1_sub_448_n180;
  tri   P1_sub_448_n179;
  tri   P1_sub_448_n178;
  tri   P1_sub_448_n177;
  tri   P1_sub_448_n176;
  tri   P1_sub_448_n175;
  tri   P1_sub_448_n174;
  tri   P1_sub_448_n173;
  tri   P1_sub_448_n172;
  tri   P1_sub_448_n171;
  tri   P1_sub_448_n170;
  tri   P1_sub_448_n169;
  tri   P1_sub_448_n168;
  tri   P1_sub_448_n167;
  tri   P1_sub_448_n166;
  tri   P1_sub_448_n165;
  tri   P1_sub_448_n164;
  tri   P1_sub_448_n163;
  tri   P1_sub_448_n162;
  tri   P1_sub_448_n161;
  tri   P1_sub_448_n160;
  tri   P1_sub_448_n159;
  tri   P1_sub_448_n158;
  tri   P1_sub_448_n157;
  tri   P1_sub_448_n154;
  tri   P1_sub_448_n153;
  tri   P1_sub_448_n151;
  tri   P1_sub_448_n150;
  tri   P1_sub_448_n149;
  tri   P1_sub_448_n148;
  tri   P1_sub_448_n147;
  tri   P1_sub_448_n146;
  tri   P1_sub_448_n145;
  tri   P1_sub_448_n144;
  tri   P1_sub_448_n143;
  tri   P1_sub_448_n142;
  tri   P1_sub_448_n141;
  tri   P1_sub_448_n140;
  tri   P1_sub_448_n139;
  tri   P1_sub_448_n125;
  tri   P1_sub_448_n138;
  tri   P1_sub_448_n137;
  tri   P1_sub_448_n136;
  tri   P1_sub_448_n135;
  tri   P1_sub_448_n134;
  tri   P1_sub_448_n133;
  tri   P1_sub_448_n132;
  tri   P1_sub_448_n131;
  tri   P1_sub_448_n130;
  tri   P1_sub_448_n129;
  tri   P1_sub_448_n115;
  tri   P1_sub_448_n121;
  tri   P1_sub_448_n128;
  tri   P1_sub_448_n127;
  tri   P1_sub_448_n122;
  tri   P1_sub_448_n124;
  tri   P1_sub_448_n126;
  tri   P1_sub_448_n279;
  tri   P1_sub_448_n278;
  tri   P1_sub_448_n156;
  tri   P1_sub_448_n276;
  tri   P1_sub_448_n275;
  tri   P1_sub_448_n274;
  tri   P1_sub_448_n53;
  tri   P1_sub_448_n56;
  tri   P1_sub_448_n273;
  tri   P1_sub_448_n272;
  tri   P1_sub_448_n271;
  tri   P1_sub_448_n46;
  tri   P1_sub_448_n49;
  tri   P1_sub_448_n270;
  tri   P1_sub_448_n269;
  tri   P1_sub_448_n268;
  tri   P1_sub_448_n39;
  tri   P1_sub_448_n42;
  tri   P1_sub_448_n267;
  tri   P1_sub_448_n266;
  tri   P1_sub_448_n265;
  tri   P1_sub_448_n32;
  tri   P1_sub_448_n35;
  tri   P1_sub_448_n264;
  tri   P1_sub_448_n263;
  tri   P1_sub_448_n262;
  tri   P1_sub_448_n25;
  tri   P1_sub_448_n28;
  tri   P1_sub_448_n261;
  tri   P1_sub_448_n260;
  tri   P1_sub_448_n259;
  tri   P1_sub_448_n18;
  tri   P1_sub_448_n21;
  tri   P1_sub_448_n258;
  tri   P1_sub_448_n257;
  tri   P1_sub_448_n256;
  tri   P1_sub_448_n11;
  tri   P1_sub_448_n14;
  tri   P1_sub_448_n255;
  tri   P1_sub_448_n254;
  tri   P1_sub_448_n253;
  tri   P1_sub_448_n4;
  tri   P1_sub_448_n7;
  tri   P1_sub_448_n252;
  tri   P1_sub_448_n251;
  tri   P1_sub_448_n250;
  tri   P1_sub_448_n249;
  tri   P1_sub_448_n248;
  tri   P1_sub_448_n247;
  tri   P1_sub_448_n246;
  tri   P1_sub_448_n245;
  tri   P1_sub_448_n244;
  tri   P1_sub_448_n243;
  tri   P1_sub_448_n242;
  tri   P1_sub_448_n241;
  tri   P1_sub_448_n240;
  tri   P1_sub_448_n239;
  tri   P1_sub_448_n238;
  tri   P1_sub_448_n237;
  tri   P1_sub_448_n236;
  tri   P1_sub_448_n235;
  tri   P1_sub_448_n234;
  tri   P1_sub_448_n233;
  tri   P1_sub_448_n232;
  tri   P1_sub_448_n231;
  tri   P1_sub_448_n230;
  tri   P1_sub_448_n229;
  tri   P1_sub_448_n228;
  tri   P1_sub_448_n227;
  tri   P1_sub_448_n226;
  tri   P1_sub_448_n225;
  tri   P1_sub_448_n224;
  tri   P1_sub_448_n223;
  tri   P1_sub_448_n222;
  tri   P1_sub_448_n221;
  tri   P1_sub_448_n220;
  tri   P1_sub_448_n219;
  tri   P1_sub_448_n218;
  tri   P1_sub_448_n217;
  tri   P1_sub_448_n203;
  tri   P1_sub_448_n209;
  tri   P1_sub_448_n216;
  tri   P1_sub_448_n215;
  tri   P1_sub_448_n210;
  tri   P1_sub_448_n214;
  tri   P1_sub_448_n211;
  tri   P1_sub_448_n213;
  tri   P1_sub_448_n212;
  tri   P1_sub_448_n277;
  tri   P1_sub_448_n281;
  tri   P1_sub_448_n280;
  tri   P1_sub_448_n152;
  tri   P1_add_468_n55;
  tri   P1_add_468_n54;
  tri   P1_add_468_n53;
  tri   P1_add_468_n51;
  tri   P1_add_468_n50;
  tri   P1_add_468_n48;
  tri   P1_add_468_n47;
  tri   P1_add_468_n46;
  tri   P1_add_468_n44;
  tri   P1_add_468_n43;
  tri   P1_add_468_n41;
  tri   P1_add_468_n40;
  tri   P1_add_468_n39;
  tri   P1_add_468_n37;
  tri   P1_add_468_n36;
  tri   P1_add_468_n34;
  tri   P1_add_468_n33;
  tri   P1_add_468_n32;
  tri   P1_add_468_n30;
  tri   P1_add_468_n29;
  tri   P1_add_468_n27;
  tri   P1_add_468_n26;
  tri   P1_add_468_n25;
  tri   P1_add_468_n23;
  tri   P1_add_468_n22;
  tri   P1_add_468_n20;
  tri   P1_add_468_n19;
  tri   P1_add_468_n18;
  tri   P1_add_468_n16;
  tri   P1_add_468_n15;
  tri   P1_add_468_n13;
  tri   P1_add_468_n12;
  tri   P1_add_468_n11;
  tri   P1_add_468_n9;
  tri   P1_add_468_n8;
  tri   P1_add_468_n6;
  tri   P1_add_468_n5;
  tri   P1_add_468_n4;
  tri   P1_add_468_n2;
  tri   P1_add_468_n1;
  tri   P1_add_468_n142;
  tri   P1_add_468_n140;
  tri   P1_add_468_n139;
  tri   P1_add_468_n138;
  tri   P1_add_468_n136;
  tri   P1_add_468_n135;
  tri   P1_add_468_n134;
  tri   P1_add_468_n132;
  tri   P1_add_468_n131;
  tri   P1_add_468_n130;
  tri   P1_add_468_n129;
  tri   P1_add_468_n128;
  tri   P1_add_468_n127;
  tri   P1_add_468_n126;
  tri   P1_add_468_n125;
  tri   P1_add_468_n124;
  tri   P1_add_468_n122;
  tri   P1_add_468_n121;
  tri   P1_add_468_n120;
  tri   P1_add_468_n119;
  tri   P1_add_468_n118;
  tri   P1_add_468_n117;
  tri   P1_add_468_n116;
  tri   P1_add_468_n115;
  tri   P1_add_468_n114;
  tri   P1_add_468_n112;
  tri   P1_add_468_n111;
  tri   P1_add_468_n110;
  tri   P1_add_468_n109;
  tri   P1_add_468_n108;
  tri   P1_add_468_n107;
  tri   P1_add_468_n106;
  tri   P1_add_468_n105;
  tri   P1_add_468_n104;
  tri   P1_add_468_n102;
  tri   P1_add_468_n101;
  tri   P1_add_468_n100;
  tri   P1_add_468_n99;
  tri   P1_add_468_n98;
  tri   P1_add_468_n97;
  tri   P1_add_468_n96;
  tri   P1_add_468_n95;
  tri   P1_add_468_n94;
  tri   P1_add_468_n92;
  tri   P1_add_468_n91;
  tri   P1_add_468_n90;
  tri   P1_add_468_n89;
  tri   P1_add_468_n88;
  tri   P1_add_468_n87;
  tri   P1_add_468_n86;
  tri   P1_add_468_n85;
  tri   P1_add_468_n84;
  tri   P1_add_468_n82;
  tri   P1_add_468_n81;
  tri   P1_add_468_n80;
  tri   P1_add_468_n79;
  tri   P1_add_468_n78;
  tri   P1_add_468_n77;
  tri   P1_add_468_n76;
  tri   P1_add_468_n75;
  tri   P1_add_468_n74;
  tri   P1_add_468_n72;
  tri   P1_add_468_n71;
  tri   P1_add_468_n70;
  tri   P1_add_468_n69;
  tri   P1_add_468_n68;
  tri   P1_add_468_n66;
  tri   P1_add_468_n65;
  tri   P1_add_468_n64;
  tri   P1_add_468_n63;
  tri   P1_add_468_n62;
  tri   P1_add_468_n61;
  tri   P1_add_468_n60;
  tri   P1_add_468_n59;
  tri   P1_add_468_n58;
  tri   P1_add_468_n57;
  tri   P1_add_468_n227;
  tri   P1_add_468_n226;
  tri   P1_add_468_n225;
  tri   P1_add_468_n223;
  tri   P1_add_468_n222;
  tri   P1_add_468_n221;
  tri   P1_add_468_n219;
  tri   P1_add_468_n218;
  tri   P1_add_468_n217;
  tri   P1_add_468_n216;
  tri   P1_add_468_n215;
  tri   P1_add_468_n214;
  tri   P1_add_468_n213;
  tri   P1_add_468_n212;
  tri   P1_add_468_n211;
  tri   P1_add_468_n209;
  tri   P1_add_468_n208;
  tri   P1_add_468_n207;
  tri   P1_add_468_n206;
  tri   P1_add_468_n205;
  tri   P1_add_468_n204;
  tri   P1_add_468_n203;
  tri   P1_add_468_n202;
  tri   P1_add_468_n201;
  tri   P1_add_468_n199;
  tri   P1_add_468_n198;
  tri   P1_add_468_n197;
  tri   P1_add_468_n196;
  tri   P1_add_468_n195;
  tri   P1_add_468_n194;
  tri   P1_add_468_n193;
  tri   P1_add_468_n192;
  tri   P1_add_468_n191;
  tri   P1_add_468_n189;
  tri   P1_add_468_n188;
  tri   P1_add_468_n187;
  tri   P1_add_468_n186;
  tri   P1_add_468_n185;
  tri   P1_add_468_n184;
  tri   P1_add_468_n183;
  tri   P1_add_468_n182;
  tri   P1_add_468_n181;
  tri   P1_add_468_n179;
  tri   P1_add_468_n178;
  tri   P1_add_468_n177;
  tri   P1_add_468_n176;
  tri   P1_add_468_n175;
  tri   P1_add_468_n174;
  tri   P1_add_468_n173;
  tri   P1_add_468_n172;
  tri   P1_add_468_n171;
  tri   P1_add_468_n169;
  tri   P1_add_468_n168;
  tri   P1_add_468_n167;
  tri   P1_add_468_n166;
  tri   P1_add_468_n165;
  tri   P1_add_468_n164;
  tri   P1_add_468_n163;
  tri   P1_add_468_n162;
  tri   P1_add_468_n161;
  tri   P1_add_468_n159;
  tri   P1_add_468_n158;
  tri   P1_add_468_n157;
  tri   P1_add_468_n156;
  tri   P1_add_468_n155;
  tri   P1_add_468_n153;
  tri   P1_add_468_n152;
  tri   P1_add_468_n150;
  tri   P1_add_468_n149;
  tri   P1_add_468_n148;
  tri   P1_add_468_n147;
  tri   P1_add_468_n146;
  tri   P1_add_468_n137;
  tri   P1_add_468_n145;
  tri   P1_add_468_n144;
  tri   P1_add_468_n141;
  tri   P1_add_468_n279;
  tri   P1_add_468_n278;
  tri   P1_add_468_n151;
  tri   P1_add_468_n277;
  tri   P1_add_468_n276;
  tri   P1_add_468_n275;
  tri   P1_add_468_n52;
  tri   P1_add_468_n274;
  tri   P1_add_468_n273;
  tri   P1_add_468_n272;
  tri   P1_add_468_n45;
  tri   P1_add_468_n271;
  tri   P1_add_468_n270;
  tri   P1_add_468_n269;
  tri   P1_add_468_n38;
  tri   P1_add_468_n268;
  tri   P1_add_468_n267;
  tri   P1_add_468_n266;
  tri   P1_add_468_n31;
  tri   P1_add_468_n265;
  tri   P1_add_468_n264;
  tri   P1_add_468_n263;
  tri   P1_add_468_n24;
  tri   P1_add_468_n262;
  tri   P1_add_468_n261;
  tri   P1_add_468_n260;
  tri   P1_add_468_n17;
  tri   P1_add_468_n259;
  tri   P1_add_468_n258;
  tri   P1_add_468_n257;
  tri   P1_add_468_n10;
  tri   P1_add_468_n256;
  tri   P1_add_468_n255;
  tri   P1_add_468_n254;
  tri   P1_add_468_n3;
  tri   P1_add_468_n253;
  tri   P1_add_468_n252;
  tri   P1_add_468_n251;
  tri   P1_add_468_n249;
  tri   P1_add_468_n248;
  tri   P1_add_468_n247;
  tri   P1_add_468_n246;
  tri   P1_add_468_n245;
  tri   P1_add_468_n244;
  tri   P1_add_468_n243;
  tri   P1_add_468_n242;
  tri   P1_add_468_n241;
  tri   P1_add_468_n239;
  tri   P1_add_468_n238;
  tri   P1_add_468_n237;
  tri   P1_add_468_n236;
  tri   P1_add_468_n235;
  tri   P1_add_468_n234;
  tri   P1_add_468_n233;
  tri   P1_add_468_n224;
  tri   P1_add_468_n232;
  tri   P1_add_468_n231;
  tri   P1_add_468_n228;
  tri   P1_add_468_n229;
  tri   r845_n27;
  tri   r845_n26;
  tri   r845_n25;
  tri   r845_n23;
  tri   r845_n22;
  tri   r845_n20;
  tri   r845_n19;
  tri   r845_n18;
  tri   r845_n16;
  tri   r845_n15;
  tri   r845_n13;
  tri   r845_n12;
  tri   r845_n11;
  tri   r845_n9;
  tri   r845_n8;
  tri   r845_n6;
  tri   r845_n5;
  tri   r845_n4;
  tri   r845_n2;
  tri   r845_n1;
  tri   r845_n115;
  tri   r845_n112;
  tri   r845_n111;
  tri   r845_n110;
  tri   r845_n109;
  tri   r845_n108;
  tri   r845_n107;
  tri   r845_n106;
  tri   r845_n105;
  tri   r845_n104;
  tri   r845_n102;
  tri   r845_n101;
  tri   r845_n100;
  tri   r845_n99;
  tri   r845_n98;
  tri   r845_n97;
  tri   r845_n96;
  tri   r845_n95;
  tri   r845_n94;
  tri   r845_n92;
  tri   r845_n91;
  tri   r845_n90;
  tri   r845_n89;
  tri   r845_n88;
  tri   r845_n87;
  tri   r845_n86;
  tri   r845_n85;
  tri   r845_n84;
  tri   r845_n82;
  tri   r845_n81;
  tri   r845_n80;
  tri   r845_n79;
  tri   r845_n78;
  tri   r845_n77;
  tri   r845_n76;
  tri   r845_n75;
  tri   r845_n74;
  tri   r845_n72;
  tri   r845_n71;
  tri   r845_n70;
  tri   r845_n69;
  tri   r845_n68;
  tri   r845_n66;
  tri   r845_n65;
  tri   r845_n64;
  tri   r845_n63;
  tri   r845_n62;
  tri   r845_n61;
  tri   r845_n60;
  tri   r845_n59;
  tri   r845_n58;
  tri   r845_n57;
  tri   r845_n55;
  tri   r845_n54;
  tri   r845_n53;
  tri   r845_n51;
  tri   r845_n50;
  tri   r845_n48;
  tri   r845_n47;
  tri   r845_n46;
  tri   r845_n44;
  tri   r845_n43;
  tri   r845_n41;
  tri   r845_n40;
  tri   r845_n39;
  tri   r845_n37;
  tri   r845_n36;
  tri   r845_n34;
  tri   r845_n33;
  tri   r845_n32;
  tri   r845_n30;
  tri   r845_n29;
  tri   r845_n199;
  tri   r845_n198;
  tri   r845_n197;
  tri   r845_n196;
  tri   r845_n195;
  tri   r845_n194;
  tri   r845_n193;
  tri   r845_n192;
  tri   r845_n191;
  tri   r845_n189;
  tri   r845_n188;
  tri   r845_n187;
  tri   r845_n186;
  tri   r845_n185;
  tri   r845_n184;
  tri   r845_n183;
  tri   r845_n182;
  tri   r845_n181;
  tri   r845_n179;
  tri   r845_n178;
  tri   r845_n177;
  tri   r845_n176;
  tri   r845_n175;
  tri   r845_n174;
  tri   r845_n173;
  tri   r845_n172;
  tri   r845_n171;
  tri   r845_n169;
  tri   r845_n168;
  tri   r845_n167;
  tri   r845_n166;
  tri   r845_n165;
  tri   r845_n163;
  tri   r845_n162;
  tri   r845_n160;
  tri   r845_n159;
  tri   r845_n158;
  tri   r845_n157;
  tri   r845_n156;
  tri   r845_n155;
  tri   r845_n154;
  tri   r845_n152;
  tri   r845_n151;
  tri   r845_n150;
  tri   r845_n149;
  tri   r845_n148;
  tri   r845_n147;
  tri   r845_n146;
  tri   r845_n145;
  tri   r845_n144;
  tri   r845_n142;
  tri   r845_n141;
  tri   r845_n140;
  tri   r845_n139;
  tri   r845_n138;
  tri   r845_n137;
  tri   r845_n136;
  tri   r845_n135;
  tri   r845_n134;
  tri   r845_n132;
  tri   r845_n131;
  tri   r845_n130;
  tri   r845_n129;
  tri   r845_n128;
  tri   r845_n127;
  tri   r845_n126;
  tri   r845_n125;
  tri   r845_n124;
  tri   r845_n122;
  tri   r845_n121;
  tri   r845_n120;
  tri   r845_n119;
  tri   r845_n118;
  tri   r845_n114;
  tri   r845_n116;
  tri   r845_n117;
  tri   r845_n281;
  tri   r845_n280;
  tri   r845_n279;
  tri   r845_n38;
  tri   r845_n278;
  tri   r845_n277;
  tri   r845_n276;
  tri   r845_n31;
  tri   r845_n275;
  tri   r845_n274;
  tri   r845_n273;
  tri   r845_n24;
  tri   r845_n272;
  tri   r845_n271;
  tri   r845_n270;
  tri   r845_n17;
  tri   r845_n269;
  tri   r845_n268;
  tri   r845_n267;
  tri   r845_n10;
  tri   r845_n266;
  tri   r845_n265;
  tri   r845_n264;
  tri   r845_n3;
  tri   r845_n263;
  tri   r845_n262;
  tri   r845_n261;
  tri   r845_n259;
  tri   r845_n258;
  tri   r845_n257;
  tri   r845_n256;
  tri   r845_n255;
  tri   r845_n254;
  tri   r845_n253;
  tri   r845_n252;
  tri   r845_n251;
  tri   r845_n249;
  tri   r845_n248;
  tri   r845_n247;
  tri   r845_n246;
  tri   r845_n245;
  tri   r845_n244;
  tri   r845_n243;
  tri   r845_n242;
  tri   r845_n241;
  tri   r845_n239;
  tri   r845_n238;
  tri   r845_n237;
  tri   r845_n236;
  tri   r845_n235;
  tri   r845_n234;
  tri   r845_n233;
  tri   r845_n232;
  tri   r845_n231;
  tri   r845_n229;
  tri   r845_n228;
  tri   r845_n227;
  tri   r845_n226;
  tri   r845_n225;
  tri   r845_n224;
  tri   r845_n223;
  tri   r845_n222;
  tri   r845_n221;
  tri   r845_n219;
  tri   r845_n218;
  tri   r845_n217;
  tri   r845_n216;
  tri   r845_n215;
  tri   r845_n214;
  tri   r845_n213;
  tri   r845_n212;
  tri   r845_n211;
  tri   r845_n209;
  tri   r845_n208;
  tri   r845_n207;
  tri   r845_n206;
  tri   r845_n205;
  tri   r845_n201;
  tri   r845_n204;
  tri   r845_n202;
  tri   r845_n203;
  tri   r845_n289;
  tri   r845_n288;
  tri   r845_n161;
  tri   r845_n287;
  tri   r845_n286;
  tri   r845_n285;
  tri   r845_n52;
  tri   r845_n284;
  tri   r845_n45;
  tri   r845_n283;
  tri   r845_n282;
  tri   r847_n78;
  tri   r847_n77;
  tri   r847_n74;
  tri   r847_n73;
  tri   r847_n72;
  tri   r847_n71;
  tri   r847_n70;
  tri   r847_n69;
  tri   r847_n67;
  tri   r847_n66;
  tri   r847_n65;
  tri   r847_n63;
  tri   r847_n62;
  tri   r847_n61;
  tri   r847_n59;
  tri   r847_n60;
  tri   r847_n58;
  tri   r847_n57;
  tri   r847_n55;
  tri   r847_n54;
  tri   r847_n52;
  tri   r847_n51;
  tri   r847_n50;
  tri   r847_n48;
  tri   r847_n47;
  tri   r847_n45;
  tri   r847_n44;
  tri   r847_n43;
  tri   r847_n41;
  tri   r847_n40;
  tri   r847_n38;
  tri   r847_n37;
  tri   r847_n36;
  tri   r847_n34;
  tri   r847_n33;
  tri   r847_n31;
  tri   r847_n30;
  tri   r847_n29;
  tri   r847_n27;
  tri   r847_n26;
  tri   r847_n24;
  tri   r847_n23;
  tri   r847_n22;
  tri   r847_n20;
  tri   r847_n19;
  tri   r847_n17;
  tri   r847_n16;
  tri   r847_n15;
  tri   r847_n13;
  tri   r847_n12;
  tri   r847_n10;
  tri   r847_n9;
  tri   r847_n8;
  tri   r847_n6;
  tri   r847_n5;
  tri   r847_n3;
  tri   r847_n2;
  tri   r847_n1;
  tri   r847_n161;
  tri   r847_n160;
  tri   r847_n159;
  tri   r847_n158;
  tri   r847_n157;
  tri   r847_n154;
  tri   r847_n153;
  tri   r847_n152;
  tri   r847_n151;
  tri   r847_n150;
  tri   r847_n149;
  tri   r847_n148;
  tri   r847_n147;
  tri   r847_n146;
  tri   r847_n145;
  tri   r847_n144;
  tri   r847_n143;
  tri   r847_n142;
  tri   r847_n141;
  tri   r847_n140;
  tri   r847_n139;
  tri   r847_n138;
  tri   r847_n137;
  tri   r847_n136;
  tri   r847_n135;
  tri   r847_n134;
  tri   r847_n133;
  tri   r847_n132;
  tri   r847_n131;
  tri   r847_n130;
  tri   r847_n129;
  tri   r847_n128;
  tri   r847_n127;
  tri   r847_n126;
  tri   r847_n125;
  tri   r847_n124;
  tri   r847_n123;
  tri   r847_n122;
  tri   r847_n121;
  tri   r847_n120;
  tri   r847_n119;
  tri   r847_n118;
  tri   r847_n117;
  tri   r847_n116;
  tri   r847_n115;
  tri   r847_n114;
  tri   r847_n113;
  tri   r847_n112;
  tri   r847_n111;
  tri   r847_n110;
  tri   r847_n109;
  tri   r847_n108;
  tri   r847_n107;
  tri   r847_n106;
  tri   r847_n105;
  tri   r847_n104;
  tri   r847_n103;
  tri   r847_n102;
  tri   r847_n101;
  tri   r847_n100;
  tri   r847_n99;
  tri   r847_n98;
  tri   r847_n97;
  tri   r847_n96;
  tri   r847_n95;
  tri   r847_n94;
  tri   r847_n93;
  tri   r847_n92;
  tri   r847_n91;
  tri   r847_n90;
  tri   r847_n89;
  tri   r847_n75;
  tri   r847_n88;
  tri   r847_n87;
  tri   r847_n86;
  tri   r847_n85;
  tri   r847_n84;
  tri   r847_n83;
  tri   r847_n82;
  tri   r847_n81;
  tri   r847_n76;
  tri   r847_n80;
  tri   r847_n79;
  tri   r847_n64;
  tri   r847_n248;
  tri   r847_n247;
  tri   r847_n246;
  tri   r847_n245;
  tri   r847_n242;
  tri   r847_n241;
  tri   r847_n240;
  tri   r847_n239;
  tri   r847_n238;
  tri   r847_n237;
  tri   r847_n236;
  tri   r847_n235;
  tri   r847_n234;
  tri   r847_n233;
  tri   r847_n232;
  tri   r847_n231;
  tri   r847_n230;
  tri   r847_n229;
  tri   r847_n228;
  tri   r847_n227;
  tri   r847_n226;
  tri   r847_n225;
  tri   r847_n224;
  tri   r847_n223;
  tri   r847_n222;
  tri   r847_n221;
  tri   r847_n220;
  tri   r847_n219;
  tri   r847_n218;
  tri   r847_n217;
  tri   r847_n216;
  tri   r847_n215;
  tri   r847_n214;
  tri   r847_n213;
  tri   r847_n212;
  tri   r847_n211;
  tri   r847_n210;
  tri   r847_n209;
  tri   r847_n208;
  tri   r847_n207;
  tri   r847_n206;
  tri   r847_n205;
  tri   r847_n204;
  tri   r847_n203;
  tri   r847_n202;
  tri   r847_n201;
  tri   r847_n200;
  tri   r847_n199;
  tri   r847_n198;
  tri   r847_n197;
  tri   r847_n196;
  tri   r847_n195;
  tri   r847_n194;
  tri   r847_n193;
  tri   r847_n192;
  tri   r847_n191;
  tri   r847_n190;
  tri   r847_n189;
  tri   r847_n188;
  tri   r847_n187;
  tri   r847_n186;
  tri   r847_n185;
  tri   r847_n184;
  tri   r847_n183;
  tri   r847_n182;
  tri   r847_n181;
  tri   r847_n180;
  tri   r847_n179;
  tri   r847_n178;
  tri   r847_n177;
  tri   r847_n155;
  tri   r847_n176;
  tri   r847_n175;
  tri   r847_n174;
  tri   r847_n173;
  tri   r847_n172;
  tri   r847_n171;
  tri   r847_n170;
  tri   r847_n169;
  tri   r847_n156;
  tri   r847_n168;
  tri   r847_n167;
  tri   r847_n163;
  tri   r847_n164;
  tri   r847_n291;
  tri   r847_n290;
  tri   r847_n289;
  tri   r847_n288;
  tri   r847_n162;
  tri   r847_n287;
  tri   r847_n166;
  tri   r847_n286;
  tri   r847_n285;
  tri   r847_n284;
  tri   r847_n53;
  tri   r847_n56;
  tri   r847_n283;
  tri   r847_n282;
  tri   r847_n281;
  tri   r847_n46;
  tri   r847_n49;
  tri   r847_n280;
  tri   r847_n279;
  tri   r847_n278;
  tri   r847_n39;
  tri   r847_n42;
  tri   r847_n277;
  tri   r847_n276;
  tri   r847_n275;
  tri   r847_n32;
  tri   r847_n35;
  tri   r847_n274;
  tri   r847_n273;
  tri   r847_n272;
  tri   r847_n25;
  tri   r847_n28;
  tri   r847_n271;
  tri   r847_n270;
  tri   r847_n269;
  tri   r847_n18;
  tri   r847_n21;
  tri   r847_n268;
  tri   r847_n267;
  tri   r847_n266;
  tri   r847_n11;
  tri   r847_n14;
  tri   r847_n265;
  tri   r847_n264;
  tri   r847_n263;
  tri   r847_n4;
  tri   r847_n7;
  tri   r847_n262;
  tri   r847_n261;
  tri   r847_n260;
  tri   r847_n259;
  tri   r847_n258;
  tri   r847_n257;
  tri   r847_n243;
  tri   r847_n249;
  tri   r847_n256;
  tri   r847_n255;
  tri   r847_n254;
  tri   r847_n253;
  tri   r847_n252;
  tri   r847_n244;
  tri   r847_n251;
  tri   r847_n250;
  tri   r849_n16;
  tri   r849_n15;
  tri   r849_n13;
  tri   r849_n12;
  tri   r849_n11;
  tri   r849_n9;
  tri   r849_n8;
  tri   r849_n6;
  tri   r849_n5;
  tri   r849_n4;
  tri   r849_n2;
  tri   r849_n1;
  tri   r849_n106;
  tri   r849_n105;
  tri   r849_n102;
  tri   r849_n101;
  tri   r849_n100;
  tri   r849_n99;
  tri   r849_n98;
  tri   r849_n97;
  tri   r849_n96;
  tri   r849_n95;
  tri   r849_n94;
  tri   r849_n92;
  tri   r849_n91;
  tri   r849_n90;
  tri   r849_n89;
  tri   r849_n88;
  tri   r849_n87;
  tri   r849_n86;
  tri   r849_n85;
  tri   r849_n84;
  tri   r849_n82;
  tri   r849_n81;
  tri   r849_n80;
  tri   r849_n79;
  tri   r849_n78;
  tri   r849_n77;
  tri   r849_n76;
  tri   r849_n75;
  tri   r849_n74;
  tri   r849_n72;
  tri   r849_n71;
  tri   r849_n70;
  tri   r849_n69;
  tri   r849_n68;
  tri   r849_n66;
  tri   r849_n65;
  tri   r849_n64;
  tri   r849_n63;
  tri   r849_n62;
  tri   r849_n61;
  tri   r849_n60;
  tri   r849_n59;
  tri   r849_n58;
  tri   r849_n57;
  tri   r849_n55;
  tri   r849_n54;
  tri   r849_n53;
  tri   r849_n51;
  tri   r849_n50;
  tri   r849_n48;
  tri   r849_n47;
  tri   r849_n46;
  tri   r849_n44;
  tri   r849_n43;
  tri   r849_n41;
  tri   r849_n40;
  tri   r849_n39;
  tri   r849_n37;
  tri   r849_n36;
  tri   r849_n34;
  tri   r849_n33;
  tri   r849_n32;
  tri   r849_n30;
  tri   r849_n29;
  tri   r849_n27;
  tri   r849_n26;
  tri   r849_n25;
  tri   r849_n23;
  tri   r849_n22;
  tri   r849_n18;
  tri   r849_n20;
  tri   r849_n19;
  tri   r849_n192;
  tri   r849_n189;
  tri   r849_n188;
  tri   r849_n187;
  tri   r849_n186;
  tri   r849_n185;
  tri   r849_n184;
  tri   r849_n183;
  tri   r849_n182;
  tri   r849_n181;
  tri   r849_n179;
  tri   r849_n178;
  tri   r849_n177;
  tri   r849_n176;
  tri   r849_n175;
  tri   r849_n174;
  tri   r849_n173;
  tri   r849_n172;
  tri   r849_n171;
  tri   r849_n169;
  tri   r849_n168;
  tri   r849_n167;
  tri   r849_n166;
  tri   r849_n165;
  tri   r849_n163;
  tri   r849_n162;
  tri   r849_n160;
  tri   r849_n159;
  tri   r849_n158;
  tri   r849_n157;
  tri   r849_n156;
  tri   r849_n155;
  tri   r849_n154;
  tri   r849_n152;
  tri   r849_n151;
  tri   r849_n150;
  tri   r849_n149;
  tri   r849_n148;
  tri   r849_n147;
  tri   r849_n146;
  tri   r849_n145;
  tri   r849_n144;
  tri   r849_n142;
  tri   r849_n141;
  tri   r849_n140;
  tri   r849_n139;
  tri   r849_n138;
  tri   r849_n137;
  tri   r849_n136;
  tri   r849_n135;
  tri   r849_n134;
  tri   r849_n132;
  tri   r849_n131;
  tri   r849_n130;
  tri   r849_n129;
  tri   r849_n128;
  tri   r849_n127;
  tri   r849_n126;
  tri   r849_n125;
  tri   r849_n124;
  tri   r849_n122;
  tri   r849_n121;
  tri   r849_n120;
  tri   r849_n119;
  tri   r849_n118;
  tri   r849_n117;
  tri   r849_n116;
  tri   r849_n115;
  tri   r849_n114;
  tri   r849_n112;
  tri   r849_n111;
  tri   r849_n110;
  tri   r849_n109;
  tri   r849_n108;
  tri   r849_n104;
  tri   r849_n107;
  tri   r849_n274;
  tri   r849_n24;
  tri   r849_n272;
  tri   r849_n271;
  tri   r849_n270;
  tri   r849_n17;
  tri   r849_n269;
  tri   r849_n268;
  tri   r849_n267;
  tri   r849_n10;
  tri   r849_n266;
  tri   r849_n265;
  tri   r849_n264;
  tri   r849_n3;
  tri   r849_n263;
  tri   r849_n262;
  tri   r849_n261;
  tri   r849_n259;
  tri   r849_n258;
  tri   r849_n257;
  tri   r849_n256;
  tri   r849_n255;
  tri   r849_n254;
  tri   r849_n253;
  tri   r849_n252;
  tri   r849_n251;
  tri   r849_n249;
  tri   r849_n248;
  tri   r849_n247;
  tri   r849_n246;
  tri   r849_n245;
  tri   r849_n244;
  tri   r849_n243;
  tri   r849_n242;
  tri   r849_n241;
  tri   r849_n239;
  tri   r849_n238;
  tri   r849_n237;
  tri   r849_n236;
  tri   r849_n235;
  tri   r849_n234;
  tri   r849_n233;
  tri   r849_n232;
  tri   r849_n231;
  tri   r849_n229;
  tri   r849_n228;
  tri   r849_n227;
  tri   r849_n226;
  tri   r849_n225;
  tri   r849_n224;
  tri   r849_n223;
  tri   r849_n222;
  tri   r849_n221;
  tri   r849_n219;
  tri   r849_n218;
  tri   r849_n217;
  tri   r849_n216;
  tri   r849_n215;
  tri   r849_n214;
  tri   r849_n213;
  tri   r849_n212;
  tri   r849_n211;
  tri   r849_n209;
  tri   r849_n208;
  tri   r849_n207;
  tri   r849_n206;
  tri   r849_n205;
  tri   r849_n204;
  tri   r849_n203;
  tri   r849_n202;
  tri   r849_n201;
  tri   r849_n199;
  tri   r849_n198;
  tri   r849_n197;
  tri   r849_n196;
  tri   r849_n195;
  tri   r849_n191;
  tri   r849_n193;
  tri   r849_n194;
  tri   r849_n289;
  tri   r849_n288;
  tri   r849_n161;
  tri   r849_n287;
  tri   r849_n286;
  tri   r849_n285;
  tri   r849_n52;
  tri   r849_n284;
  tri   r849_n283;
  tri   r849_n282;
  tri   r849_n45;
  tri   r849_n281;
  tri   r849_n280;
  tri   r849_n279;
  tri   r849_n38;
  tri   r849_n278;
  tri   r849_n277;
  tri   r849_n276;
  tri   r849_n273;
  tri   r849_n275;
  tri   r849_n31;
  tri   r851_n67;
  tri   r851_n66;
  tri   r851_n63;
  tri   r851_n62;
  tri   r851_n61;
  tri   r851_n59;
  tri   r851_n60;
  tri   r851_n58;
  tri   r851_n57;
  tri   r851_n55;
  tri   r851_n54;
  tri   r851_n52;
  tri   r851_n51;
  tri   r851_n50;
  tri   r851_n48;
  tri   r851_n47;
  tri   r851_n45;
  tri   r851_n44;
  tri   r851_n43;
  tri   r851_n41;
  tri   r851_n40;
  tri   r851_n38;
  tri   r851_n37;
  tri   r851_n36;
  tri   r851_n34;
  tri   r851_n33;
  tri   r851_n31;
  tri   r851_n30;
  tri   r851_n29;
  tri   r851_n27;
  tri   r851_n26;
  tri   r851_n24;
  tri   r851_n23;
  tri   r851_n22;
  tri   r851_n20;
  tri   r851_n19;
  tri   r851_n17;
  tri   r851_n16;
  tri   r851_n15;
  tri   r851_n13;
  tri   r851_n12;
  tri   r851_n10;
  tri   r851_n9;
  tri   r851_n8;
  tri   r851_n6;
  tri   r851_n5;
  tri   r851_n3;
  tri   r851_n2;
  tri   r851_n1;
  tri   r851_n153;
  tri   r851_n150;
  tri   r851_n149;
  tri   r851_n148;
  tri   r851_n147;
  tri   r851_n146;
  tri   r851_n144;
  tri   r851_n143;
  tri   r851_n142;
  tri   r851_n141;
  tri   r851_n140;
  tri   r851_n139;
  tri   r851_n138;
  tri   r851_n137;
  tri   r851_n136;
  tri   r851_n135;
  tri   r851_n134;
  tri   r851_n133;
  tri   r851_n132;
  tri   r851_n131;
  tri   r851_n130;
  tri   r851_n129;
  tri   r851_n128;
  tri   r851_n127;
  tri   r851_n126;
  tri   r851_n125;
  tri   r851_n124;
  tri   r851_n123;
  tri   r851_n122;
  tri   r851_n121;
  tri   r851_n120;
  tri   r851_n119;
  tri   r851_n118;
  tri   r851_n117;
  tri   r851_n116;
  tri   r851_n115;
  tri   r851_n114;
  tri   r851_n113;
  tri   r851_n112;
  tri   r851_n111;
  tri   r851_n110;
  tri   r851_n109;
  tri   r851_n108;
  tri   r851_n107;
  tri   r851_n106;
  tri   r851_n105;
  tri   r851_n104;
  tri   r851_n103;
  tri   r851_n102;
  tri   r851_n101;
  tri   r851_n100;
  tri   r851_n99;
  tri   r851_n98;
  tri   r851_n97;
  tri   r851_n96;
  tri   r851_n95;
  tri   r851_n94;
  tri   r851_n93;
  tri   r851_n92;
  tri   r851_n91;
  tri   r851_n90;
  tri   r851_n89;
  tri   r851_n88;
  tri   r851_n87;
  tri   r851_n86;
  tri   r851_n85;
  tri   r851_n84;
  tri   r851_n83;
  tri   r851_n82;
  tri   r851_n81;
  tri   r851_n80;
  tri   r851_n79;
  tri   r851_n64;
  tri   r851_n78;
  tri   r851_n77;
  tri   r851_n76;
  tri   r851_n75;
  tri   r851_n74;
  tri   r851_n73;
  tri   r851_n72;
  tri   r851_n71;
  tri   r851_n65;
  tri   r851_n70;
  tri   r851_n69;
  tri   r851_n238;
  tri   r851_n237;
  tri   r851_n236;
  tri   r851_n235;
  tri   r851_n234;
  tri   r851_n232;
  tri   r851_n231;
  tri   r851_n230;
  tri   r851_n229;
  tri   r851_n228;
  tri   r851_n227;
  tri   r851_n226;
  tri   r851_n225;
  tri   r851_n224;
  tri   r851_n223;
  tri   r851_n222;
  tri   r851_n221;
  tri   r851_n220;
  tri   r851_n219;
  tri   r851_n218;
  tri   r851_n217;
  tri   r851_n216;
  tri   r851_n215;
  tri   r851_n214;
  tri   r851_n213;
  tri   r851_n212;
  tri   r851_n211;
  tri   r851_n210;
  tri   r851_n209;
  tri   r851_n208;
  tri   r851_n207;
  tri   r851_n206;
  tri   r851_n205;
  tri   r851_n204;
  tri   r851_n203;
  tri   r851_n202;
  tri   r851_n201;
  tri   r851_n200;
  tri   r851_n199;
  tri   r851_n198;
  tri   r851_n197;
  tri   r851_n196;
  tri   r851_n195;
  tri   r851_n194;
  tri   r851_n193;
  tri   r851_n192;
  tri   r851_n191;
  tri   r851_n190;
  tri   r851_n189;
  tri   r851_n188;
  tri   r851_n187;
  tri   r851_n186;
  tri   r851_n185;
  tri   r851_n184;
  tri   r851_n183;
  tri   r851_n182;
  tri   r851_n181;
  tri   r851_n180;
  tri   r851_n179;
  tri   r851_n178;
  tri   r851_n177;
  tri   r851_n155;
  tri   r851_n176;
  tri   r851_n175;
  tri   r851_n174;
  tri   r851_n173;
  tri   r851_n172;
  tri   r851_n171;
  tri   r851_n170;
  tri   r851_n169;
  tri   r851_n168;
  tri   r851_n167;
  tri   r851_n164;
  tri   r851_n163;
  tri   r851_n161;
  tri   r851_n160;
  tri   r851_n159;
  tri   r851_n145;
  tri   r851_n151;
  tri   r851_n158;
  tri   r851_n157;
  tri   r851_n152;
  tri   r851_n154;
  tri   r851_n156;
  tri   r851_n291;
  tri   r851_n290;
  tri   r851_n289;
  tri   r851_n288;
  tri   r851_n162;
  tri   r851_n287;
  tri   r851_n166;
  tri   r851_n286;
  tri   r851_n285;
  tri   r851_n284;
  tri   r851_n53;
  tri   r851_n56;
  tri   r851_n283;
  tri   r851_n282;
  tri   r851_n281;
  tri   r851_n46;
  tri   r851_n49;
  tri   r851_n280;
  tri   r851_n279;
  tri   r851_n278;
  tri   r851_n39;
  tri   r851_n42;
  tri   r851_n277;
  tri   r851_n276;
  tri   r851_n275;
  tri   r851_n32;
  tri   r851_n35;
  tri   r851_n274;
  tri   r851_n273;
  tri   r851_n272;
  tri   r851_n25;
  tri   r851_n28;
  tri   r851_n271;
  tri   r851_n270;
  tri   r851_n269;
  tri   r851_n18;
  tri   r851_n21;
  tri   r851_n268;
  tri   r851_n267;
  tri   r851_n266;
  tri   r851_n11;
  tri   r851_n14;
  tri   r851_n265;
  tri   r851_n264;
  tri   r851_n263;
  tri   r851_n4;
  tri   r851_n7;
  tri   r851_n262;
  tri   r851_n261;
  tri   r851_n260;
  tri   r851_n259;
  tri   r851_n258;
  tri   r851_n257;
  tri   r851_n256;
  tri   r851_n255;
  tri   r851_n254;
  tri   r851_n253;
  tri   r851_n252;
  tri   r851_n251;
  tri   r851_n250;
  tri   r851_n249;
  tri   r851_n248;
  tri   r851_n247;
  tri   r851_n233;
  tri   r851_n239;
  tri   r851_n246;
  tri   r851_n245;
  tri   r851_n240;
  tri   r851_n244;
  tri   r851_n241;
  tri   r851_n243;
  tri   r851_n242;
  tri   r854_n6;
  tri   r854_n5;
  tri   r854_n4;
  tri   r854_n2;
  tri   r854_n1;
  tri   r854_n96;
  tri   r854_n95;
  tri   r854_n94;
  tri   r854_n92;
  tri   r854_n91;
  tri   r854_n90;
  tri   r854_n89;
  tri   r854_n88;
  tri   r854_n87;
  tri   r854_n86;
  tri   r854_n85;
  tri   r854_n84;
  tri   r854_n82;
  tri   r854_n81;
  tri   r854_n80;
  tri   r854_n79;
  tri   r854_n78;
  tri   r854_n77;
  tri   r854_n76;
  tri   r854_n75;
  tri   r854_n74;
  tri   r854_n72;
  tri   r854_n71;
  tri   r854_n70;
  tri   r854_n69;
  tri   r854_n68;
  tri   r854_n66;
  tri   r854_n65;
  tri   r854_n64;
  tri   r854_n63;
  tri   r854_n62;
  tri   r854_n61;
  tri   r854_n60;
  tri   r854_n59;
  tri   r854_n58;
  tri   r854_n57;
  tri   r854_n55;
  tri   r854_n54;
  tri   r854_n53;
  tri   r854_n51;
  tri   r854_n50;
  tri   r854_n48;
  tri   r854_n47;
  tri   r854_n46;
  tri   r854_n44;
  tri   r854_n43;
  tri   r854_n41;
  tri   r854_n40;
  tri   r854_n39;
  tri   r854_n37;
  tri   r854_n36;
  tri   r854_n34;
  tri   r854_n33;
  tri   r854_n32;
  tri   r854_n30;
  tri   r854_n29;
  tri   r854_n27;
  tri   r854_n26;
  tri   r854_n25;
  tri   r854_n23;
  tri   r854_n22;
  tri   r854_n20;
  tri   r854_n19;
  tri   r854_n18;
  tri   r854_n16;
  tri   r854_n15;
  tri   r854_n13;
  tri   r854_n12;
  tri   r854_n11;
  tri   r854_n9;
  tri   r854_n8;
  tri   r854_n183;
  tri   r854_n182;
  tri   r854_n179;
  tri   r854_n178;
  tri   r854_n177;
  tri   r854_n176;
  tri   r854_n175;
  tri   r854_n174;
  tri   r854_n173;
  tri   r854_n172;
  tri   r854_n171;
  tri   r854_n169;
  tri   r854_n168;
  tri   r854_n167;
  tri   r854_n166;
  tri   r854_n165;
  tri   r854_n163;
  tri   r854_n162;
  tri   r854_n160;
  tri   r854_n159;
  tri   r854_n158;
  tri   r854_n157;
  tri   r854_n156;
  tri   r854_n155;
  tri   r854_n154;
  tri   r854_n152;
  tri   r854_n151;
  tri   r854_n150;
  tri   r854_n149;
  tri   r854_n148;
  tri   r854_n147;
  tri   r854_n146;
  tri   r854_n145;
  tri   r854_n144;
  tri   r854_n142;
  tri   r854_n141;
  tri   r854_n140;
  tri   r854_n139;
  tri   r854_n138;
  tri   r854_n137;
  tri   r854_n136;
  tri   r854_n135;
  tri   r854_n134;
  tri   r854_n132;
  tri   r854_n131;
  tri   r854_n130;
  tri   r854_n129;
  tri   r854_n128;
  tri   r854_n127;
  tri   r854_n126;
  tri   r854_n125;
  tri   r854_n124;
  tri   r854_n122;
  tri   r854_n121;
  tri   r854_n120;
  tri   r854_n119;
  tri   r854_n118;
  tri   r854_n117;
  tri   r854_n116;
  tri   r854_n115;
  tri   r854_n114;
  tri   r854_n112;
  tri   r854_n111;
  tri   r854_n110;
  tri   r854_n109;
  tri   r854_n108;
  tri   r854_n107;
  tri   r854_n106;
  tri   r854_n105;
  tri   r854_n104;
  tri   r854_n102;
  tri   r854_n101;
  tri   r854_n100;
  tri   r854_n97;
  tri   r854_n99;
  tri   r854_n98;
  tri   r854_n266;
  tri   r854_n265;
  tri   r854_n264;
  tri   r854_n3;
  tri   r854_n263;
  tri   r854_n262;
  tri   r854_n261;
  tri   r854_n259;
  tri   r854_n258;
  tri   r854_n257;
  tri   r854_n256;
  tri   r854_n255;
  tri   r854_n254;
  tri   r854_n253;
  tri   r854_n252;
  tri   r854_n251;
  tri   r854_n249;
  tri   r854_n248;
  tri   r854_n247;
  tri   r854_n246;
  tri   r854_n245;
  tri   r854_n244;
  tri   r854_n243;
  tri   r854_n242;
  tri   r854_n241;
  tri   r854_n239;
  tri   r854_n238;
  tri   r854_n237;
  tri   r854_n236;
  tri   r854_n235;
  tri   r854_n234;
  tri   r854_n233;
  tri   r854_n232;
  tri   r854_n231;
  tri   r854_n229;
  tri   r854_n228;
  tri   r854_n227;
  tri   r854_n226;
  tri   r854_n225;
  tri   r854_n224;
  tri   r854_n223;
  tri   r854_n222;
  tri   r854_n221;
  tri   r854_n219;
  tri   r854_n218;
  tri   r854_n217;
  tri   r854_n216;
  tri   r854_n215;
  tri   r854_n214;
  tri   r854_n213;
  tri   r854_n212;
  tri   r854_n211;
  tri   r854_n209;
  tri   r854_n208;
  tri   r854_n207;
  tri   r854_n206;
  tri   r854_n205;
  tri   r854_n204;
  tri   r854_n203;
  tri   r854_n202;
  tri   r854_n201;
  tri   r854_n199;
  tri   r854_n198;
  tri   r854_n197;
  tri   r854_n196;
  tri   r854_n195;
  tri   r854_n194;
  tri   r854_n193;
  tri   r854_n192;
  tri   r854_n191;
  tri   r854_n189;
  tri   r854_n188;
  tri   r854_n187;
  tri   r854_n186;
  tri   r854_n185;
  tri   r854_n181;
  tri   r854_n184;
  tri   r854_n289;
  tri   r854_n288;
  tri   r854_n161;
  tri   r854_n287;
  tri   r854_n286;
  tri   r854_n285;
  tri   r854_n52;
  tri   r854_n284;
  tri   r854_n283;
  tri   r854_n282;
  tri   r854_n45;
  tri   r854_n281;
  tri   r854_n280;
  tri   r854_n279;
  tri   r854_n38;
  tri   r854_n278;
  tri   r854_n277;
  tri   r854_n276;
  tri   r854_n31;
  tri   r854_n275;
  tri   r854_n274;
  tri   r854_n273;
  tri   r854_n24;
  tri   r854_n272;
  tri   r854_n271;
  tri   r854_n270;
  tri   r854_n17;
  tri   r854_n269;
  tri   r854_n10;
  tri   r854_n268;
  tri   r854_n267;
  tri   r855_n62;
  tri   r855_n61;
  tri   r855_n60;
  tri   r855_n57;
  tri   r855_n56;
  tri   r855_n55;
  tri   r855_n54;
  tri   r855_n53;
  tri   r855_n52;
  tri   r855_n50;
  tri   r855_n49;
  tri   r855_n48;
  tri   r855_n47;
  tri   r855_n46;
  tri   r855_n45;
  tri   r855_n44;
  tri   r855_n42;
  tri   r855_n41;
  tri   r855_n40;
  tri   r855_n39;
  tri   r855_n38;
  tri   r855_n37;
  tri   r855_n36;
  tri   r855_n35;
  tri   r855_n34;
  tri   r855_n32;
  tri   r855_n31;
  tri   r855_n29;
  tri   r855_n28;
  tri   r855_n27;
  tri   r855_n24;
  tri   r855_n23;
  tri   r855_n22;
  tri   r855_n21;
  tri   r855_n20;
  tri   r855_n17;
  tri   r855_n16;
  tri   r855_n15;
  tri   r855_n14;
  tri   r855_n13;
  tri   r855_n10;
  tri   r855_n9;
  tri   r855_n8;
  tri   r855_n7;
  tri   r855_n6;
  tri   r855_n3;
  tri   r855_n2;
  tri   r855_n1;
  tri   r855_n124;
  tri   r855_n123;
  tri   r855_n121;
  tri   r855_n120;
  tri   r855_n26;
  tri   r855_n119;
  tri   r855_n19;
  tri   r855_n118;
  tri   r855_n12;
  tri   r855_n117;
  tri   r855_n5;
  tri   r855_n116;
  tri   r855_n115;
  tri   r855_n114;
  tri   r855_n113;
  tri   r855_n112;
  tri   r855_n111;
  tri   r855_n109;
  tri   r855_n108;
  tri   r855_n107;
  tri   r855_n106;
  tri   r855_n105;
  tri   r855_n104;
  tri   r855_n103;
  tri   r855_n101;
  tri   r855_n100;
  tri   r855_n99;
  tri   r855_n98;
  tri   r855_n97;
  tri   r855_n96;
  tri   r855_n95;
  tri   r855_n93;
  tri   r855_n92;
  tri   r855_n91;
  tri   r855_n90;
  tri   r855_n89;
  tri   r855_n88;
  tri   r855_n87;
  tri   r855_n85;
  tri   r855_n84;
  tri   r855_n83;
  tri   r855_n82;
  tri   r855_n81;
  tri   r855_n80;
  tri   r855_n79;
  tri   r855_n78;
  tri   r855_n77;
  tri   r855_n76;
  tri   r855_n74;
  tri   r855_n73;
  tri   r855_n72;
  tri   r855_n71;
  tri   r855_n70;
  tri   r855_n69;
  tri   r855_n68;
  tri   r855_n66;
  tri   r855_n65;
  tri   r855_n58;
  tri   r855_n64;
  tri   r855_n63;
  tri   r855_n11;
  tri   r855_n30;
  tri   r855_n51;
  tri   r855_n125;
  tri   r855_n128;
  tri   r855_n131;
  tri   r855_n134;
  tri   r855_n146;
  tri   r860_n107;
  tri   r860_n103;
  tri   r860_n102;
  tri   r860_n101;
  tri   r860_n100;
  tri   r860_n97;
  tri   r860_n96;
  tri   r860_n93;
  tri   r860_n92;
  tri   r860_n88;
  tri   r860_n87;
  tri   r860_n86;
  tri   r860_n85;
  tri   r860_n82;
  tri   r860_n81;
  tri   r860_n78;
  tri   r860_n77;
  tri   r860_n73;
  tri   r860_n72;
  tri   r860_n71;
  tri   r860_n70;
  tri   r860_n67;
  tri   r860_n66;
  tri   r860_n63;
  tri   r860_n62;
  tri   r860_n58;
  tri   r860_n57;
  tri   r860_n56;
  tri   r860_n55;
  tri   r860_n52;
  tri   r860_n51;
  tri   r860_n48;
  tri   r860_n47;
  tri   r860_n43;
  tri   r860_n42;
  tri   r860_n41;
  tri   r860_n40;
  tri   r860_n37;
  tri   r860_n36;
  tri   r860_n33;
  tri   r860_n32;
  tri   r860_n28;
  tri   r860_n27;
  tri   r860_n26;
  tri   r860_n25;
  tri   r860_n22;
  tri   r860_n21;
  tri   r860_n18;
  tri   r860_n17;
  tri   r860_n13;
  tri   r860_n12;
  tri   r860_n11;
  tri   r860_n10;
  tri   r860_n7;
  tri   r860_n5;
  tri   r860_n3;
  tri   r860_n2;
  tri   r860_n68;
  tri   r860_n198;
  tri   r860_n197;
  tri   r860_n195;
  tri   r860_n59;
  tri   r860_n61;
  tri   r860_n193;
  tri   r860_n192;
  tri   r860_n191;
  tri   r860_n190;
  tri   r860_n189;
  tri   r860_n188;
  tri   r860_n186;
  tri   r860_n53;
  tri   r860_n185;
  tri   r860_n184;
  tri   r860_n183;
  tri   r860_n182;
  tri   r860_n180;
  tri   r860_n44;
  tri   r860_n46;
  tri   r860_n178;
  tri   r860_n177;
  tri   r860_n176;
  tri   r860_n175;
  tri   r860_n174;
  tri   r860_n173;
  tri   r860_n171;
  tri   r860_n38;
  tri   r860_n170;
  tri   r860_n169;
  tri   r860_n168;
  tri   r860_n167;
  tri   r860_n165;
  tri   r860_n29;
  tri   r860_n31;
  tri   r860_n163;
  tri   r860_n162;
  tri   r860_n161;
  tri   r860_n160;
  tri   r860_n159;
  tri   r860_n158;
  tri   r860_n156;
  tri   r860_n23;
  tri   r860_n155;
  tri   r860_n154;
  tri   r860_n153;
  tri   r860_n152;
  tri   r860_n150;
  tri   r860_n14;
  tri   r860_n16;
  tri   r860_n148;
  tri   r860_n147;
  tri   r860_n146;
  tri   r860_n145;
  tri   r860_n144;
  tri   r860_n143;
  tri   r860_n6;
  tri   r860_n8;
  tri   r860_n140;
  tri   r860_n139;
  tri   r860_n138;
  tri   r860_n1;
  tri   r860_n136;
  tri   r860_n135;
  tri   r860_n133;
  tri   r860_n20;
  tri   r860_n131;
  tri   r860_n35;
  tri   r860_n129;
  tri   r860_n50;
  tri   r860_n65;
  tri   r860_n80;
  tri   r860_n95;
  tri   r860_n119;
  tri   r860_n118;
  tri   r860_n117;
  tri   r860_n115;
  tri   r860_n114;
  tri   r860_n112;
  tri   r860_n108;
  tri   r860_n111;
  tri   r860_n110;
  tri   r860_n60;
  tri   r860_n54;
  tri   r860_n128;
  tri   r860_n64;
  tri   r860_n196;
  tri   r860_n79;
  tri   r860_n94;
  tri   r860_n109;
  tri   r860_n120;
  tri   r860_n251;
  tri   r860_n250;
  tri   r860_n249;
  tri   r860_n248;
  tri   r860_n246;
  tri   r860_n121;
  tri   r860_n113;
  tri   r860_n245;
  tri   r860_n244;
  tri   r860_n243;
  tri   r860_n242;
  tri   r860_n241;
  tri   r860_n240;
  tri   r860_n122;
  tri   r860_n104;
  tri   r860_n106;
  tri   r860_n238;
  tri   r860_n237;
  tri   r860_n236;
  tri   r860_n235;
  tri   r860_n234;
  tri   r860_n99;
  tri   r860_n233;
  tri   r860_n105;
  tri   r860_n231;
  tri   r860_n123;
  tri   r860_n98;
  tri   r860_n230;
  tri   r860_n229;
  tri   r860_n228;
  tri   r860_n227;
  tri   r860_n226;
  tri   r860_n225;
  tri   r860_n124;
  tri   r860_n89;
  tri   r860_n91;
  tri   r860_n223;
  tri   r860_n222;
  tri   r860_n221;
  tri   r860_n220;
  tri   r860_n219;
  tri   r860_n84;
  tri   r860_n218;
  tri   r860_n90;
  tri   r860_n216;
  tri   r860_n125;
  tri   r860_n83;
  tri   r860_n215;
  tri   r860_n214;
  tri   r860_n213;
  tri   r860_n212;
  tri   r860_n211;
  tri   r860_n210;
  tri   r860_n126;
  tri   r860_n74;
  tri   r860_n76;
  tri   r860_n208;
  tri   r860_n207;
  tri   r860_n206;
  tri   r860_n205;
  tri   r860_n204;
  tri   r860_n69;
  tri   r860_n203;
  tri   r860_n75;
  tri   r860_n200;
  tri   r860_n127;
  tri   r860_n199;
  tri   r860_n201;
  tri   r860_n4;
  tri   r860_n15;
  tri   r860_n9;
  tri   r860_n134;
  tri   r860_n19;
  tri   r860_n151;
  tri   r860_n30;
  tri   r860_n24;
  tri   r860_n132;
  tri   r860_n34;
  tri   r860_n166;
  tri   r860_n45;
  tri   r860_n39;
  tri   r860_n130;
  tri   r860_n49;
  tri   r860_n181;
  tri   r860_n297;
  tri   r860_n300;
  tri   r860_n303;
  tri   r860_n309;
  tri   add_1095_n189;
  tri   add_1095_n188;
  tri   add_1095_n190;
  tri   add_1095_n183;
  tri   add_1095_n184;
  tri   add_1095_n182;
  tri   add_1095_n185;
  tri   add_1095_n186;
  tri   add_1095_n187;
  tri   add_1095_n177;
  tri   add_1095_n178;
  tri   add_1095_n176;
  tri   add_1095_n179;
  tri   add_1095_n180;
  tri   add_1095_n181;
  tri   add_1095_n171;
  tri   add_1095_n172;
  tri   add_1095_n170;
  tri   add_1095_n173;
  tri   add_1095_n174;
  tri   add_1095_n175;
  tri   add_1095_n165;
  tri   add_1095_n166;
  tri   add_1095_n164;
  tri   add_1095_n167;
  tri   add_1095_n168;
  tri   add_1095_n169;
  tri   add_1095_n157;
  tri   add_1095_n159;
  tri   add_1095_n158;
  tri   add_1095_n160;
  tri   add_1095_n161;
  tri   add_1095_n162;
  tri   add_1095_n163;
  tri   add_1095_n150;
  tri   add_1095_n152;
  tri   add_1095_n153;
  tri   add_1095_n151;
  tri   add_1095_n154;
  tri   add_1095_n156;
  tri   add_1095_n155;
  tri   add_1095_n142;
  tri   add_1095_n143;
  tri   add_1095_n141;
  tri   add_1095_n146;
  tri   add_1095_n144;
  tri   add_1095_n145;
  tri   add_1095_n147;
  tri   add_1095_n149;
  tri   add_1095_n148;
  tri   add_1095_n136;
  tri   add_1095_n135;
  tri   add_1095_n137;
  tri   add_1095_n139;
  tri   add_1095_n138;
  tri   add_1095_n140;
  tri   add_1095_n129;
  tri   add_1095_n128;
  tri   add_1095_n130;
  tri   add_1095_n131;
  tri   add_1095_n132;
  tri   add_1095_n133;
  tri   add_1095_n134;
  tri   add_1095_n122;
  tri   add_1095_n123;
  tri   add_1095_n121;
  tri   add_1095_n125;
  tri   add_1095_n126;
  tri   add_1095_n127;
  tri   add_1095_n124;
  tri   add_1095_n113;
  tri   add_1095_n116;
  tri   add_1095_n114;
  tri   add_1095_n115;
  tri   add_1095_n117;
  tri   add_1095_n118;
  tri   add_1095_n119;
  tri   add_1095_n120;
  tri   add_1095_n106;
  tri   add_1095_n105;
  tri   add_1095_n107;
  tri   add_1095_n109;
  tri   add_1095_n108;
  tri   add_1095_n110;
  tri   add_1095_n112;
  tri   add_1095_n111;
  tri   add_1095_n99;
  tri   add_1095_n98;
  tri   add_1095_n100;
  tri   add_1095_n102;
  tri   add_1095_n103;
  tri   add_1095_n101;
  tri   add_1095_n104;
  tri   add_1095_n92;
  tri   add_1095_n93;
  tri   add_1095_n91;
  tri   add_1095_n96;
  tri   add_1095_n97;
  tri   add_1095_n94;
  tri   add_1095_n95;
  tri   add_1095_n86;
  tri   add_1095_n84;
  tri   add_1095_n85;
  tri   add_1095_n87;
  tri   add_1095_n89;
  tri   add_1095_n88;
  tri   add_1095_n90;
  tri   add_1095_n77;
  tri   add_1095_n79;
  tri   add_1095_n78;
  tri   add_1095_n80;
  tri   add_1095_n81;
  tri   add_1095_n82;
  tri   add_1095_n83;
  tri   add_1095_n70;
  tri   add_1095_n71;
  tri   add_1095_n73;
  tri   add_1095_n72;
  tri   add_1095_n74;
  tri   add_1095_n76;
  tri   add_1095_n75;
  tri   add_1095_n62;
  tri   add_1095_n61;
  tri   add_1095_n63;
  tri   add_1095_n65;
  tri   add_1095_n67;
  tri   add_1095_n64;
  tri   add_1095_n66;
  tri   add_1095_n69;
  tri   add_1095_n68;
  tri   add_1095_n52;
  tri   add_1095_n53;
  tri   add_1095_n55;
  tri   add_1095_n54;
  tri   add_1095_n56;
  tri   add_1095_n57;
  tri   add_1095_n58;
  tri   add_1095_n59;
  tri   add_1095_n60;
  tri   add_1095_n44;
  tri   add_1095_n45;
  tri   add_1095_n43;
  tri   add_1095_n46;
  tri   add_1095_n48;
  tri   add_1095_n47;
  tri   add_1095_n49;
  tri   add_1095_n51;
  tri   add_1095_n50;
  tri   add_1095_n37;
  tri   add_1095_n38;
  tri   add_1095_n36;
  tri   add_1095_n39;
  tri   add_1095_n41;
  tri   add_1095_n40;
  tri   add_1095_n42;
  tri   add_1095_n30;
  tri   add_1095_n31;
  tri   add_1095_n29;
  tri   add_1095_n32;
  tri   add_1095_n34;
  tri   add_1095_n33;
  tri   add_1095_n35;
  tri   add_1095_n21;
  tri   add_1095_n23;
  tri   add_1095_n24;
  tri   add_1095_n22;
  tri   add_1095_n25;
  tri   add_1095_n26;
  tri   add_1095_n27;
  tri   add_1095_n28;
  tri   add_1095_n13;
  tri   add_1095_n12;
  tri   add_1095_n14;
  tri   add_1095_n16;
  tri   add_1095_n17;
  tri   add_1095_n15;
  tri   add_1095_n18;
  tri   add_1095_n20;
  tri   add_1095_n19;
  tri   add_1095_n6;
  tri   add_1095_n5;
  tri   add_1095_n7;
  tri   add_1095_n9;
  tri   add_1095_n11;
  tri   add_1095_n10;
  tri   add_1095_n8;
  tri   add_1095_n1;
  tri   add_1095_n2;
  tri   add_1095_n4;
  tri   add_1095_n3;
  tri   P2_sub_621_n33;
  tri   P2_sub_621_n32;
  tri   P2_sub_621_n31;
  tri   P2_sub_621_n29;
  tri   P2_sub_621_n28;
  tri   P2_sub_621_n27;
  tri   P2_sub_621_n26;
  tri   P2_sub_621_n25;
  tri   P2_sub_621_n24;
  tri   P2_sub_621_n23;
  tri   P2_sub_621_n22;
  tri   P2_sub_621_n20;
  tri   P2_sub_621_n19;
  tri   P2_sub_621_n18;
  tri   P2_sub_621_n16;
  tri   P2_sub_621_n15;
  tri   P2_sub_621_n14;
  tri   P2_sub_621_n13;
  tri   P2_sub_621_n12;
  tri   P2_sub_621_n11;
  tri   P2_sub_621_n10;
  tri   P2_sub_621_n9;
  tri   P2_sub_621_n7;
  tri   P2_sub_621_n6;
  tri   P2_sub_621_n5;
  tri   P2_sub_621_n3;
  tri   P2_sub_621_n2;
  tri   P2_sub_621_n107;
  tri   P2_sub_621_n106;
  tri   P2_sub_621_n105;
  tri   P2_sub_621_n104;
  tri   P2_sub_621_n103;
  tri   P2_sub_621_n102;
  tri   P2_sub_621_n101;
  tri   P2_sub_621_n100;
  tri   P2_sub_621_n99;
  tri   P2_sub_621_n98;
  tri   P2_sub_621_n97;
  tri   P2_sub_621_n96;
  tri   P2_sub_621_n95;
  tri   P2_sub_621_n94;
  tri   P2_sub_621_n93;
  tri   P2_sub_621_n92;
  tri   P2_sub_621_n91;
  tri   P2_sub_621_n90;
  tri   P2_sub_621_n89;
  tri   P2_sub_621_n88;
  tri   P2_sub_621_n87;
  tri   P2_sub_621_n86;
  tri   P2_sub_621_n85;
  tri   P2_sub_621_n84;
  tri   P2_sub_621_n83;
  tri   P2_sub_621_n82;
  tri   P2_sub_621_n81;
  tri   P2_sub_621_n80;
  tri   P2_sub_621_n79;
  tri   P2_sub_621_n78;
  tri   P2_sub_621_n77;
  tri   P2_sub_621_n76;
  tri   P2_sub_621_n75;
  tri   P2_sub_621_n73;
  tri   P2_sub_621_n72;
  tri   P2_sub_621_n71;
  tri   P2_sub_621_n70;
  tri   P2_sub_621_n69;
  tri   P2_sub_621_n68;
  tri   P2_sub_621_n67;
  tri   P2_sub_621_n66;
  tri   P2_sub_621_n65;
  tri   P2_sub_621_n64;
  tri   P2_sub_621_n63;
  tri   P2_sub_621_n62;
  tri   P2_sub_621_n61;
  tri   P2_sub_621_n60;
  tri   P2_sub_621_n59;
  tri   P2_sub_621_n58;
  tri   P2_sub_621_n57;
  tri   P2_sub_621_n56;
  tri   P2_sub_621_n55;
  tri   P2_sub_621_n54;
  tri   P2_sub_621_n53;
  tri   P2_sub_621_n52;
  tri   P2_sub_621_n51;
  tri   P2_sub_621_n50;
  tri   P2_sub_621_n49;
  tri   P2_sub_621_n48;
  tri   P2_sub_621_n47;
  tri   P2_sub_621_n46;
  tri   P2_sub_621_n45;
  tri   P2_sub_621_n44;
  tri   P2_sub_621_n43;
  tri   P2_sub_621_n42;
  tri   P2_sub_621_n41;
  tri   P2_sub_621_n40;
  tri   P2_sub_621_n39;
  tri   P2_sub_621_n38;
  tri   P2_sub_621_n37;
  tri   P2_sub_621_n36;
  tri   P2_sub_621_n34;
  tri   P2_sub_621_n30;
  tri   P2_sub_621_n35;
  tri   P2_sub_621_n115;
  tri   P2_sub_621_n21;
  tri   P2_sub_621_n114;
  tri   P2_sub_621_n17;
  tri   P2_sub_621_n113;
  tri   P2_sub_621_n8;
  tri   P2_sub_621_n112;
  tri   P2_sub_621_n108;
  tri   P2_sub_621_n4;
  tri   P2_sub_621_n111;
  tri   P2_sub_621_n110;
  tri   P2_sub_621_n109;
  tri   r837_n75;
  tri   r837_n74;
  tri   r837_n71;
  tri   r837_n70;
  tri   r837_n69;
  tri   r837_n67;
  tri   r837_n68;
  tri   r837_n66;
  tri   r837_n65;
  tri   r837_n62;
  tri   r837_n61;
  tri   r837_n59;
  tri   r837_n58;
  tri   r837_n57;
  tri   r837_n55;
  tri   r837_n54;
  tri   r837_n52;
  tri   r837_n51;
  tri   r837_n50;
  tri   r837_n48;
  tri   r837_n47;
  tri   r837_n45;
  tri   r837_n44;
  tri   r837_n43;
  tri   r837_n41;
  tri   r837_n40;
  tri   r837_n38;
  tri   r837_n37;
  tri   r837_n36;
  tri   r837_n34;
  tri   r837_n33;
  tri   r837_n31;
  tri   r837_n30;
  tri   r837_n29;
  tri   r837_n27;
  tri   r837_n26;
  tri   r837_n24;
  tri   r837_n23;
  tri   r837_n22;
  tri   r837_n20;
  tri   r837_n19;
  tri   r837_n17;
  tri   r837_n16;
  tri   r837_n15;
  tri   r837_n13;
  tri   r837_n12;
  tri   r837_n10;
  tri   r837_n9;
  tri   r837_n8;
  tri   r837_n6;
  tri   r837_n5;
  tri   r837_n3;
  tri   r837_n2;
  tri   r837_n1;
  tri   r837_n158;
  tri   r837_n157;
  tri   r837_n156;
  tri   r837_n155;
  tri   r837_n154;
  tri   r837_n152;
  tri   r837_n151;
  tri   r837_n150;
  tri   r837_n149;
  tri   r837_n148;
  tri   r837_n147;
  tri   r837_n146;
  tri   r837_n145;
  tri   r837_n144;
  tri   r837_n142;
  tri   r837_n141;
  tri   r837_n140;
  tri   r837_n139;
  tri   r837_n138;
  tri   r837_n137;
  tri   r837_n136;
  tri   r837_n135;
  tri   r837_n134;
  tri   r837_n132;
  tri   r837_n131;
  tri   r837_n130;
  tri   r837_n129;
  tri   r837_n128;
  tri   r837_n127;
  tri   r837_n126;
  tri   r837_n125;
  tri   r837_n124;
  tri   r837_n122;
  tri   r837_n121;
  tri   r837_n120;
  tri   r837_n119;
  tri   r837_n118;
  tri   r837_n117;
  tri   r837_n116;
  tri   r837_n115;
  tri   r837_n114;
  tri   r837_n112;
  tri   r837_n111;
  tri   r837_n110;
  tri   r837_n109;
  tri   r837_n108;
  tri   r837_n107;
  tri   r837_n106;
  tri   r837_n105;
  tri   r837_n104;
  tri   r837_n102;
  tri   r837_n101;
  tri   r837_n100;
  tri   r837_n99;
  tri   r837_n98;
  tri   r837_n97;
  tri   r837_n96;
  tri   r837_n95;
  tri   r837_n94;
  tri   r837_n92;
  tri   r837_n91;
  tri   r837_n90;
  tri   r837_n89;
  tri   r837_n88;
  tri   r837_n87;
  tri   r837_n86;
  tri   r837_n85;
  tri   r837_n84;
  tri   r837_n82;
  tri   r837_n81;
  tri   r837_n80;
  tri   r837_n79;
  tri   r837_n73;
  tri   r837_n78;
  tri   r837_n77;
  tri   r837_n191;
  tri   r837_n190;
  tri   r837_n159;
  tri   r837_n189;
  tri   r837_n188;
  tri   r837_n60;
  tri   r837_n187;
  tri   r837_n186;
  tri   r837_n185;
  tri   r837_n184;
  tri   r837_n53;
  tri   r837_n183;
  tri   r837_n182;
  tri   r837_n181;
  tri   r837_n46;
  tri   r837_n180;
  tri   r837_n179;
  tri   r837_n178;
  tri   r837_n39;
  tri   r837_n177;
  tri   r837_n176;
  tri   r837_n175;
  tri   r837_n32;
  tri   r837_n174;
  tri   r837_n173;
  tri   r837_n172;
  tri   r837_n25;
  tri   r837_n171;
  tri   r837_n170;
  tri   r837_n169;
  tri   r837_n18;
  tri   r837_n168;
  tri   r837_n167;
  tri   r837_n166;
  tri   r837_n11;
  tri   r837_n14;
  tri   r837_n165;
  tri   r837_n164;
  tri   r837_n163;
  tri   r837_n160;
  tri   r837_n4;
  tri   r837_n161;
  tri   r837_n162;
  tri   r838_n98;
  tri   r838_n96;
  tri   r838_n95;
  tri   r838_n92;
  tri   r838_n91;
  tri   r838_n90;
  tri   r838_n89;
  tri   r838_n88;
  tri   r838_n87;
  tri   r838_n86;
  tri   r838_n85;
  tri   r838_n84;
  tri   r838_n82;
  tri   r838_n81;
  tri   r838_n80;
  tri   r838_n79;
  tri   r838_n78;
  tri   r838_n77;
  tri   r838_n75;
  tri   r838_n74;
  tri   r838_n73;
  tri   r838_n71;
  tri   r838_n70;
  tri   r838_n69;
  tri   r838_n67;
  tri   r838_n68;
  tri   r838_n66;
  tri   r838_n65;
  tri   r838_n62;
  tri   r838_n61;
  tri   r838_n59;
  tri   r838_n58;
  tri   r838_n57;
  tri   r838_n55;
  tri   r838_n54;
  tri   r838_n52;
  tri   r838_n51;
  tri   r838_n50;
  tri   r838_n48;
  tri   r838_n47;
  tri   r838_n45;
  tri   r838_n44;
  tri   r838_n43;
  tri   r838_n41;
  tri   r838_n40;
  tri   r838_n38;
  tri   r838_n37;
  tri   r838_n36;
  tri   r838_n34;
  tri   r838_n33;
  tri   r838_n31;
  tri   r838_n30;
  tri   r838_n29;
  tri   r838_n27;
  tri   r838_n26;
  tri   r838_n24;
  tri   r838_n23;
  tri   r838_n22;
  tri   r838_n20;
  tri   r838_n19;
  tri   r838_n17;
  tri   r838_n16;
  tri   r838_n15;
  tri   r838_n13;
  tri   r838_n12;
  tri   r838_n10;
  tri   r838_n9;
  tri   r838_n8;
  tri   r838_n6;
  tri   r838_n5;
  tri   r838_n3;
  tri   r838_n2;
  tri   r838_n1;
  tri   r838_n32;
  tri   r838_n174;
  tri   r838_n173;
  tri   r838_n172;
  tri   r838_n25;
  tri   r838_n171;
  tri   r838_n170;
  tri   r838_n169;
  tri   r838_n18;
  tri   r838_n168;
  tri   r838_n167;
  tri   r838_n166;
  tri   r838_n11;
  tri   r838_n165;
  tri   r838_n164;
  tri   r838_n163;
  tri   r838_n4;
  tri   r838_n162;
  tri   r838_n161;
  tri   r838_n160;
  tri   r838_n158;
  tri   r838_n157;
  tri   r838_n156;
  tri   r838_n155;
  tri   r838_n154;
  tri   r838_n152;
  tri   r838_n151;
  tri   r838_n150;
  tri   r838_n149;
  tri   r838_n148;
  tri   r838_n147;
  tri   r838_n146;
  tri   r838_n145;
  tri   r838_n144;
  tri   r838_n142;
  tri   r838_n141;
  tri   r838_n140;
  tri   r838_n139;
  tri   r838_n138;
  tri   r838_n137;
  tri   r838_n136;
  tri   r838_n135;
  tri   r838_n134;
  tri   r838_n132;
  tri   r838_n131;
  tri   r838_n130;
  tri   r838_n129;
  tri   r838_n128;
  tri   r838_n127;
  tri   r838_n126;
  tri   r838_n125;
  tri   r838_n124;
  tri   r838_n122;
  tri   r838_n121;
  tri   r838_n120;
  tri   r838_n119;
  tri   r838_n118;
  tri   r838_n117;
  tri   r838_n116;
  tri   r838_n115;
  tri   r838_n114;
  tri   r838_n112;
  tri   r838_n111;
  tri   r838_n110;
  tri   r838_n109;
  tri   r838_n108;
  tri   r838_n107;
  tri   r838_n106;
  tri   r838_n105;
  tri   r838_n104;
  tri   r838_n102;
  tri   r838_n101;
  tri   r838_n100;
  tri   r838_n97;
  tri   r838_n94;
  tri   r838_n99;
  tri   r838_n191;
  tri   r838_n190;
  tri   r838_n159;
  tri   r838_n189;
  tri   r838_n188;
  tri   r838_n60;
  tri   r838_n187;
  tri   r838_n186;
  tri   r838_n185;
  tri   r838_n184;
  tri   r838_n53;
  tri   r838_n183;
  tri   r838_n182;
  tri   r838_n181;
  tri   r838_n46;
  tri   r838_n180;
  tri   r838_n179;
  tri   r838_n178;
  tri   r838_n175;
  tri   r838_n39;
  tri   r838_n176;
  tri   r838_n177;
  tri   P2_sub_632_n54;
  tri   P2_sub_632_n53;
  tri   P2_sub_632_n52;
  tri   P2_sub_632_n51;
  tri   P2_sub_632_n50;
  tri   P2_sub_632_n49;
  tri   P2_sub_632_n48;
  tri   P2_sub_632_n47;
  tri   P2_sub_632_n46;
  tri   P2_sub_632_n45;
  tri   P2_sub_632_n44;
  tri   P2_sub_632_n43;
  tri   P2_sub_632_n42;
  tri   P2_sub_632_n41;
  tri   P2_sub_632_n40;
  tri   P2_sub_632_n39;
  tri   P2_sub_632_n38;
  tri   P2_sub_632_n37;
  tri   P2_sub_632_n36;
  tri   P2_sub_632_n35;
  tri   P2_sub_632_n34;
  tri   P2_sub_632_n33;
  tri   P2_sub_632_n32;
  tri   P2_sub_632_n31;
  tri   P2_sub_632_n30;
  tri   P2_sub_632_n29;
  tri   P2_sub_632_n28;
  tri   P2_sub_632_n27;
  tri   P2_sub_632_n26;
  tri   P2_sub_632_n25;
  tri   P2_sub_632_n24;
  tri   P2_sub_632_n23;
  tri   P2_sub_632_n22;
  tri   P2_sub_632_n21;
  tri   P2_sub_632_n20;
  tri   P2_sub_632_n19;
  tri   P2_sub_632_n18;
  tri   P2_sub_632_n17;
  tri   P2_sub_632_n16;
  tri   P2_sub_632_n14;
  tri   P2_sub_632_n12;
  tri   P2_sub_632_n10;
  tri   P2_sub_632_n8;
  tri   P2_sub_632_n7;
  tri   P2_sub_632_n6;
  tri   P2_sub_632_n5;
  tri   P2_sub_632_n15;
  tri   P2_sub_632_n13;
  tri   P2_sub_632_n9;
  tri   P2_sub_632_n11;
  tri   add_1108_n309;
  tri   add_1108_n308;
  tri   add_1108_n310;
  tri   add_1108_n303;
  tri   add_1108_n304;
  tri   add_1108_n302;
  tri   add_1108_n305;
  tri   add_1108_n306;
  tri   add_1108_n307;
  tri   add_1108_n297;
  tri   add_1108_n298;
  tri   add_1108_n296;
  tri   add_1108_n299;
  tri   add_1108_n300;
  tri   add_1108_n301;
  tri   add_1108_n291;
  tri   add_1108_n292;
  tri   add_1108_n290;
  tri   add_1108_n293;
  tri   add_1108_n294;
  tri   add_1108_n295;
  tri   add_1108_n285;
  tri   add_1108_n286;
  tri   add_1108_n284;
  tri   add_1108_n287;
  tri   add_1108_n288;
  tri   add_1108_n289;
  tri   add_1108_n277;
  tri   add_1108_n279;
  tri   add_1108_n278;
  tri   add_1108_n280;
  tri   add_1108_n281;
  tri   add_1108_n282;
  tri   add_1108_n283;
  tri   add_1108_n270;
  tri   add_1108_n272;
  tri   add_1108_n273;
  tri   add_1108_n271;
  tri   add_1108_n274;
  tri   add_1108_n276;
  tri   add_1108_n275;
  tri   add_1108_n262;
  tri   add_1108_n263;
  tri   add_1108_n261;
  tri   add_1108_n266;
  tri   add_1108_n264;
  tri   add_1108_n265;
  tri   add_1108_n267;
  tri   add_1108_n269;
  tri   add_1108_n268;
  tri   add_1108_n256;
  tri   add_1108_n255;
  tri   add_1108_n257;
  tri   add_1108_n259;
  tri   add_1108_n258;
  tri   add_1108_n260;
  tri   add_1108_n249;
  tri   add_1108_n248;
  tri   add_1108_n250;
  tri   add_1108_n251;
  tri   add_1108_n252;
  tri   add_1108_n253;
  tri   add_1108_n254;
  tri   add_1108_n242;
  tri   add_1108_n243;
  tri   add_1108_n241;
  tri   add_1108_n245;
  tri   add_1108_n246;
  tri   add_1108_n247;
  tri   add_1108_n244;
  tri   add_1108_n233;
  tri   add_1108_n236;
  tri   add_1108_n234;
  tri   add_1108_n235;
  tri   add_1108_n237;
  tri   add_1108_n238;
  tri   add_1108_n239;
  tri   add_1108_n240;
  tri   add_1108_n226;
  tri   add_1108_n225;
  tri   add_1108_n227;
  tri   add_1108_n229;
  tri   add_1108_n228;
  tri   add_1108_n230;
  tri   add_1108_n232;
  tri   add_1108_n231;
  tri   add_1108_n219;
  tri   add_1108_n218;
  tri   add_1108_n220;
  tri   add_1108_n222;
  tri   add_1108_n223;
  tri   add_1108_n221;
  tri   add_1108_n224;
  tri   add_1108_n212;
  tri   add_1108_n213;
  tri   add_1108_n211;
  tri   add_1108_n216;
  tri   add_1108_n217;
  tri   add_1108_n214;
  tri   add_1108_n215;
  tri   add_1108_n206;
  tri   add_1108_n204;
  tri   add_1108_n205;
  tri   add_1108_n207;
  tri   add_1108_n209;
  tri   add_1108_n208;
  tri   add_1108_n210;
  tri   add_1108_n197;
  tri   add_1108_n199;
  tri   add_1108_n198;
  tri   add_1108_n200;
  tri   add_1108_n201;
  tri   add_1108_n202;
  tri   add_1108_n203;
  tri   add_1108_n190;
  tri   add_1108_n192;
  tri   add_1108_n193;
  tri   add_1108_n191;
  tri   add_1108_n194;
  tri   add_1108_n196;
  tri   add_1108_n195;
  tri   add_1108_n183;
  tri   add_1108_n182;
  tri   add_1108_n184;
  tri   add_1108_n186;
  tri   add_1108_n185;
  tri   add_1108_n187;
  tri   add_1108_n189;
  tri   add_1108_n188;
  tri   add_1108_n175;
  tri   add_1108_n176;
  tri   add_1108_n174;
  tri   add_1108_n177;
  tri   add_1108_n178;
  tri   add_1108_n179;
  tri   add_1108_n180;
  tri   add_1108_n181;
  tri   add_1108_n166;
  tri   add_1108_n169;
  tri   add_1108_n167;
  tri   add_1108_n168;
  tri   add_1108_n170;
  tri   add_1108_n171;
  tri   add_1108_n172;
  tri   add_1108_n173;
  tri   add_1108_n159;
  tri   add_1108_n158;
  tri   add_1108_n160;
  tri   add_1108_n162;
  tri   add_1108_n161;
  tri   add_1108_n163;
  tri   add_1108_n165;
  tri   add_1108_n164;
  tri   add_1108_n152;
  tri   add_1108_n151;
  tri   add_1108_n153;
  tri   add_1108_n155;
  tri   add_1108_n156;
  tri   add_1108_n154;
  tri   add_1108_n157;
  tri   add_1108_n145;
  tri   add_1108_n146;
  tri   add_1108_n144;
  tri   add_1108_n149;
  tri   add_1108_n150;
  tri   add_1108_n147;
  tri   add_1108_n148;
  tri   add_1108_n139;
  tri   add_1108_n137;
  tri   add_1108_n138;
  tri   add_1108_n140;
  tri   add_1108_n142;
  tri   add_1108_n141;
  tri   add_1108_n143;
  tri   add_1108_n130;
  tri   add_1108_n132;
  tri   add_1108_n131;
  tri   add_1108_n133;
  tri   add_1108_n134;
  tri   add_1108_n135;
  tri   add_1108_n136;
  tri   add_1108_n123;
  tri   add_1108_n125;
  tri   add_1108_n126;
  tri   add_1108_n124;
  tri   add_1108_n127;
  tri   add_1108_n129;
  tri   add_1108_n128;
  tri   add_1108_n115;
  tri   add_1108_n116;
  tri   add_1108_n114;
  tri   add_1108_n119;
  tri   add_1108_n117;
  tri   add_1108_n118;
  tri   add_1108_n120;
  tri   add_1108_n122;
  tri   add_1108_n121;
  tri   add_1108_n109;
  tri   add_1108_n108;
  tri   add_1108_n110;
  tri   add_1108_n112;
  tri   add_1108_n111;
  tri   add_1108_n113;
  tri   add_1108_n102;
  tri   add_1108_n101;
  tri   add_1108_n103;
  tri   add_1108_n104;
  tri   add_1108_n105;
  tri   add_1108_n106;
  tri   add_1108_n107;
  tri   add_1108_n95;
  tri   add_1108_n96;
  tri   add_1108_n94;
  tri   add_1108_n98;
  tri   add_1108_n99;
  tri   add_1108_n100;
  tri   add_1108_n97;
  tri   add_1108_n86;
  tri   add_1108_n89;
  tri   add_1108_n87;
  tri   add_1108_n88;
  tri   add_1108_n90;
  tri   add_1108_n91;
  tri   add_1108_n92;
  tri   add_1108_n93;
  tri   add_1108_n79;
  tri   add_1108_n78;
  tri   add_1108_n80;
  tri   add_1108_n82;
  tri   add_1108_n81;
  tri   add_1108_n83;
  tri   add_1108_n85;
  tri   add_1108_n84;
  tri   add_1108_n72;
  tri   add_1108_n73;
  tri   add_1108_n71;
  tri   add_1108_n74;
  tri   add_1108_n76;
  tri   add_1108_n75;
  tri   add_1108_n77;
  tri   add_1108_n65;
  tri   add_1108_n64;
  tri   add_1108_n66;
  tri   add_1108_n67;
  tri   add_1108_n68;
  tri   add_1108_n69;
  tri   add_1108_n70;
  tri   add_1108_n59;
  tri   add_1108_n58;
  tri   add_1108_n60;
  tri   add_1108_n61;
  tri   add_1108_n62;
  tri   add_1108_n63;
  tri   add_1108_n57;
  tri   add_1108_n49;
  tri   add_1108_n51;
  tri   add_1108_n53;
  tri   add_1108_n50;
  tri   add_1108_n52;
  tri   add_1108_n54;
  tri   add_1108_n55;
  tri   add_1108_n56;
  tri   add_1108_n41;
  tri   add_1108_n40;
  tri   add_1108_n42;
  tri   add_1108_n44;
  tri   add_1108_n45;
  tri   add_1108_n43;
  tri   add_1108_n46;
  tri   add_1108_n48;
  tri   add_1108_n47;
  tri   add_1108_n34;
  tri   add_1108_n33;
  tri   add_1108_n35;
  tri   add_1108_n37;
  tri   add_1108_n39;
  tri   add_1108_n38;
  tri   add_1108_n36;
  tri   add_1108_n24;
  tri   add_1108_n25;
  tri   add_1108_n27;
  tri   add_1108_n26;
  tri   add_1108_n28;
  tri   add_1108_n29;
  tri   add_1108_n30;
  tri   add_1108_n32;
  tri   add_1108_n31;
  tri   add_1108_n16;
  tri   add_1108_n17;
  tri   add_1108_n15;
  tri   add_1108_n18;
  tri   add_1108_n20;
  tri   add_1108_n19;
  tri   add_1108_n21;
  tri   add_1108_n23;
  tri   add_1108_n22;
  tri   add_1108_n9;
  tri   add_1108_n10;
  tri   add_1108_n8;
  tri   add_1108_n11;
  tri   add_1108_n13;
  tri   add_1108_n12;
  tri   add_1108_n14;
  tri   add_1108_n2;
  tri   add_1108_n3;
  tri   add_1108_n1;
  tri   add_1108_n4;
  tri   add_1108_n6;
  tri   add_1108_n5;
  tri   add_1108_n7;
  tri   r839_n94;
  tri   r839_n93;
  tri   r839_n92;
  tri   r839_n91;
  tri   r839_n90;
  tri   r839_n89;
  tri   r839_n88;
  tri   r839_n87;
  tri   r839_n86;
  tri   r839_n84;
  tri   r839_n83;
  tri   r839_n82;
  tri   r839_n81;
  tri   r839_n80;
  tri   r839_n79;
  tri   r839_n78;
  tri   r839_n77;
  tri   r839_n76;
  tri   r839_n75;
  tri   r839_n74;
  tri   r839_n73;
  tri   r839_n72;
  tri   r839_n71;
  tri   r839_n70;
  tri   r839_n69;
  tri   r839_n67;
  tri   r839_n66;
  tri   r839_n65;
  tri   r839_n64;
  tri   r839_n63;
  tri   r839_n62;
  tri   r839_n61;
  tri   r839_n59;
  tri   r839_n60;
  tri   r839_n58;
  tri   r839_n57;
  tri   r839_n55;
  tri   r839_n54;
  tri   r839_n52;
  tri   r839_n51;
  tri   r839_n50;
  tri   r839_n48;
  tri   r839_n47;
  tri   r839_n45;
  tri   r839_n44;
  tri   r839_n43;
  tri   r839_n41;
  tri   r839_n40;
  tri   r839_n38;
  tri   r839_n37;
  tri   r839_n36;
  tri   r839_n34;
  tri   r839_n33;
  tri   r839_n31;
  tri   r839_n30;
  tri   r839_n29;
  tri   r839_n27;
  tri   r839_n26;
  tri   r839_n24;
  tri   r839_n23;
  tri   r839_n22;
  tri   r839_n20;
  tri   r839_n19;
  tri   r839_n17;
  tri   r839_n16;
  tri   r839_n15;
  tri   r839_n13;
  tri   r839_n12;
  tri   r839_n10;
  tri   r839_n9;
  tri   r839_n8;
  tri   r839_n6;
  tri   r839_n5;
  tri   r839_n3;
  tri   r839_n2;
  tri   r839_n1;
  tri   r839_n182;
  tri   r839_n181;
  tri   r839_n180;
  tri   r839_n178;
  tri   r839_n177;
  tri   r839_n176;
  tri   r839_n175;
  tri   r839_n174;
  tri   r839_n172;
  tri   r839_n171;
  tri   r839_n170;
  tri   r839_n169;
  tri   r839_n168;
  tri   r839_n167;
  tri   r839_n164;
  tri   r839_n163;
  tri   r839_n161;
  tri   r839_n160;
  tri   r839_n159;
  tri   r839_n158;
  tri   r839_n157;
  tri   r839_n156;
  tri   r839_n155;
  tri   r839_n154;
  tri   r839_n153;
  tri   r839_n152;
  tri   r839_n151;
  tri   r839_n150;
  tri   r839_n149;
  tri   r839_n148;
  tri   r839_n147;
  tri   r839_n146;
  tri   r839_n145;
  tri   r839_n144;
  tri   r839_n143;
  tri   r839_n142;
  tri   r839_n141;
  tri   r839_n140;
  tri   r839_n139;
  tri   r839_n138;
  tri   r839_n137;
  tri   r839_n136;
  tri   r839_n135;
  tri   r839_n134;
  tri   r839_n133;
  tri   r839_n132;
  tri   r839_n131;
  tri   r839_n130;
  tri   r839_n129;
  tri   r839_n128;
  tri   r839_n127;
  tri   r839_n126;
  tri   r839_n125;
  tri   r839_n124;
  tri   r839_n123;
  tri   r839_n122;
  tri   r839_n121;
  tri   r839_n120;
  tri   r839_n119;
  tri   r839_n118;
  tri   r839_n117;
  tri   r839_n116;
  tri   r839_n115;
  tri   r839_n114;
  tri   r839_n113;
  tri   r839_n112;
  tri   r839_n111;
  tri   r839_n110;
  tri   r839_n109;
  tri   r839_n95;
  tri   r839_n108;
  tri   r839_n107;
  tri   r839_n106;
  tri   r839_n105;
  tri   r839_n104;
  tri   r839_n103;
  tri   r839_n102;
  tri   r839_n101;
  tri   r839_n96;
  tri   r839_n100;
  tri   r839_n99;
  tri   r839_n97;
  tri   r839_n98;
  tri   r839_n85;
  tri   r839_n14;
  tri   r839_n265;
  tri   r839_n264;
  tri   r839_n4;
  tri   r839_n7;
  tri   r839_n262;
  tri   r839_n261;
  tri   r839_n260;
  tri   r839_n258;
  tri   r839_n257;
  tri   r839_n256;
  tri   r839_n255;
  tri   r839_n254;
  tri   r839_n252;
  tri   r839_n251;
  tri   r839_n250;
  tri   r839_n249;
  tri   r839_n248;
  tri   r839_n247;
  tri   r839_n246;
  tri   r839_n245;
  tri   r839_n244;
  tri   r839_n243;
  tri   r839_n242;
  tri   r839_n241;
  tri   r839_n240;
  tri   r839_n239;
  tri   r839_n238;
  tri   r839_n237;
  tri   r839_n236;
  tri   r839_n235;
  tri   r839_n234;
  tri   r839_n233;
  tri   r839_n232;
  tri   r839_n231;
  tri   r839_n230;
  tri   r839_n229;
  tri   r839_n228;
  tri   r839_n227;
  tri   r839_n226;
  tri   r839_n225;
  tri   r839_n224;
  tri   r839_n223;
  tri   r839_n222;
  tri   r839_n221;
  tri   r839_n220;
  tri   r839_n219;
  tri   r839_n218;
  tri   r839_n217;
  tri   r839_n216;
  tri   r839_n215;
  tri   r839_n214;
  tri   r839_n213;
  tri   r839_n212;
  tri   r839_n211;
  tri   r839_n210;
  tri   r839_n209;
  tri   r839_n208;
  tri   r839_n207;
  tri   r839_n206;
  tri   r839_n205;
  tri   r839_n204;
  tri   r839_n203;
  tri   r839_n202;
  tri   r839_n201;
  tri   r839_n200;
  tri   r839_n199;
  tri   r839_n198;
  tri   r839_n197;
  tri   r839_n183;
  tri   r839_n196;
  tri   r839_n195;
  tri   r839_n194;
  tri   r839_n193;
  tri   r839_n192;
  tri   r839_n191;
  tri   r839_n190;
  tri   r839_n189;
  tri   r839_n184;
  tri   r839_n188;
  tri   r839_n187;
  tri   r839_n173;
  tri   r839_n179;
  tri   r839_n186;
  tri   r839_n185;
  tri   r839_n291;
  tri   r839_n290;
  tri   r839_n253;
  tri   r839_n259;
  tri   r839_n289;
  tri   r839_n288;
  tri   r839_n162;
  tri   r839_n287;
  tri   r839_n166;
  tri   r839_n286;
  tri   r839_n285;
  tri   r839_n284;
  tri   r839_n53;
  tri   r839_n56;
  tri   r839_n283;
  tri   r839_n282;
  tri   r839_n281;
  tri   r839_n46;
  tri   r839_n49;
  tri   r839_n280;
  tri   r839_n279;
  tri   r839_n278;
  tri   r839_n39;
  tri   r839_n42;
  tri   r839_n277;
  tri   r839_n276;
  tri   r839_n275;
  tri   r839_n32;
  tri   r839_n35;
  tri   r839_n274;
  tri   r839_n273;
  tri   r839_n272;
  tri   r839_n25;
  tri   r839_n28;
  tri   r839_n271;
  tri   r839_n270;
  tri   r839_n269;
  tri   r839_n18;
  tri   r839_n21;
  tri   r839_n268;
  tri   r839_n267;
  tri   r839_n266;
  tri   r839_n263;
  tri   r839_n11;
  tri   r841_n44;
  tri   r841_n41;
  tri   r841_n40;
  tri   r841_n38;
  tri   r841_n37;
  tri   r841_n36;
  tri   r841_n34;
  tri   r841_n33;
  tri   r841_n31;
  tri   r841_n30;
  tri   r841_n29;
  tri   r841_n27;
  tri   r841_n26;
  tri   r841_n24;
  tri   r841_n23;
  tri   r841_n22;
  tri   r841_n20;
  tri   r841_n19;
  tri   r841_n17;
  tri   r841_n16;
  tri   r841_n15;
  tri   r841_n13;
  tri   r841_n12;
  tri   r841_n10;
  tri   r841_n9;
  tri   r841_n8;
  tri   r841_n6;
  tri   r841_n5;
  tri   r841_n3;
  tri   r841_n2;
  tri   r841_n1;
  tri   r841_n134;
  tri   r841_n133;
  tri   r841_n130;
  tri   r841_n129;
  tri   r841_n128;
  tri   r841_n127;
  tri   r841_n126;
  tri   r841_n124;
  tri   r841_n123;
  tri   r841_n122;
  tri   r841_n121;
  tri   r841_n120;
  tri   r841_n119;
  tri   r841_n118;
  tri   r841_n117;
  tri   r841_n116;
  tri   r841_n115;
  tri   r841_n114;
  tri   r841_n113;
  tri   r841_n112;
  tri   r841_n111;
  tri   r841_n110;
  tri   r841_n109;
  tri   r841_n108;
  tri   r841_n107;
  tri   r841_n106;
  tri   r841_n105;
  tri   r841_n104;
  tri   r841_n103;
  tri   r841_n102;
  tri   r841_n101;
  tri   r841_n100;
  tri   r841_n99;
  tri   r841_n98;
  tri   r841_n97;
  tri   r841_n96;
  tri   r841_n95;
  tri   r841_n94;
  tri   r841_n93;
  tri   r841_n92;
  tri   r841_n91;
  tri   r841_n90;
  tri   r841_n89;
  tri   r841_n88;
  tri   r841_n87;
  tri   r841_n86;
  tri   r841_n85;
  tri   r841_n84;
  tri   r841_n83;
  tri   r841_n82;
  tri   r841_n81;
  tri   r841_n80;
  tri   r841_n79;
  tri   r841_n78;
  tri   r841_n77;
  tri   r841_n76;
  tri   r841_n75;
  tri   r841_n74;
  tri   r841_n73;
  tri   r841_n72;
  tri   r841_n71;
  tri   r841_n70;
  tri   r841_n69;
  tri   r841_n67;
  tri   r841_n66;
  tri   r841_n65;
  tri   r841_n64;
  tri   r841_n63;
  tri   r841_n62;
  tri   r841_n61;
  tri   r841_n59;
  tri   r841_n60;
  tri   r841_n58;
  tri   r841_n57;
  tri   r841_n55;
  tri   r841_n54;
  tri   r841_n52;
  tri   r841_n51;
  tri   r841_n50;
  tri   r841_n48;
  tri   r841_n47;
  tri   r841_n43;
  tri   r841_n45;
  tri   r841_n221;
  tri   r841_n218;
  tri   r841_n217;
  tri   r841_n216;
  tri   r841_n215;
  tri   r841_n214;
  tri   r841_n212;
  tri   r841_n211;
  tri   r841_n210;
  tri   r841_n209;
  tri   r841_n208;
  tri   r841_n207;
  tri   r841_n206;
  tri   r841_n205;
  tri   r841_n204;
  tri   r841_n203;
  tri   r841_n202;
  tri   r841_n201;
  tri   r841_n200;
  tri   r841_n199;
  tri   r841_n198;
  tri   r841_n197;
  tri   r841_n196;
  tri   r841_n195;
  tri   r841_n194;
  tri   r841_n193;
  tri   r841_n192;
  tri   r841_n191;
  tri   r841_n190;
  tri   r841_n189;
  tri   r841_n188;
  tri   r841_n187;
  tri   r841_n186;
  tri   r841_n185;
  tri   r841_n184;
  tri   r841_n183;
  tri   r841_n182;
  tri   r841_n181;
  tri   r841_n180;
  tri   r841_n179;
  tri   r841_n178;
  tri   r841_n177;
  tri   r841_n176;
  tri   r841_n175;
  tri   r841_n174;
  tri   r841_n173;
  tri   r841_n172;
  tri   r841_n171;
  tri   r841_n170;
  tri   r841_n169;
  tri   r841_n168;
  tri   r841_n167;
  tri   r841_n164;
  tri   r841_n163;
  tri   r841_n161;
  tri   r841_n160;
  tri   r841_n159;
  tri   r841_n158;
  tri   r841_n157;
  tri   r841_n156;
  tri   r841_n155;
  tri   r841_n154;
  tri   r841_n153;
  tri   r841_n152;
  tri   r841_n151;
  tri   r841_n150;
  tri   r841_n149;
  tri   r841_n135;
  tri   r841_n148;
  tri   r841_n147;
  tri   r841_n146;
  tri   r841_n145;
  tri   r841_n144;
  tri   r841_n143;
  tri   r841_n142;
  tri   r841_n141;
  tri   r841_n140;
  tri   r841_n139;
  tri   r841_n125;
  tri   r841_n131;
  tri   r841_n138;
  tri   r841_n137;
  tri   r841_n132;
  tri   r841_n136;
  tri   r841_n289;
  tri   r841_n288;
  tri   r841_n166;
  tri   r841_n286;
  tri   r841_n285;
  tri   r841_n284;
  tri   r841_n53;
  tri   r841_n56;
  tri   r841_n283;
  tri   r841_n282;
  tri   r841_n281;
  tri   r841_n46;
  tri   r841_n49;
  tri   r841_n280;
  tri   r841_n279;
  tri   r841_n278;
  tri   r841_n39;
  tri   r841_n42;
  tri   r841_n277;
  tri   r841_n276;
  tri   r841_n275;
  tri   r841_n32;
  tri   r841_n35;
  tri   r841_n274;
  tri   r841_n273;
  tri   r841_n272;
  tri   r841_n25;
  tri   r841_n28;
  tri   r841_n271;
  tri   r841_n270;
  tri   r841_n269;
  tri   r841_n18;
  tri   r841_n21;
  tri   r841_n268;
  tri   r841_n267;
  tri   r841_n266;
  tri   r841_n11;
  tri   r841_n14;
  tri   r841_n265;
  tri   r841_n264;
  tri   r841_n263;
  tri   r841_n4;
  tri   r841_n7;
  tri   r841_n262;
  tri   r841_n261;
  tri   r841_n260;
  tri   r841_n259;
  tri   r841_n258;
  tri   r841_n257;
  tri   r841_n256;
  tri   r841_n255;
  tri   r841_n254;
  tri   r841_n253;
  tri   r841_n252;
  tri   r841_n251;
  tri   r841_n250;
  tri   r841_n249;
  tri   r841_n248;
  tri   r841_n247;
  tri   r841_n246;
  tri   r841_n245;
  tri   r841_n244;
  tri   r841_n243;
  tri   r841_n242;
  tri   r841_n241;
  tri   r841_n240;
  tri   r841_n239;
  tri   r841_n238;
  tri   r841_n237;
  tri   r841_n223;
  tri   r841_n236;
  tri   r841_n235;
  tri   r841_n234;
  tri   r841_n233;
  tri   r841_n232;
  tri   r841_n231;
  tri   r841_n230;
  tri   r841_n229;
  tri   r841_n228;
  tri   r841_n227;
  tri   r841_n213;
  tri   r841_n219;
  tri   r841_n226;
  tri   r841_n225;
  tri   r841_n220;
  tri   r841_n222;
  tri   r841_n224;
  tri   r841_n287;
  tri   r841_n162;
  tri   r841_n290;
  tri   r841_n291;
  tri   r843_n76;
  tri   r843_n75;
  tri   r843_n74;
  tri   r843_n72;
  tri   r843_n71;
  tri   r843_n70;
  tri   r843_n69;
  tri   r843_n68;
  tri   r843_n66;
  tri   r843_n65;
  tri   r843_n64;
  tri   r843_n63;
  tri   r843_n62;
  tri   r843_n61;
  tri   r843_n60;
  tri   r843_n59;
  tri   r843_n58;
  tri   r843_n57;
  tri   r843_n55;
  tri   r843_n54;
  tri   r843_n53;
  tri   r843_n51;
  tri   r843_n50;
  tri   r843_n48;
  tri   r843_n47;
  tri   r843_n46;
  tri   r843_n44;
  tri   r843_n43;
  tri   r843_n41;
  tri   r843_n40;
  tri   r843_n39;
  tri   r843_n37;
  tri   r843_n36;
  tri   r843_n34;
  tri   r843_n33;
  tri   r843_n32;
  tri   r843_n30;
  tri   r843_n29;
  tri   r843_n27;
  tri   r843_n26;
  tri   r843_n25;
  tri   r843_n23;
  tri   r843_n22;
  tri   r843_n20;
  tri   r843_n19;
  tri   r843_n18;
  tri   r843_n16;
  tri   r843_n15;
  tri   r843_n13;
  tri   r843_n12;
  tri   r843_n11;
  tri   r843_n9;
  tri   r843_n8;
  tri   r843_n6;
  tri   r843_n5;
  tri   r843_n4;
  tri   r843_n2;
  tri   r843_n1;
  tri   r843_n163;
  tri   r843_n162;
  tri   r843_n160;
  tri   r843_n159;
  tri   r843_n158;
  tri   r843_n156;
  tri   r843_n155;
  tri   r843_n154;
  tri   r843_n152;
  tri   r843_n151;
  tri   r843_n150;
  tri   r843_n149;
  tri   r843_n148;
  tri   r843_n147;
  tri   r843_n146;
  tri   r843_n145;
  tri   r843_n144;
  tri   r843_n142;
  tri   r843_n141;
  tri   r843_n140;
  tri   r843_n139;
  tri   r843_n138;
  tri   r843_n137;
  tri   r843_n136;
  tri   r843_n135;
  tri   r843_n134;
  tri   r843_n132;
  tri   r843_n131;
  tri   r843_n130;
  tri   r843_n129;
  tri   r843_n128;
  tri   r843_n127;
  tri   r843_n126;
  tri   r843_n125;
  tri   r843_n124;
  tri   r843_n122;
  tri   r843_n121;
  tri   r843_n120;
  tri   r843_n119;
  tri   r843_n118;
  tri   r843_n117;
  tri   r843_n116;
  tri   r843_n115;
  tri   r843_n114;
  tri   r843_n112;
  tri   r843_n111;
  tri   r843_n110;
  tri   r843_n109;
  tri   r843_n108;
  tri   r843_n107;
  tri   r843_n106;
  tri   r843_n105;
  tri   r843_n104;
  tri   r843_n102;
  tri   r843_n101;
  tri   r843_n100;
  tri   r843_n99;
  tri   r843_n98;
  tri   r843_n97;
  tri   r843_n96;
  tri   r843_n95;
  tri   r843_n94;
  tri   r843_n92;
  tri   r843_n91;
  tri   r843_n90;
  tri   r843_n89;
  tri   r843_n88;
  tri   r843_n87;
  tri   r843_n86;
  tri   r843_n85;
  tri   r843_n84;
  tri   r843_n82;
  tri   r843_n81;
  tri   r843_n78;
  tri   r843_n79;
  tri   r843_n80;
  tri   r843_n77;
  tri   r843_n249;
  tri   r843_n247;
  tri   r843_n246;
  tri   r843_n245;
  tri   r843_n243;
  tri   r843_n242;
  tri   r843_n241;
  tri   r843_n239;
  tri   r843_n238;
  tri   r843_n237;
  tri   r843_n236;
  tri   r843_n235;
  tri   r843_n234;
  tri   r843_n233;
  tri   r843_n232;
  tri   r843_n231;
  tri   r843_n229;
  tri   r843_n228;
  tri   r843_n227;
  tri   r843_n226;
  tri   r843_n225;
  tri   r843_n224;
  tri   r843_n223;
  tri   r843_n222;
  tri   r843_n221;
  tri   r843_n219;
  tri   r843_n218;
  tri   r843_n217;
  tri   r843_n216;
  tri   r843_n215;
  tri   r843_n214;
  tri   r843_n213;
  tri   r843_n212;
  tri   r843_n211;
  tri   r843_n209;
  tri   r843_n208;
  tri   r843_n207;
  tri   r843_n206;
  tri   r843_n205;
  tri   r843_n204;
  tri   r843_n203;
  tri   r843_n202;
  tri   r843_n201;
  tri   r843_n199;
  tri   r843_n198;
  tri   r843_n197;
  tri   r843_n196;
  tri   r843_n195;
  tri   r843_n194;
  tri   r843_n193;
  tri   r843_n192;
  tri   r843_n191;
  tri   r843_n189;
  tri   r843_n188;
  tri   r843_n187;
  tri   r843_n186;
  tri   r843_n185;
  tri   r843_n184;
  tri   r843_n183;
  tri   r843_n182;
  tri   r843_n181;
  tri   r843_n179;
  tri   r843_n178;
  tri   r843_n177;
  tri   r843_n176;
  tri   r843_n175;
  tri   r843_n174;
  tri   r843_n173;
  tri   r843_n172;
  tri   r843_n171;
  tri   r843_n169;
  tri   r843_n168;
  tri   r843_n167;
  tri   r843_n157;
  tri   r843_n166;
  tri   r843_n165;
  tri   r843_n289;
  tri   r843_n288;
  tri   r843_n161;
  tri   r843_n287;
  tri   r843_n286;
  tri   r843_n285;
  tri   r843_n52;
  tri   r843_n284;
  tri   r843_n283;
  tri   r843_n282;
  tri   r843_n45;
  tri   r843_n281;
  tri   r843_n280;
  tri   r843_n279;
  tri   r843_n38;
  tri   r843_n278;
  tri   r843_n277;
  tri   r843_n276;
  tri   r843_n31;
  tri   r843_n275;
  tri   r843_n274;
  tri   r843_n273;
  tri   r843_n24;
  tri   r843_n272;
  tri   r843_n271;
  tri   r843_n270;
  tri   r843_n17;
  tri   r843_n269;
  tri   r843_n268;
  tri   r843_n267;
  tri   r843_n10;
  tri   r843_n266;
  tri   r843_n265;
  tri   r843_n264;
  tri   r843_n3;
  tri   r843_n263;
  tri   r843_n262;
  tri   r843_n261;
  tri   r843_n259;
  tri   r843_n258;
  tri   r843_n257;
  tri   r843_n256;
  tri   r843_n255;
  tri   r843_n254;
  tri   r843_n253;
  tri   r843_n244;
  tri   r843_n252;
  tri   r843_n251;
  tri   r843_n248;
  tri   r800_n6;
  tri   r800_n3;
  tri   r800_n2;
  tri   r800_n1;
  tri   r800_n104;
  tri   r800_n103;
  tri   r800_n100;
  tri   r800_n99;
  tri   r800_n98;
  tri   r800_n97;
  tri   r800_n96;
  tri   r800_n94;
  tri   r800_n93;
  tri   r800_n92;
  tri   r800_n91;
  tri   r800_n90;
  tri   r800_n89;
  tri   r800_n88;
  tri   r800_n87;
  tri   r800_n86;
  tri   r800_n85;
  tri   r800_n84;
  tri   r800_n83;
  tri   r800_n82;
  tri   r800_n81;
  tri   r800_n80;
  tri   r800_n79;
  tri   r800_n78;
  tri   r800_n77;
  tri   r800_n76;
  tri   r800_n75;
  tri   r800_n74;
  tri   r800_n73;
  tri   r800_n72;
  tri   r800_n71;
  tri   r800_n70;
  tri   r800_n69;
  tri   r800_n67;
  tri   r800_n66;
  tri   r800_n65;
  tri   r800_n64;
  tri   r800_n63;
  tri   r800_n62;
  tri   r800_n61;
  tri   r800_n59;
  tri   r800_n60;
  tri   r800_n58;
  tri   r800_n57;
  tri   r800_n55;
  tri   r800_n54;
  tri   r800_n52;
  tri   r800_n51;
  tri   r800_n50;
  tri   r800_n48;
  tri   r800_n47;
  tri   r800_n45;
  tri   r800_n44;
  tri   r800_n43;
  tri   r800_n41;
  tri   r800_n40;
  tri   r800_n38;
  tri   r800_n37;
  tri   r800_n36;
  tri   r800_n34;
  tri   r800_n33;
  tri   r800_n31;
  tri   r800_n30;
  tri   r800_n29;
  tri   r800_n27;
  tri   r800_n26;
  tri   r800_n24;
  tri   r800_n23;
  tri   r800_n22;
  tri   r800_n20;
  tri   r800_n19;
  tri   r800_n17;
  tri   r800_n16;
  tri   r800_n15;
  tri   r800_n13;
  tri   r800_n12;
  tri   r800_n10;
  tri   r800_n9;
  tri   r800_n8;
  tri   r800_n5;
  tri   r800_n191;
  tri   r800_n188;
  tri   r800_n187;
  tri   r800_n186;
  tri   r800_n185;
  tri   r800_n184;
  tri   r800_n182;
  tri   r800_n181;
  tri   r800_n180;
  tri   r800_n179;
  tri   r800_n178;
  tri   r800_n177;
  tri   r800_n176;
  tri   r800_n175;
  tri   r800_n174;
  tri   r800_n173;
  tri   r800_n172;
  tri   r800_n171;
  tri   r800_n170;
  tri   r800_n169;
  tri   r800_n168;
  tri   r800_n167;
  tri   r800_n164;
  tri   r800_n163;
  tri   r800_n161;
  tri   r800_n160;
  tri   r800_n159;
  tri   r800_n158;
  tri   r800_n157;
  tri   r800_n156;
  tri   r800_n155;
  tri   r800_n154;
  tri   r800_n153;
  tri   r800_n152;
  tri   r800_n151;
  tri   r800_n150;
  tri   r800_n149;
  tri   r800_n148;
  tri   r800_n147;
  tri   r800_n146;
  tri   r800_n145;
  tri   r800_n144;
  tri   r800_n143;
  tri   r800_n142;
  tri   r800_n141;
  tri   r800_n140;
  tri   r800_n139;
  tri   r800_n138;
  tri   r800_n137;
  tri   r800_n136;
  tri   r800_n135;
  tri   r800_n134;
  tri   r800_n133;
  tri   r800_n132;
  tri   r800_n131;
  tri   r800_n130;
  tri   r800_n129;
  tri   r800_n128;
  tri   r800_n127;
  tri   r800_n126;
  tri   r800_n125;
  tri   r800_n124;
  tri   r800_n123;
  tri   r800_n122;
  tri   r800_n121;
  tri   r800_n120;
  tri   r800_n119;
  tri   r800_n105;
  tri   r800_n118;
  tri   r800_n117;
  tri   r800_n116;
  tri   r800_n115;
  tri   r800_n114;
  tri   r800_n113;
  tri   r800_n112;
  tri   r800_n111;
  tri   r800_n110;
  tri   r800_n109;
  tri   r800_n95;
  tri   r800_n101;
  tri   r800_n108;
  tri   r800_n107;
  tri   r800_n102;
  tri   r800_n106;
  tri   r800_n28;
  tri   r800_n270;
  tri   r800_n18;
  tri   r800_n21;
  tri   r800_n268;
  tri   r800_n267;
  tri   r800_n266;
  tri   r800_n11;
  tri   r800_n14;
  tri   r800_n265;
  tri   r800_n264;
  tri   r800_n263;
  tri   r800_n4;
  tri   r800_n7;
  tri   r800_n262;
  tri   r800_n261;
  tri   r800_n260;
  tri   r800_n258;
  tri   r800_n257;
  tri   r800_n256;
  tri   r800_n255;
  tri   r800_n254;
  tri   r800_n252;
  tri   r800_n251;
  tri   r800_n250;
  tri   r800_n249;
  tri   r800_n248;
  tri   r800_n247;
  tri   r800_n246;
  tri   r800_n245;
  tri   r800_n244;
  tri   r800_n243;
  tri   r800_n242;
  tri   r800_n241;
  tri   r800_n240;
  tri   r800_n239;
  tri   r800_n238;
  tri   r800_n237;
  tri   r800_n236;
  tri   r800_n235;
  tri   r800_n234;
  tri   r800_n233;
  tri   r800_n232;
  tri   r800_n231;
  tri   r800_n230;
  tri   r800_n229;
  tri   r800_n228;
  tri   r800_n227;
  tri   r800_n226;
  tri   r800_n225;
  tri   r800_n224;
  tri   r800_n223;
  tri   r800_n222;
  tri   r800_n221;
  tri   r800_n220;
  tri   r800_n219;
  tri   r800_n218;
  tri   r800_n217;
  tri   r800_n216;
  tri   r800_n215;
  tri   r800_n214;
  tri   r800_n213;
  tri   r800_n212;
  tri   r800_n211;
  tri   r800_n210;
  tri   r800_n209;
  tri   r800_n208;
  tri   r800_n207;
  tri   r800_n193;
  tri   r800_n206;
  tri   r800_n205;
  tri   r800_n204;
  tri   r800_n203;
  tri   r800_n202;
  tri   r800_n201;
  tri   r800_n200;
  tri   r800_n199;
  tri   r800_n198;
  tri   r800_n197;
  tri   r800_n183;
  tri   r800_n189;
  tri   r800_n196;
  tri   r800_n195;
  tri   r800_n190;
  tri   r800_n192;
  tri   r800_n194;
  tri   r800_n291;
  tri   r800_n290;
  tri   r800_n253;
  tri   r800_n259;
  tri   r800_n289;
  tri   r800_n288;
  tri   r800_n162;
  tri   r800_n287;
  tri   r800_n166;
  tri   r800_n286;
  tri   r800_n285;
  tri   r800_n284;
  tri   r800_n53;
  tri   r800_n56;
  tri   r800_n283;
  tri   r800_n282;
  tri   r800_n281;
  tri   r800_n46;
  tri   r800_n49;
  tri   r800_n280;
  tri   r800_n279;
  tri   r800_n278;
  tri   r800_n39;
  tri   r800_n42;
  tri   r800_n277;
  tri   r800_n276;
  tri   r800_n275;
  tri   r800_n32;
  tri   r800_n35;
  tri   r800_n274;
  tri   r800_n273;
  tri   r800_n272;
  tri   r800_n269;
  tri   r800_n271;
  tri   r800_n25;
  tri   r802_n55;
  tri   r802_n52;
  tri   r802_n51;
  tri   r802_n50;
  tri   r802_n48;
  tri   r802_n47;
  tri   r802_n45;
  tri   r802_n44;
  tri   r802_n43;
  tri   r802_n41;
  tri   r802_n40;
  tri   r802_n38;
  tri   r802_n37;
  tri   r802_n36;
  tri   r802_n34;
  tri   r802_n33;
  tri   r802_n31;
  tri   r802_n30;
  tri   r802_n29;
  tri   r802_n27;
  tri   r802_n26;
  tri   r802_n24;
  tri   r802_n23;
  tri   r802_n22;
  tri   r802_n20;
  tri   r802_n19;
  tri   r802_n17;
  tri   r802_n16;
  tri   r802_n15;
  tri   r802_n13;
  tri   r802_n12;
  tri   r802_n10;
  tri   r802_n9;
  tri   r802_n8;
  tri   r802_n6;
  tri   r802_n5;
  tri   r802_n3;
  tri   r802_n2;
  tri   r802_n1;
  tri   r802_n140;
  tri   r802_n139;
  tri   r802_n138;
  tri   r802_n137;
  tri   r802_n136;
  tri   r802_n134;
  tri   r802_n133;
  tri   r802_n132;
  tri   r802_n131;
  tri   r802_n130;
  tri   r802_n129;
  tri   r802_n128;
  tri   r802_n127;
  tri   r802_n126;
  tri   r802_n125;
  tri   r802_n124;
  tri   r802_n123;
  tri   r802_n122;
  tri   r802_n121;
  tri   r802_n120;
  tri   r802_n119;
  tri   r802_n118;
  tri   r802_n117;
  tri   r802_n116;
  tri   r802_n115;
  tri   r802_n114;
  tri   r802_n113;
  tri   r802_n112;
  tri   r802_n111;
  tri   r802_n110;
  tri   r802_n109;
  tri   r802_n108;
  tri   r802_n107;
  tri   r802_n106;
  tri   r802_n105;
  tri   r802_n104;
  tri   r802_n103;
  tri   r802_n102;
  tri   r802_n101;
  tri   r802_n100;
  tri   r802_n99;
  tri   r802_n98;
  tri   r802_n97;
  tri   r802_n96;
  tri   r802_n95;
  tri   r802_n94;
  tri   r802_n93;
  tri   r802_n92;
  tri   r802_n91;
  tri   r802_n90;
  tri   r802_n89;
  tri   r802_n88;
  tri   r802_n87;
  tri   r802_n86;
  tri   r802_n85;
  tri   r802_n84;
  tri   r802_n83;
  tri   r802_n82;
  tri   r802_n81;
  tri   r802_n80;
  tri   r802_n79;
  tri   r802_n78;
  tri   r802_n77;
  tri   r802_n76;
  tri   r802_n75;
  tri   r802_n74;
  tri   r802_n73;
  tri   r802_n72;
  tri   r802_n71;
  tri   r802_n70;
  tri   r802_n69;
  tri   r802_n67;
  tri   r802_n66;
  tri   r802_n65;
  tri   r802_n64;
  tri   r802_n63;
  tri   r802_n62;
  tri   r802_n61;
  tri   r802_n59;
  tri   r802_n60;
  tri   r802_n58;
  tri   r802_n57;
  tri   r802_n54;
  tri   r802_n228;
  tri   r802_n227;
  tri   r802_n226;
  tri   r802_n225;
  tri   r802_n222;
  tri   r802_n221;
  tri   r802_n220;
  tri   r802_n219;
  tri   r802_n218;
  tri   r802_n217;
  tri   r802_n216;
  tri   r802_n215;
  tri   r802_n214;
  tri   r802_n213;
  tri   r802_n212;
  tri   r802_n211;
  tri   r802_n210;
  tri   r802_n209;
  tri   r802_n208;
  tri   r802_n207;
  tri   r802_n206;
  tri   r802_n205;
  tri   r802_n204;
  tri   r802_n203;
  tri   r802_n202;
  tri   r802_n201;
  tri   r802_n200;
  tri   r802_n199;
  tri   r802_n198;
  tri   r802_n197;
  tri   r802_n196;
  tri   r802_n195;
  tri   r802_n194;
  tri   r802_n193;
  tri   r802_n192;
  tri   r802_n191;
  tri   r802_n190;
  tri   r802_n189;
  tri   r802_n188;
  tri   r802_n187;
  tri   r802_n186;
  tri   r802_n185;
  tri   r802_n184;
  tri   r802_n183;
  tri   r802_n182;
  tri   r802_n181;
  tri   r802_n180;
  tri   r802_n179;
  tri   r802_n178;
  tri   r802_n177;
  tri   r802_n176;
  tri   r802_n175;
  tri   r802_n174;
  tri   r802_n173;
  tri   r802_n172;
  tri   r802_n171;
  tri   r802_n170;
  tri   r802_n169;
  tri   r802_n168;
  tri   r802_n167;
  tri   r802_n164;
  tri   r802_n163;
  tri   r802_n161;
  tri   r802_n160;
  tri   r802_n159;
  tri   r802_n158;
  tri   r802_n157;
  tri   r802_n156;
  tri   r802_n155;
  tri   r802_n154;
  tri   r802_n153;
  tri   r802_n152;
  tri   r802_n151;
  tri   r802_n150;
  tri   r802_n149;
  tri   r802_n135;
  tri   r802_n141;
  tri   r802_n148;
  tri   r802_n147;
  tri   r802_n142;
  tri   r802_n146;
  tri   r802_n143;
  tri   r802_n145;
  tri   r802_n144;
  tri   r802_n291;
  tri   r802_n290;
  tri   r802_n289;
  tri   r802_n288;
  tri   r802_n162;
  tri   r802_n287;
  tri   r802_n166;
  tri   r802_n286;
  tri   r802_n285;
  tri   r802_n284;
  tri   r802_n53;
  tri   r802_n56;
  tri   r802_n283;
  tri   r802_n282;
  tri   r802_n281;
  tri   r802_n46;
  tri   r802_n49;
  tri   r802_n280;
  tri   r802_n279;
  tri   r802_n278;
  tri   r802_n39;
  tri   r802_n42;
  tri   r802_n277;
  tri   r802_n276;
  tri   r802_n275;
  tri   r802_n32;
  tri   r802_n35;
  tri   r802_n274;
  tri   r802_n273;
  tri   r802_n272;
  tri   r802_n25;
  tri   r802_n28;
  tri   r802_n271;
  tri   r802_n270;
  tri   r802_n269;
  tri   r802_n18;
  tri   r802_n21;
  tri   r802_n268;
  tri   r802_n267;
  tri   r802_n266;
  tri   r802_n11;
  tri   r802_n14;
  tri   r802_n265;
  tri   r802_n264;
  tri   r802_n263;
  tri   r802_n4;
  tri   r802_n7;
  tri   r802_n262;
  tri   r802_n261;
  tri   r802_n260;
  tri   r802_n259;
  tri   r802_n258;
  tri   r802_n257;
  tri   r802_n256;
  tri   r802_n255;
  tri   r802_n254;
  tri   r802_n253;
  tri   r802_n252;
  tri   r802_n251;
  tri   r802_n250;
  tri   r802_n249;
  tri   r802_n248;
  tri   r802_n247;
  tri   r802_n246;
  tri   r802_n245;
  tri   r802_n244;
  tri   r802_n243;
  tri   r802_n242;
  tri   r802_n241;
  tri   r802_n240;
  tri   r802_n239;
  tri   r802_n238;
  tri   r802_n237;
  tri   r802_n223;
  tri   r802_n229;
  tri   r802_n236;
  tri   r802_n235;
  tri   r802_n234;
  tri   r802_n233;
  tri   r802_n232;
  tri   r802_n224;
  tri   r802_n231;
  tri   r802_n230;
  tri   r804_n86;
  tri   r804_n85;
  tri   r804_n82;
  tri   r804_n81;
  tri   r804_n80;
  tri   r804_n79;
  tri   r804_n78;
  tri   r804_n77;
  tri   r804_n76;
  tri   r804_n75;
  tri   r804_n74;
  tri   r804_n72;
  tri   r804_n71;
  tri   r804_n70;
  tri   r804_n69;
  tri   r804_n68;
  tri   r804_n66;
  tri   r804_n65;
  tri   r804_n64;
  tri   r804_n63;
  tri   r804_n62;
  tri   r804_n61;
  tri   r804_n60;
  tri   r804_n59;
  tri   r804_n58;
  tri   r804_n57;
  tri   r804_n55;
  tri   r804_n54;
  tri   r804_n53;
  tri   r804_n51;
  tri   r804_n50;
  tri   r804_n48;
  tri   r804_n47;
  tri   r804_n46;
  tri   r804_n44;
  tri   r804_n43;
  tri   r804_n41;
  tri   r804_n40;
  tri   r804_n39;
  tri   r804_n37;
  tri   r804_n36;
  tri   r804_n34;
  tri   r804_n33;
  tri   r804_n32;
  tri   r804_n30;
  tri   r804_n29;
  tri   r804_n27;
  tri   r804_n26;
  tri   r804_n25;
  tri   r804_n23;
  tri   r804_n22;
  tri   r804_n20;
  tri   r804_n19;
  tri   r804_n18;
  tri   r804_n16;
  tri   r804_n15;
  tri   r804_n13;
  tri   r804_n12;
  tri   r804_n11;
  tri   r804_n9;
  tri   r804_n8;
  tri   r804_n6;
  tri   r804_n5;
  tri   r804_n4;
  tri   r804_n2;
  tri   r804_n1;
  tri   r804_n172;
  tri   r804_n169;
  tri   r804_n168;
  tri   r804_n167;
  tri   r804_n166;
  tri   r804_n165;
  tri   r804_n163;
  tri   r804_n162;
  tri   r804_n160;
  tri   r804_n159;
  tri   r804_n158;
  tri   r804_n157;
  tri   r804_n156;
  tri   r804_n155;
  tri   r804_n154;
  tri   r804_n152;
  tri   r804_n151;
  tri   r804_n150;
  tri   r804_n149;
  tri   r804_n148;
  tri   r804_n147;
  tri   r804_n146;
  tri   r804_n145;
  tri   r804_n144;
  tri   r804_n142;
  tri   r804_n141;
  tri   r804_n140;
  tri   r804_n139;
  tri   r804_n138;
  tri   r804_n137;
  tri   r804_n136;
  tri   r804_n135;
  tri   r804_n134;
  tri   r804_n132;
  tri   r804_n131;
  tri   r804_n130;
  tri   r804_n129;
  tri   r804_n128;
  tri   r804_n127;
  tri   r804_n126;
  tri   r804_n125;
  tri   r804_n124;
  tri   r804_n122;
  tri   r804_n121;
  tri   r804_n120;
  tri   r804_n119;
  tri   r804_n118;
  tri   r804_n117;
  tri   r804_n116;
  tri   r804_n115;
  tri   r804_n114;
  tri   r804_n112;
  tri   r804_n111;
  tri   r804_n110;
  tri   r804_n109;
  tri   r804_n108;
  tri   r804_n107;
  tri   r804_n106;
  tri   r804_n105;
  tri   r804_n104;
  tri   r804_n102;
  tri   r804_n101;
  tri   r804_n100;
  tri   r804_n99;
  tri   r804_n98;
  tri   r804_n97;
  tri   r804_n96;
  tri   r804_n95;
  tri   r804_n94;
  tri   r804_n92;
  tri   r804_n91;
  tri   r804_n90;
  tri   r804_n89;
  tri   r804_n88;
  tri   r804_n84;
  tri   r804_n87;
  tri   r804_n256;
  tri   r804_n255;
  tri   r804_n253;
  tri   r804_n252;
  tri   r804_n251;
  tri   r804_n249;
  tri   r804_n248;
  tri   r804_n247;
  tri   r804_n246;
  tri   r804_n245;
  tri   r804_n244;
  tri   r804_n243;
  tri   r804_n242;
  tri   r804_n241;
  tri   r804_n239;
  tri   r804_n238;
  tri   r804_n237;
  tri   r804_n236;
  tri   r804_n235;
  tri   r804_n234;
  tri   r804_n233;
  tri   r804_n232;
  tri   r804_n231;
  tri   r804_n229;
  tri   r804_n228;
  tri   r804_n227;
  tri   r804_n226;
  tri   r804_n225;
  tri   r804_n224;
  tri   r804_n223;
  tri   r804_n222;
  tri   r804_n221;
  tri   r804_n219;
  tri   r804_n218;
  tri   r804_n217;
  tri   r804_n216;
  tri   r804_n215;
  tri   r804_n214;
  tri   r804_n213;
  tri   r804_n212;
  tri   r804_n211;
  tri   r804_n209;
  tri   r804_n208;
  tri   r804_n207;
  tri   r804_n206;
  tri   r804_n205;
  tri   r804_n204;
  tri   r804_n203;
  tri   r804_n202;
  tri   r804_n201;
  tri   r804_n199;
  tri   r804_n198;
  tri   r804_n197;
  tri   r804_n196;
  tri   r804_n195;
  tri   r804_n194;
  tri   r804_n193;
  tri   r804_n192;
  tri   r804_n191;
  tri   r804_n189;
  tri   r804_n188;
  tri   r804_n187;
  tri   r804_n186;
  tri   r804_n185;
  tri   r804_n184;
  tri   r804_n183;
  tri   r804_n182;
  tri   r804_n181;
  tri   r804_n179;
  tri   r804_n178;
  tri   r804_n177;
  tri   r804_n176;
  tri   r804_n175;
  tri   r804_n171;
  tri   r804_n173;
  tri   r804_n174;
  tri   r804_n289;
  tri   r804_n288;
  tri   r804_n161;
  tri   r804_n287;
  tri   r804_n286;
  tri   r804_n285;
  tri   r804_n52;
  tri   r804_n284;
  tri   r804_n283;
  tri   r804_n282;
  tri   r804_n45;
  tri   r804_n281;
  tri   r804_n280;
  tri   r804_n279;
  tri   r804_n38;
  tri   r804_n278;
  tri   r804_n277;
  tri   r804_n276;
  tri   r804_n31;
  tri   r804_n275;
  tri   r804_n274;
  tri   r804_n273;
  tri   r804_n24;
  tri   r804_n272;
  tri   r804_n271;
  tri   r804_n270;
  tri   r804_n17;
  tri   r804_n269;
  tri   r804_n268;
  tri   r804_n267;
  tri   r804_n10;
  tri   r804_n266;
  tri   r804_n265;
  tri   r804_n264;
  tri   r804_n3;
  tri   r804_n263;
  tri   r804_n254;
  tri   r804_n262;
  tri   r804_n261;
  tri   r804_n257;
  tri   r804_n259;
  tri   r804_n258;
  tri   r806_n41;
  tri   r806_n40;
  tri   r806_n38;
  tri   r806_n37;
  tri   r806_n36;
  tri   r806_n34;
  tri   r806_n33;
  tri   r806_n31;
  tri   r806_n30;
  tri   r806_n29;
  tri   r806_n27;
  tri   r806_n26;
  tri   r806_n24;
  tri   r806_n23;
  tri   r806_n22;
  tri   r806_n20;
  tri   r806_n19;
  tri   r806_n17;
  tri   r806_n16;
  tri   r806_n15;
  tri   r806_n13;
  tri   r806_n12;
  tri   r806_n10;
  tri   r806_n9;
  tri   r806_n8;
  tri   r806_n6;
  tri   r806_n5;
  tri   r806_n3;
  tri   r806_n2;
  tri   r806_n1;
  tri   r806_n133;
  tri   r806_n130;
  tri   r806_n129;
  tri   r806_n128;
  tri   r806_n127;
  tri   r806_n126;
  tri   r806_n124;
  tri   r806_n123;
  tri   r806_n122;
  tri   r806_n121;
  tri   r806_n120;
  tri   r806_n119;
  tri   r806_n118;
  tri   r806_n117;
  tri   r806_n116;
  tri   r806_n115;
  tri   r806_n114;
  tri   r806_n113;
  tri   r806_n112;
  tri   r806_n111;
  tri   r806_n110;
  tri   r806_n109;
  tri   r806_n108;
  tri   r806_n107;
  tri   r806_n106;
  tri   r806_n105;
  tri   r806_n104;
  tri   r806_n103;
  tri   r806_n102;
  tri   r806_n101;
  tri   r806_n100;
  tri   r806_n99;
  tri   r806_n98;
  tri   r806_n97;
  tri   r806_n96;
  tri   r806_n95;
  tri   r806_n94;
  tri   r806_n93;
  tri   r806_n92;
  tri   r806_n91;
  tri   r806_n90;
  tri   r806_n89;
  tri   r806_n88;
  tri   r806_n87;
  tri   r806_n86;
  tri   r806_n85;
  tri   r806_n84;
  tri   r806_n83;
  tri   r806_n82;
  tri   r806_n81;
  tri   r806_n80;
  tri   r806_n79;
  tri   r806_n78;
  tri   r806_n77;
  tri   r806_n76;
  tri   r806_n75;
  tri   r806_n74;
  tri   r806_n73;
  tri   r806_n72;
  tri   r806_n71;
  tri   r806_n70;
  tri   r806_n69;
  tri   r806_n67;
  tri   r806_n66;
  tri   r806_n65;
  tri   r806_n64;
  tri   r806_n63;
  tri   r806_n62;
  tri   r806_n61;
  tri   r806_n59;
  tri   r806_n60;
  tri   r806_n58;
  tri   r806_n57;
  tri   r806_n55;
  tri   r806_n54;
  tri   r806_n52;
  tri   r806_n51;
  tri   r806_n50;
  tri   r806_n48;
  tri   r806_n47;
  tri   r806_n43;
  tri   r806_n44;
  tri   r806_n45;
  tri   r806_n218;
  tri   r806_n217;
  tri   r806_n216;
  tri   r806_n215;
  tri   r806_n214;
  tri   r806_n212;
  tri   r806_n211;
  tri   r806_n210;
  tri   r806_n209;
  tri   r806_n208;
  tri   r806_n207;
  tri   r806_n206;
  tri   r806_n205;
  tri   r806_n204;
  tri   r806_n203;
  tri   r806_n202;
  tri   r806_n201;
  tri   r806_n200;
  tri   r806_n199;
  tri   r806_n198;
  tri   r806_n197;
  tri   r806_n196;
  tri   r806_n195;
  tri   r806_n194;
  tri   r806_n193;
  tri   r806_n192;
  tri   r806_n191;
  tri   r806_n190;
  tri   r806_n189;
  tri   r806_n188;
  tri   r806_n187;
  tri   r806_n186;
  tri   r806_n185;
  tri   r806_n184;
  tri   r806_n183;
  tri   r806_n182;
  tri   r806_n181;
  tri   r806_n180;
  tri   r806_n179;
  tri   r806_n178;
  tri   r806_n177;
  tri   r806_n176;
  tri   r806_n175;
  tri   r806_n174;
  tri   r806_n173;
  tri   r806_n172;
  tri   r806_n171;
  tri   r806_n170;
  tri   r806_n169;
  tri   r806_n168;
  tri   r806_n167;
  tri   r806_n164;
  tri   r806_n163;
  tri   r806_n161;
  tri   r806_n160;
  tri   r806_n159;
  tri   r806_n158;
  tri   r806_n157;
  tri   r806_n156;
  tri   r806_n155;
  tri   r806_n154;
  tri   r806_n153;
  tri   r806_n152;
  tri   r806_n151;
  tri   r806_n150;
  tri   r806_n149;
  tri   r806_n135;
  tri   r806_n148;
  tri   r806_n147;
  tri   r806_n146;
  tri   r806_n145;
  tri   r806_n144;
  tri   r806_n143;
  tri   r806_n142;
  tri   r806_n141;
  tri   r806_n140;
  tri   r806_n139;
  tri   r806_n125;
  tri   r806_n131;
  tri   r806_n138;
  tri   r806_n137;
  tri   r806_n132;
  tri   r806_n134;
  tri   r806_n136;
  tri   r806_n289;
  tri   r806_n288;
  tri   r806_n166;
  tri   r806_n286;
  tri   r806_n285;
  tri   r806_n284;
  tri   r806_n53;
  tri   r806_n56;
  tri   r806_n283;
  tri   r806_n282;
  tri   r806_n281;
  tri   r806_n46;
  tri   r806_n49;
  tri   r806_n280;
  tri   r806_n279;
  tri   r806_n278;
  tri   r806_n39;
  tri   r806_n42;
  tri   r806_n277;
  tri   r806_n276;
  tri   r806_n275;
  tri   r806_n32;
  tri   r806_n35;
  tri   r806_n274;
  tri   r806_n273;
  tri   r806_n272;
  tri   r806_n25;
  tri   r806_n28;
  tri   r806_n271;
  tri   r806_n270;
  tri   r806_n269;
  tri   r806_n18;
  tri   r806_n21;
  tri   r806_n268;
  tri   r806_n267;
  tri   r806_n266;
  tri   r806_n11;
  tri   r806_n14;
  tri   r806_n265;
  tri   r806_n264;
  tri   r806_n263;
  tri   r806_n4;
  tri   r806_n7;
  tri   r806_n262;
  tri   r806_n261;
  tri   r806_n260;
  tri   r806_n259;
  tri   r806_n258;
  tri   r806_n257;
  tri   r806_n256;
  tri   r806_n255;
  tri   r806_n254;
  tri   r806_n253;
  tri   r806_n252;
  tri   r806_n251;
  tri   r806_n250;
  tri   r806_n249;
  tri   r806_n248;
  tri   r806_n247;
  tri   r806_n246;
  tri   r806_n245;
  tri   r806_n244;
  tri   r806_n243;
  tri   r806_n242;
  tri   r806_n241;
  tri   r806_n240;
  tri   r806_n239;
  tri   r806_n238;
  tri   r806_n237;
  tri   r806_n236;
  tri   r806_n235;
  tri   r806_n234;
  tri   r806_n233;
  tri   r806_n232;
  tri   r806_n231;
  tri   r806_n230;
  tri   r806_n229;
  tri   r806_n228;
  tri   r806_n227;
  tri   r806_n213;
  tri   r806_n219;
  tri   r806_n226;
  tri   r806_n225;
  tri   r806_n220;
  tri   r806_n224;
  tri   r806_n221;
  tri   r806_n223;
  tri   r806_n222;
  tri   r806_n287;
  tri   r806_n291;
  tri   r806_n290;
  tri   r806_n162;
  tri   r808_n76;
  tri   r808_n75;
  tri   r808_n74;
  tri   r808_n72;
  tri   r808_n71;
  tri   r808_n70;
  tri   r808_n69;
  tri   r808_n68;
  tri   r808_n66;
  tri   r808_n65;
  tri   r808_n64;
  tri   r808_n63;
  tri   r808_n62;
  tri   r808_n61;
  tri   r808_n60;
  tri   r808_n59;
  tri   r808_n58;
  tri   r808_n57;
  tri   r808_n55;
  tri   r808_n54;
  tri   r808_n53;
  tri   r808_n51;
  tri   r808_n50;
  tri   r808_n48;
  tri   r808_n47;
  tri   r808_n46;
  tri   r808_n44;
  tri   r808_n43;
  tri   r808_n41;
  tri   r808_n40;
  tri   r808_n39;
  tri   r808_n37;
  tri   r808_n36;
  tri   r808_n34;
  tri   r808_n33;
  tri   r808_n32;
  tri   r808_n30;
  tri   r808_n29;
  tri   r808_n27;
  tri   r808_n26;
  tri   r808_n25;
  tri   r808_n23;
  tri   r808_n22;
  tri   r808_n20;
  tri   r808_n19;
  tri   r808_n18;
  tri   r808_n16;
  tri   r808_n15;
  tri   r808_n13;
  tri   r808_n12;
  tri   r808_n11;
  tri   r808_n9;
  tri   r808_n8;
  tri   r808_n6;
  tri   r808_n5;
  tri   r808_n4;
  tri   r808_n2;
  tri   r808_n1;
  tri   r808_n163;
  tri   r808_n160;
  tri   r808_n159;
  tri   r808_n158;
  tri   r808_n156;
  tri   r808_n155;
  tri   r808_n154;
  tri   r808_n152;
  tri   r808_n151;
  tri   r808_n150;
  tri   r808_n149;
  tri   r808_n148;
  tri   r808_n147;
  tri   r808_n146;
  tri   r808_n145;
  tri   r808_n144;
  tri   r808_n142;
  tri   r808_n141;
  tri   r808_n140;
  tri   r808_n139;
  tri   r808_n138;
  tri   r808_n137;
  tri   r808_n136;
  tri   r808_n135;
  tri   r808_n134;
  tri   r808_n132;
  tri   r808_n131;
  tri   r808_n130;
  tri   r808_n129;
  tri   r808_n128;
  tri   r808_n127;
  tri   r808_n126;
  tri   r808_n125;
  tri   r808_n124;
  tri   r808_n122;
  tri   r808_n121;
  tri   r808_n120;
  tri   r808_n119;
  tri   r808_n118;
  tri   r808_n117;
  tri   r808_n116;
  tri   r808_n115;
  tri   r808_n114;
  tri   r808_n112;
  tri   r808_n111;
  tri   r808_n110;
  tri   r808_n109;
  tri   r808_n108;
  tri   r808_n107;
  tri   r808_n106;
  tri   r808_n105;
  tri   r808_n104;
  tri   r808_n102;
  tri   r808_n101;
  tri   r808_n100;
  tri   r808_n99;
  tri   r808_n98;
  tri   r808_n97;
  tri   r808_n96;
  tri   r808_n95;
  tri   r808_n94;
  tri   r808_n92;
  tri   r808_n91;
  tri   r808_n90;
  tri   r808_n89;
  tri   r808_n88;
  tri   r808_n87;
  tri   r808_n86;
  tri   r808_n85;
  tri   r808_n84;
  tri   r808_n82;
  tri   r808_n81;
  tri   r808_n80;
  tri   r808_n77;
  tri   r808_n79;
  tri   r808_n78;
  tri   r808_n247;
  tri   r808_n246;
  tri   r808_n245;
  tri   r808_n243;
  tri   r808_n242;
  tri   r808_n241;
  tri   r808_n239;
  tri   r808_n238;
  tri   r808_n237;
  tri   r808_n236;
  tri   r808_n235;
  tri   r808_n234;
  tri   r808_n233;
  tri   r808_n232;
  tri   r808_n231;
  tri   r808_n229;
  tri   r808_n228;
  tri   r808_n227;
  tri   r808_n226;
  tri   r808_n225;
  tri   r808_n224;
  tri   r808_n223;
  tri   r808_n222;
  tri   r808_n221;
  tri   r808_n219;
  tri   r808_n218;
  tri   r808_n217;
  tri   r808_n216;
  tri   r808_n215;
  tri   r808_n214;
  tri   r808_n213;
  tri   r808_n212;
  tri   r808_n211;
  tri   r808_n209;
  tri   r808_n208;
  tri   r808_n207;
  tri   r808_n206;
  tri   r808_n205;
  tri   r808_n204;
  tri   r808_n203;
  tri   r808_n202;
  tri   r808_n201;
  tri   r808_n199;
  tri   r808_n198;
  tri   r808_n197;
  tri   r808_n196;
  tri   r808_n195;
  tri   r808_n194;
  tri   r808_n193;
  tri   r808_n192;
  tri   r808_n191;
  tri   r808_n189;
  tri   r808_n188;
  tri   r808_n187;
  tri   r808_n186;
  tri   r808_n185;
  tri   r808_n184;
  tri   r808_n183;
  tri   r808_n182;
  tri   r808_n181;
  tri   r808_n179;
  tri   r808_n178;
  tri   r808_n177;
  tri   r808_n176;
  tri   r808_n175;
  tri   r808_n174;
  tri   r808_n173;
  tri   r808_n172;
  tri   r808_n171;
  tri   r808_n169;
  tri   r808_n168;
  tri   r808_n167;
  tri   r808_n157;
  tri   r808_n166;
  tri   r808_n165;
  tri   r808_n162;
  tri   r808_n289;
  tri   r808_n288;
  tri   r808_n161;
  tri   r808_n287;
  tri   r808_n286;
  tri   r808_n285;
  tri   r808_n52;
  tri   r808_n284;
  tri   r808_n283;
  tri   r808_n282;
  tri   r808_n45;
  tri   r808_n281;
  tri   r808_n280;
  tri   r808_n279;
  tri   r808_n38;
  tri   r808_n278;
  tri   r808_n277;
  tri   r808_n276;
  tri   r808_n31;
  tri   r808_n275;
  tri   r808_n274;
  tri   r808_n273;
  tri   r808_n24;
  tri   r808_n272;
  tri   r808_n271;
  tri   r808_n270;
  tri   r808_n17;
  tri   r808_n269;
  tri   r808_n268;
  tri   r808_n267;
  tri   r808_n10;
  tri   r808_n266;
  tri   r808_n265;
  tri   r808_n264;
  tri   r808_n3;
  tri   r808_n263;
  tri   r808_n262;
  tri   r808_n261;
  tri   r808_n259;
  tri   r808_n258;
  tri   r808_n257;
  tri   r808_n256;
  tri   r808_n255;
  tri   r808_n254;
  tri   r808_n253;
  tri   r808_n244;
  tri   r808_n252;
  tri   r808_n251;
  tri   r808_n248;
  tri   r808_n249;
  tri   r810_n30;
  tri   r810_n29;
  tri   r810_n27;
  tri   r810_n26;
  tri   r810_n24;
  tri   r810_n23;
  tri   r810_n22;
  tri   r810_n20;
  tri   r810_n19;
  tri   r810_n17;
  tri   r810_n16;
  tri   r810_n15;
  tri   r810_n13;
  tri   r810_n12;
  tri   r810_n10;
  tri   r810_n9;
  tri   r810_n8;
  tri   r810_n6;
  tri   r810_n5;
  tri   r810_n3;
  tri   r810_n2;
  tri   r810_n1;
  tri   r810_n124;
  tri   r810_n123;
  tri   r810_n120;
  tri   r810_n119;
  tri   r810_n118;
  tri   r810_n117;
  tri   r810_n116;
  tri   r810_n114;
  tri   r810_n113;
  tri   r810_n112;
  tri   r810_n111;
  tri   r810_n110;
  tri   r810_n109;
  tri   r810_n108;
  tri   r810_n107;
  tri   r810_n106;
  tri   r810_n105;
  tri   r810_n104;
  tri   r810_n103;
  tri   r810_n102;
  tri   r810_n101;
  tri   r810_n100;
  tri   r810_n99;
  tri   r810_n98;
  tri   r810_n97;
  tri   r810_n96;
  tri   r810_n95;
  tri   r810_n94;
  tri   r810_n93;
  tri   r810_n92;
  tri   r810_n91;
  tri   r810_n90;
  tri   r810_n89;
  tri   r810_n88;
  tri   r810_n87;
  tri   r810_n86;
  tri   r810_n85;
  tri   r810_n84;
  tri   r810_n83;
  tri   r810_n82;
  tri   r810_n81;
  tri   r810_n80;
  tri   r810_n79;
  tri   r810_n78;
  tri   r810_n77;
  tri   r810_n76;
  tri   r810_n75;
  tri   r810_n74;
  tri   r810_n73;
  tri   r810_n72;
  tri   r810_n71;
  tri   r810_n70;
  tri   r810_n69;
  tri   r810_n67;
  tri   r810_n66;
  tri   r810_n65;
  tri   r810_n64;
  tri   r810_n63;
  tri   r810_n62;
  tri   r810_n61;
  tri   r810_n59;
  tri   r810_n60;
  tri   r810_n58;
  tri   r810_n57;
  tri   r810_n55;
  tri   r810_n54;
  tri   r810_n52;
  tri   r810_n51;
  tri   r810_n50;
  tri   r810_n48;
  tri   r810_n47;
  tri   r810_n45;
  tri   r810_n44;
  tri   r810_n43;
  tri   r810_n41;
  tri   r810_n40;
  tri   r810_n38;
  tri   r810_n37;
  tri   r810_n36;
  tri   r810_n31;
  tri   r810_n34;
  tri   r810_n33;
  tri   r810_n211;
  tri   r810_n208;
  tri   r810_n207;
  tri   r810_n206;
  tri   r810_n205;
  tri   r810_n204;
  tri   r810_n202;
  tri   r810_n201;
  tri   r810_n200;
  tri   r810_n199;
  tri   r810_n198;
  tri   r810_n197;
  tri   r810_n196;
  tri   r810_n195;
  tri   r810_n194;
  tri   r810_n193;
  tri   r810_n192;
  tri   r810_n191;
  tri   r810_n190;
  tri   r810_n189;
  tri   r810_n188;
  tri   r810_n187;
  tri   r810_n186;
  tri   r810_n185;
  tri   r810_n184;
  tri   r810_n183;
  tri   r810_n182;
  tri   r810_n181;
  tri   r810_n180;
  tri   r810_n179;
  tri   r810_n178;
  tri   r810_n177;
  tri   r810_n176;
  tri   r810_n175;
  tri   r810_n174;
  tri   r810_n173;
  tri   r810_n172;
  tri   r810_n171;
  tri   r810_n170;
  tri   r810_n169;
  tri   r810_n168;
  tri   r810_n167;
  tri   r810_n164;
  tri   r810_n163;
  tri   r810_n161;
  tri   r810_n160;
  tri   r810_n159;
  tri   r810_n158;
  tri   r810_n157;
  tri   r810_n156;
  tri   r810_n155;
  tri   r810_n154;
  tri   r810_n153;
  tri   r810_n152;
  tri   r810_n151;
  tri   r810_n150;
  tri   r810_n149;
  tri   r810_n148;
  tri   r810_n147;
  tri   r810_n146;
  tri   r810_n145;
  tri   r810_n144;
  tri   r810_n143;
  tri   r810_n142;
  tri   r810_n141;
  tri   r810_n140;
  tri   r810_n139;
  tri   r810_n125;
  tri   r810_n138;
  tri   r810_n137;
  tri   r810_n136;
  tri   r810_n135;
  tri   r810_n134;
  tri   r810_n133;
  tri   r810_n132;
  tri   r810_n131;
  tri   r810_n130;
  tri   r810_n129;
  tri   r810_n115;
  tri   r810_n121;
  tri   r810_n128;
  tri   r810_n127;
  tri   r810_n122;
  tri   r810_n126;
  tri   r810_n56;
  tri   r810_n283;
  tri   r810_n282;
  tri   r810_n281;
  tri   r810_n46;
  tri   r810_n49;
  tri   r810_n280;
  tri   r810_n279;
  tri   r810_n278;
  tri   r810_n39;
  tri   r810_n42;
  tri   r810_n277;
  tri   r810_n276;
  tri   r810_n275;
  tri   r810_n32;
  tri   r810_n35;
  tri   r810_n274;
  tri   r810_n273;
  tri   r810_n272;
  tri   r810_n25;
  tri   r810_n28;
  tri   r810_n271;
  tri   r810_n270;
  tri   r810_n269;
  tri   r810_n18;
  tri   r810_n21;
  tri   r810_n268;
  tri   r810_n267;
  tri   r810_n266;
  tri   r810_n11;
  tri   r810_n14;
  tri   r810_n265;
  tri   r810_n264;
  tri   r810_n263;
  tri   r810_n4;
  tri   r810_n7;
  tri   r810_n262;
  tri   r810_n261;
  tri   r810_n260;
  tri   r810_n258;
  tri   r810_n257;
  tri   r810_n256;
  tri   r810_n255;
  tri   r810_n254;
  tri   r810_n252;
  tri   r810_n251;
  tri   r810_n250;
  tri   r810_n249;
  tri   r810_n248;
  tri   r810_n247;
  tri   r810_n246;
  tri   r810_n245;
  tri   r810_n244;
  tri   r810_n243;
  tri   r810_n242;
  tri   r810_n241;
  tri   r810_n240;
  tri   r810_n239;
  tri   r810_n238;
  tri   r810_n237;
  tri   r810_n236;
  tri   r810_n235;
  tri   r810_n234;
  tri   r810_n233;
  tri   r810_n232;
  tri   r810_n231;
  tri   r810_n230;
  tri   r810_n229;
  tri   r810_n228;
  tri   r810_n227;
  tri   r810_n213;
  tri   r810_n226;
  tri   r810_n225;
  tri   r810_n224;
  tri   r810_n223;
  tri   r810_n222;
  tri   r810_n221;
  tri   r810_n220;
  tri   r810_n219;
  tri   r810_n218;
  tri   r810_n217;
  tri   r810_n203;
  tri   r810_n209;
  tri   r810_n216;
  tri   r810_n215;
  tri   r810_n210;
  tri   r810_n212;
  tri   r810_n214;
  tri   r810_n291;
  tri   r810_n290;
  tri   r810_n253;
  tri   r810_n259;
  tri   r810_n289;
  tri   r810_n288;
  tri   r810_n162;
  tri   r810_n287;
  tri   r810_n166;
  tri   r810_n286;
  tri   r810_n53;
  tri   r810_n285;
  tri   r810_n284;
  tri   r812_n78;
  tri   r812_n77;
  tri   r812_n76;
  tri   r812_n73;
  tri   r812_n72;
  tri   r812_n71;
  tri   r812_n70;
  tri   r812_n69;
  tri   r812_n68;
  tri   r812_n66;
  tri   r812_n65;
  tri   r812_n64;
  tri   r812_n63;
  tri   r812_n62;
  tri   r812_n61;
  tri   r812_n60;
  tri   r812_n58;
  tri   r812_n57;
  tri   r812_n56;
  tri   r812_n55;
  tri   r812_n54;
  tri   r812_n53;
  tri   r812_n52;
  tri   r812_n50;
  tri   r812_n49;
  tri   r812_n48;
  tri   r812_n47;
  tri   r812_n46;
  tri   r812_n45;
  tri   r812_n44;
  tri   r812_n42;
  tri   r812_n41;
  tri   r812_n40;
  tri   r812_n39;
  tri   r812_n38;
  tri   r812_n37;
  tri   r812_n36;
  tri   r812_n35;
  tri   r812_n34;
  tri   r812_n32;
  tri   r812_n31;
  tri   r812_n29;
  tri   r812_n28;
  tri   r812_n27;
  tri   r812_n24;
  tri   r812_n23;
  tri   r812_n22;
  tri   r812_n21;
  tri   r812_n20;
  tri   r812_n17;
  tri   r812_n16;
  tri   r812_n15;
  tri   r812_n14;
  tri   r812_n13;
  tri   r812_n10;
  tri   r812_n9;
  tri   r812_n8;
  tri   r812_n7;
  tri   r812_n6;
  tri   r812_n3;
  tri   r812_n2;
  tri   r812_n1;
  tri   r812_n124;
  tri   r812_n123;
  tri   r812_n121;
  tri   r812_n120;
  tri   r812_n26;
  tri   r812_n119;
  tri   r812_n19;
  tri   r812_n118;
  tri   r812_n12;
  tri   r812_n117;
  tri   r812_n5;
  tri   r812_n116;
  tri   r812_n115;
  tri   r812_n114;
  tri   r812_n113;
  tri   r812_n112;
  tri   r812_n111;
  tri   r812_n109;
  tri   r812_n108;
  tri   r812_n107;
  tri   r812_n106;
  tri   r812_n105;
  tri   r812_n104;
  tri   r812_n103;
  tri   r812_n101;
  tri   r812_n100;
  tri   r812_n99;
  tri   r812_n98;
  tri   r812_n97;
  tri   r812_n96;
  tri   r812_n95;
  tri   r812_n93;
  tri   r812_n92;
  tri   r812_n91;
  tri   r812_n90;
  tri   r812_n89;
  tri   r812_n88;
  tri   r812_n87;
  tri   r812_n85;
  tri   r812_n84;
  tri   r812_n83;
  tri   r812_n82;
  tri   r812_n74;
  tri   r812_n79;
  tri   r812_n80;
  tri   r812_n81;
  tri   r812_n18;
  tri   r812_n33;
  tri   r812_n125;
  tri   r812_n128;
  tri   r812_n131;
  tri   r812_n135;
  tri   r812_n138;
  tri   r812_n141;
  tri   r816_n138;
  tri   r816_n136;
  tri   r816_n135;
  tri   r816_n119;
  tri   r816_n118;
  tri   r816_n117;
  tri   r816_n115;
  tri   r816_n114;
  tri   r816_n112;
  tri   r816_n111;
  tri   r816_n110;
  tri   r816_n108;
  tri   r816_n107;
  tri   r816_n103;
  tri   r816_n102;
  tri   r816_n101;
  tri   r816_n100;
  tri   r816_n97;
  tri   r816_n96;
  tri   r816_n95;
  tri   r816_n93;
  tri   r816_n92;
  tri   r816_n88;
  tri   r816_n87;
  tri   r816_n86;
  tri   r816_n85;
  tri   r816_n82;
  tri   r816_n81;
  tri   r816_n80;
  tri   r816_n78;
  tri   r816_n77;
  tri   r816_n73;
  tri   r816_n72;
  tri   r816_n71;
  tri   r816_n70;
  tri   r816_n67;
  tri   r816_n66;
  tri   r816_n65;
  tri   r816_n63;
  tri   r816_n62;
  tri   r816_n58;
  tri   r816_n57;
  tri   r816_n56;
  tri   r816_n55;
  tri   r816_n52;
  tri   r816_n51;
  tri   r816_n50;
  tri   r816_n48;
  tri   r816_n47;
  tri   r816_n43;
  tri   r816_n42;
  tri   r816_n41;
  tri   r816_n40;
  tri   r816_n37;
  tri   r816_n36;
  tri   r816_n35;
  tri   r816_n33;
  tri   r816_n32;
  tri   r816_n28;
  tri   r816_n27;
  tri   r816_n26;
  tri   r816_n25;
  tri   r816_n22;
  tri   r816_n21;
  tri   r816_n20;
  tri   r816_n18;
  tri   r816_n17;
  tri   r816_n13;
  tri   r816_n12;
  tri   r816_n11;
  tri   r816_n10;
  tri   r816_n7;
  tri   r816_n5;
  tri   r816_n3;
  tri   r816_n2;
  tri   r816_n1;
  tri   r816_n216;
  tri   r816_n83;
  tri   r816_n214;
  tri   r816_n213;
  tri   r816_n212;
  tri   r816_n210;
  tri   r816_n74;
  tri   r816_n76;
  tri   r816_n208;
  tri   r816_n207;
  tri   r816_n206;
  tri   r816_n205;
  tri   r816_n204;
  tri   r816_n203;
  tri   r816_n201;
  tri   r816_n127;
  tri   r816_n68;
  tri   r816_n200;
  tri   r816_n199;
  tri   r816_n198;
  tri   r816_n197;
  tri   r816_n195;
  tri   r816_n59;
  tri   r816_n61;
  tri   r816_n193;
  tri   r816_n192;
  tri   r816_n191;
  tri   r816_n190;
  tri   r816_n189;
  tri   r816_n188;
  tri   r816_n186;
  tri   r816_n129;
  tri   r816_n53;
  tri   r816_n185;
  tri   r816_n184;
  tri   r816_n183;
  tri   r816_n182;
  tri   r816_n180;
  tri   r816_n44;
  tri   r816_n46;
  tri   r816_n178;
  tri   r816_n177;
  tri   r816_n176;
  tri   r816_n175;
  tri   r816_n174;
  tri   r816_n173;
  tri   r816_n171;
  tri   r816_n131;
  tri   r816_n38;
  tri   r816_n170;
  tri   r816_n169;
  tri   r816_n168;
  tri   r816_n167;
  tri   r816_n165;
  tri   r816_n29;
  tri   r816_n31;
  tri   r816_n163;
  tri   r816_n162;
  tri   r816_n161;
  tri   r816_n160;
  tri   r816_n159;
  tri   r816_n158;
  tri   r816_n156;
  tri   r816_n133;
  tri   r816_n23;
  tri   r816_n155;
  tri   r816_n154;
  tri   r816_n153;
  tri   r816_n152;
  tri   r816_n150;
  tri   r816_n14;
  tri   r816_n16;
  tri   r816_n148;
  tri   r816_n147;
  tri   r816_n146;
  tri   r816_n145;
  tri   r816_n144;
  tri   r816_n143;
  tri   r816_n140;
  tri   r816_n8;
  tri   r816_n139;
  tri   r816_n6;
  tri   r816_n15;
  tri   r816_n9;
  tri   r816_n134;
  tri   r816_n19;
  tri   r816_n151;
  tri   r816_n30;
  tri   r816_n24;
  tri   r816_n132;
  tri   r816_n34;
  tri   r816_n166;
  tri   r816_n45;
  tri   r816_n39;
  tri   r816_n130;
  tri   r816_n49;
  tri   r816_n181;
  tri   r816_n60;
  tri   r816_n54;
  tri   r816_n128;
  tri   r816_n64;
  tri   r816_n196;
  tri   r816_n75;
  tri   r816_n69;
  tri   r816_n126;
  tri   r816_n79;
  tri   r816_n211;
  tri   r816_n94;
  tri   r816_n109;
  tri   r816_n120;
  tri   r816_n251;
  tri   r816_n250;
  tri   r816_n249;
  tri   r816_n248;
  tri   r816_n246;
  tri   r816_n121;
  tri   r816_n113;
  tri   r816_n245;
  tri   r816_n244;
  tri   r816_n243;
  tri   r816_n242;
  tri   r816_n241;
  tri   r816_n240;
  tri   r816_n122;
  tri   r816_n104;
  tri   r816_n106;
  tri   r816_n238;
  tri   r816_n237;
  tri   r816_n236;
  tri   r816_n235;
  tri   r816_n234;
  tri   r816_n99;
  tri   r816_n233;
  tri   r816_n105;
  tri   r816_n231;
  tri   r816_n123;
  tri   r816_n98;
  tri   r816_n230;
  tri   r816_n229;
  tri   r816_n228;
  tri   r816_n227;
  tri   r816_n226;
  tri   r816_n225;
  tri   r816_n124;
  tri   r816_n89;
  tri   r816_n91;
  tri   r816_n223;
  tri   r816_n222;
  tri   r816_n221;
  tri   r816_n220;
  tri   r816_n219;
  tri   r816_n84;
  tri   r816_n218;
  tri   r816_n90;
  tri   r816_n215;
  tri   r816_n125;
  tri   r816_n4;
  tri   r816_n276;
  tri   r816_n301;
  tri   r816_n304;
  tri   r816_n308;
  tri   P1_sub_111_n44;
  tri   P1_sub_111_n43;
  tri   P1_sub_111_n42;
  tri   P1_sub_111_n41;
  tri   P1_sub_111_n40;
  tri   P1_sub_111_n39;
  tri   P1_sub_111_n38;
  tri   P1_sub_111_n37;
  tri   P1_sub_111_n36;
  tri   P1_sub_111_n35;
  tri   P1_sub_111_n34;
  tri   P1_sub_111_n33;
  tri   P1_sub_111_n32;
  tri   P1_sub_111_n31;
  tri   P1_sub_111_n30;
  tri   P1_sub_111_n29;
  tri   P1_sub_111_n28;
  tri   P1_sub_111_n27;
  tri   P1_sub_111_n26;
  tri   P1_sub_111_n25;
  tri   P1_sub_111_n24;
  tri   P1_sub_111_n23;
  tri   P1_sub_111_n22;
  tri   P1_sub_111_n20;
  tri   P1_sub_111_n19;
  tri   P1_sub_111_n18;
  tri   P1_sub_111_n16;
  tri   P1_sub_111_n15;
  tri   P1_sub_111_n14;
  tri   P1_sub_111_n13;
  tri   P1_sub_111_n12;
  tri   P1_sub_111_n11;
  tri   P1_sub_111_n10;
  tri   P1_sub_111_n9;
  tri   P1_sub_111_n7;
  tri   P1_sub_111_n6;
  tri   P1_sub_111_n5;
  tri   P1_sub_111_n3;
  tri   P1_sub_111_n2;
  tri   P1_sub_111_n115;
  tri   P1_sub_111_n21;
  tri   P1_sub_111_n114;
  tri   P1_sub_111_n17;
  tri   P1_sub_111_n113;
  tri   P1_sub_111_n8;
  tri   P1_sub_111_n112;
  tri   P1_sub_111_n4;
  tri   P1_sub_111_n111;
  tri   P1_sub_111_n110;
  tri   P1_sub_111_n109;
  tri   P1_sub_111_n108;
  tri   P1_sub_111_n107;
  tri   P1_sub_111_n106;
  tri   P1_sub_111_n105;
  tri   P1_sub_111_n104;
  tri   P1_sub_111_n103;
  tri   P1_sub_111_n102;
  tri   P1_sub_111_n101;
  tri   P1_sub_111_n100;
  tri   P1_sub_111_n99;
  tri   P1_sub_111_n98;
  tri   P1_sub_111_n97;
  tri   P1_sub_111_n96;
  tri   P1_sub_111_n95;
  tri   P1_sub_111_n94;
  tri   P1_sub_111_n93;
  tri   P1_sub_111_n92;
  tri   P1_sub_111_n91;
  tri   P1_sub_111_n90;
  tri   P1_sub_111_n89;
  tri   P1_sub_111_n88;
  tri   P1_sub_111_n87;
  tri   P1_sub_111_n86;
  tri   P1_sub_111_n85;
  tri   P1_sub_111_n84;
  tri   P1_sub_111_n83;
  tri   P1_sub_111_n82;
  tri   P1_sub_111_n81;
  tri   P1_sub_111_n80;
  tri   P1_sub_111_n79;
  tri   P1_sub_111_n78;
  tri   P1_sub_111_n77;
  tri   P1_sub_111_n76;
  tri   P1_sub_111_n75;
  tri   P1_sub_111_n73;
  tri   P1_sub_111_n72;
  tri   P1_sub_111_n71;
  tri   P1_sub_111_n70;
  tri   P1_sub_111_n69;
  tri   P1_sub_111_n68;
  tri   P1_sub_111_n67;
  tri   P1_sub_111_n66;
  tri   P1_sub_111_n65;
  tri   P1_sub_111_n64;
  tri   P1_sub_111_n63;
  tri   P1_sub_111_n62;
  tri   P1_sub_111_n61;
  tri   P1_sub_111_n60;
  tri   P1_sub_111_n59;
  tri   P1_sub_111_n58;
  tri   P1_sub_111_n57;
  tri   P1_sub_111_n56;
  tri   P1_sub_111_n55;
  tri   P1_sub_111_n54;
  tri   P1_sub_111_n53;
  tri   P1_sub_111_n52;
  tri   P1_sub_111_n45;
  tri   P1_sub_111_n51;
  tri   P1_sub_111_n50;
  tri   P1_sub_111_n49;
  tri   P1_sub_111_n48;
  tri   P1_sub_111_n47;
  tri   P1_sub_111_n46;
  tri   r792_n77;
  tri   r792_n76;
  tri   r792_n75;
  tri   r792_n74;
  tri   r792_n73;
  tri   r792_n72;
  tri   r792_n70;
  tri   r792_n69;
  tri   r792_n68;
  tri   r792_n67;
  tri   r792_n66;
  tri   r792_n65;
  tri   r792_n64;
  tri   r792_n62;
  tri   r792_n61;
  tri   r792_n59;
  tri   r792_n58;
  tri   r792_n57;
  tri   r792_n55;
  tri   r792_n54;
  tri   r792_n53;
  tri   r792_n51;
  tri   r792_n50;
  tri   r792_n48;
  tri   r792_n47;
  tri   r792_n46;
  tri   r792_n44;
  tri   r792_n43;
  tri   r792_n41;
  tri   r792_n40;
  tri   r792_n39;
  tri   r792_n37;
  tri   r792_n36;
  tri   r792_n34;
  tri   r792_n33;
  tri   r792_n32;
  tri   r792_n30;
  tri   r792_n29;
  tri   r792_n27;
  tri   r792_n26;
  tri   r792_n25;
  tri   r792_n23;
  tri   r792_n22;
  tri   r792_n20;
  tri   r792_n19;
  tri   r792_n18;
  tri   r792_n16;
  tri   r792_n15;
  tri   r792_n13;
  tri   r792_n12;
  tri   r792_n11;
  tri   r792_n9;
  tri   r792_n8;
  tri   r792_n6;
  tri   r792_n5;
  tri   r792_n4;
  tri   r792_n2;
  tri   r792_n1;
  tri   r792_n162;
  tri   r792_n159;
  tri   r792_n158;
  tri   r792_n157;
  tri   r792_n156;
  tri   r792_n155;
  tri   r792_n154;
  tri   r792_n153;
  tri   r792_n152;
  tri   r792_n151;
  tri   r792_n149;
  tri   r792_n148;
  tri   r792_n147;
  tri   r792_n146;
  tri   r792_n145;
  tri   r792_n144;
  tri   r792_n143;
  tri   r792_n142;
  tri   r792_n141;
  tri   r792_n139;
  tri   r792_n138;
  tri   r792_n137;
  tri   r792_n136;
  tri   r792_n135;
  tri   r792_n134;
  tri   r792_n133;
  tri   r792_n132;
  tri   r792_n131;
  tri   r792_n129;
  tri   r792_n128;
  tri   r792_n127;
  tri   r792_n126;
  tri   r792_n125;
  tri   r792_n124;
  tri   r792_n123;
  tri   r792_n122;
  tri   r792_n121;
  tri   r792_n119;
  tri   r792_n118;
  tri   r792_n117;
  tri   r792_n116;
  tri   r792_n115;
  tri   r792_n114;
  tri   r792_n113;
  tri   r792_n112;
  tri   r792_n111;
  tri   r792_n109;
  tri   r792_n108;
  tri   r792_n107;
  tri   r792_n106;
  tri   r792_n105;
  tri   r792_n104;
  tri   r792_n103;
  tri   r792_n102;
  tri   r792_n101;
  tri   r792_n99;
  tri   r792_n98;
  tri   r792_n97;
  tri   r792_n96;
  tri   r792_n95;
  tri   r792_n94;
  tri   r792_n93;
  tri   r792_n92;
  tri   r792_n91;
  tri   r792_n89;
  tri   r792_n88;
  tri   r792_n87;
  tri   r792_n86;
  tri   r792_n85;
  tri   r792_n84;
  tri   r792_n83;
  tri   r792_n71;
  tri   r792_n82;
  tri   r792_n81;
  tri   r792_n78;
  tri   r792_n79;
  tri   r792_n189;
  tri   r792_n188;
  tri   r792_n60;
  tri   r792_n187;
  tri   r792_n186;
  tri   r792_n185;
  tri   r792_n52;
  tri   r792_n184;
  tri   r792_n183;
  tri   r792_n182;
  tri   r792_n45;
  tri   r792_n181;
  tri   r792_n180;
  tri   r792_n179;
  tri   r792_n38;
  tri   r792_n178;
  tri   r792_n177;
  tri   r792_n176;
  tri   r792_n31;
  tri   r792_n175;
  tri   r792_n174;
  tri   r792_n173;
  tri   r792_n24;
  tri   r792_n172;
  tri   r792_n171;
  tri   r792_n170;
  tri   r792_n17;
  tri   r792_n169;
  tri   r792_n168;
  tri   r792_n167;
  tri   r792_n10;
  tri   r792_n166;
  tri   r792_n165;
  tri   r792_n164;
  tri   r792_n161;
  tri   r792_n163;
  tri   r792_n3;
  tri   r793_n6;
  tri   r793_n5;
  tri   r793_n4;
  tri   r793_n2;
  tri   r793_n1;
  tri   r793_n99;
  tri   r793_n98;
  tri   r793_n97;
  tri   r793_n96;
  tri   r793_n95;
  tri   r793_n93;
  tri   r793_n92;
  tri   r793_n91;
  tri   r793_n89;
  tri   r793_n88;
  tri   r793_n87;
  tri   r793_n86;
  tri   r793_n85;
  tri   r793_n84;
  tri   r793_n83;
  tri   r793_n82;
  tri   r793_n81;
  tri   r793_n79;
  tri   r793_n78;
  tri   r793_n77;
  tri   r793_n76;
  tri   r793_n75;
  tri   r793_n74;
  tri   r793_n73;
  tri   r793_n72;
  tri   r793_n71;
  tri   r793_n70;
  tri   r793_n69;
  tri   r793_n68;
  tri   r793_n67;
  tri   r793_n66;
  tri   r793_n65;
  tri   r793_n64;
  tri   r793_n62;
  tri   r793_n61;
  tri   r793_n59;
  tri   r793_n58;
  tri   r793_n57;
  tri   r793_n55;
  tri   r793_n54;
  tri   r793_n53;
  tri   r793_n51;
  tri   r793_n50;
  tri   r793_n48;
  tri   r793_n47;
  tri   r793_n46;
  tri   r793_n44;
  tri   r793_n43;
  tri   r793_n41;
  tri   r793_n40;
  tri   r793_n39;
  tri   r793_n37;
  tri   r793_n36;
  tri   r793_n34;
  tri   r793_n33;
  tri   r793_n32;
  tri   r793_n30;
  tri   r793_n29;
  tri   r793_n27;
  tri   r793_n26;
  tri   r793_n25;
  tri   r793_n23;
  tri   r793_n22;
  tri   r793_n20;
  tri   r793_n19;
  tri   r793_n18;
  tri   r793_n16;
  tri   r793_n15;
  tri   r793_n13;
  tri   r793_n12;
  tri   r793_n8;
  tri   r793_n9;
  tri   r793_n11;
  tri   r793_n180;
  tri   r793_n38;
  tri   r793_n178;
  tri   r793_n177;
  tri   r793_n176;
  tri   r793_n31;
  tri   r793_n175;
  tri   r793_n174;
  tri   r793_n173;
  tri   r793_n24;
  tri   r793_n172;
  tri   r793_n171;
  tri   r793_n170;
  tri   r793_n17;
  tri   r793_n169;
  tri   r793_n168;
  tri   r793_n167;
  tri   r793_n10;
  tri   r793_n166;
  tri   r793_n165;
  tri   r793_n164;
  tri   r793_n3;
  tri   r793_n163;
  tri   r793_n162;
  tri   r793_n161;
  tri   r793_n159;
  tri   r793_n158;
  tri   r793_n157;
  tri   r793_n156;
  tri   r793_n155;
  tri   r793_n154;
  tri   r793_n153;
  tri   r793_n152;
  tri   r793_n151;
  tri   r793_n149;
  tri   r793_n148;
  tri   r793_n147;
  tri   r793_n146;
  tri   r793_n145;
  tri   r793_n144;
  tri   r793_n143;
  tri   r793_n142;
  tri   r793_n141;
  tri   r793_n139;
  tri   r793_n138;
  tri   r793_n137;
  tri   r793_n136;
  tri   r793_n135;
  tri   r793_n134;
  tri   r793_n133;
  tri   r793_n132;
  tri   r793_n131;
  tri   r793_n129;
  tri   r793_n128;
  tri   r793_n127;
  tri   r793_n126;
  tri   r793_n125;
  tri   r793_n124;
  tri   r793_n123;
  tri   r793_n122;
  tri   r793_n121;
  tri   r793_n119;
  tri   r793_n118;
  tri   r793_n117;
  tri   r793_n116;
  tri   r793_n115;
  tri   r793_n114;
  tri   r793_n113;
  tri   r793_n112;
  tri   r793_n111;
  tri   r793_n109;
  tri   r793_n108;
  tri   r793_n107;
  tri   r793_n106;
  tri   r793_n105;
  tri   r793_n104;
  tri   r793_n103;
  tri   r793_n94;
  tri   r793_n102;
  tri   r793_n101;
  tri   r793_n189;
  tri   r793_n188;
  tri   r793_n60;
  tri   r793_n187;
  tri   r793_n186;
  tri   r793_n185;
  tri   r793_n52;
  tri   r793_n184;
  tri   r793_n183;
  tri   r793_n182;
  tri   r793_n179;
  tri   r793_n181;
  tri   r793_n45;
  tri   add_1104_n309;
  tri   add_1104_n308;
  tri   add_1104_n310;
  tri   add_1104_n303;
  tri   add_1104_n304;
  tri   add_1104_n302;
  tri   add_1104_n305;
  tri   add_1104_n306;
  tri   add_1104_n307;
  tri   add_1104_n297;
  tri   add_1104_n298;
  tri   add_1104_n296;
  tri   add_1104_n299;
  tri   add_1104_n300;
  tri   add_1104_n301;
  tri   add_1104_n291;
  tri   add_1104_n292;
  tri   add_1104_n290;
  tri   add_1104_n293;
  tri   add_1104_n294;
  tri   add_1104_n295;
  tri   add_1104_n285;
  tri   add_1104_n286;
  tri   add_1104_n284;
  tri   add_1104_n287;
  tri   add_1104_n288;
  tri   add_1104_n289;
  tri   add_1104_n277;
  tri   add_1104_n279;
  tri   add_1104_n278;
  tri   add_1104_n280;
  tri   add_1104_n281;
  tri   add_1104_n282;
  tri   add_1104_n283;
  tri   add_1104_n270;
  tri   add_1104_n272;
  tri   add_1104_n273;
  tri   add_1104_n271;
  tri   add_1104_n274;
  tri   add_1104_n276;
  tri   add_1104_n275;
  tri   add_1104_n262;
  tri   add_1104_n263;
  tri   add_1104_n261;
  tri   add_1104_n266;
  tri   add_1104_n264;
  tri   add_1104_n265;
  tri   add_1104_n267;
  tri   add_1104_n269;
  tri   add_1104_n268;
  tri   add_1104_n256;
  tri   add_1104_n255;
  tri   add_1104_n257;
  tri   add_1104_n259;
  tri   add_1104_n258;
  tri   add_1104_n260;
  tri   add_1104_n249;
  tri   add_1104_n248;
  tri   add_1104_n250;
  tri   add_1104_n251;
  tri   add_1104_n252;
  tri   add_1104_n253;
  tri   add_1104_n254;
  tri   add_1104_n242;
  tri   add_1104_n243;
  tri   add_1104_n241;
  tri   add_1104_n245;
  tri   add_1104_n246;
  tri   add_1104_n247;
  tri   add_1104_n244;
  tri   add_1104_n233;
  tri   add_1104_n236;
  tri   add_1104_n234;
  tri   add_1104_n235;
  tri   add_1104_n237;
  tri   add_1104_n238;
  tri   add_1104_n239;
  tri   add_1104_n240;
  tri   add_1104_n226;
  tri   add_1104_n225;
  tri   add_1104_n227;
  tri   add_1104_n229;
  tri   add_1104_n228;
  tri   add_1104_n230;
  tri   add_1104_n232;
  tri   add_1104_n231;
  tri   add_1104_n219;
  tri   add_1104_n218;
  tri   add_1104_n220;
  tri   add_1104_n222;
  tri   add_1104_n223;
  tri   add_1104_n221;
  tri   add_1104_n224;
  tri   add_1104_n212;
  tri   add_1104_n213;
  tri   add_1104_n211;
  tri   add_1104_n216;
  tri   add_1104_n217;
  tri   add_1104_n214;
  tri   add_1104_n215;
  tri   add_1104_n206;
  tri   add_1104_n204;
  tri   add_1104_n205;
  tri   add_1104_n207;
  tri   add_1104_n209;
  tri   add_1104_n208;
  tri   add_1104_n210;
  tri   add_1104_n197;
  tri   add_1104_n199;
  tri   add_1104_n198;
  tri   add_1104_n200;
  tri   add_1104_n201;
  tri   add_1104_n202;
  tri   add_1104_n203;
  tri   add_1104_n190;
  tri   add_1104_n192;
  tri   add_1104_n193;
  tri   add_1104_n191;
  tri   add_1104_n194;
  tri   add_1104_n196;
  tri   add_1104_n195;
  tri   add_1104_n183;
  tri   add_1104_n182;
  tri   add_1104_n184;
  tri   add_1104_n186;
  tri   add_1104_n185;
  tri   add_1104_n187;
  tri   add_1104_n189;
  tri   add_1104_n188;
  tri   add_1104_n175;
  tri   add_1104_n176;
  tri   add_1104_n174;
  tri   add_1104_n177;
  tri   add_1104_n178;
  tri   add_1104_n179;
  tri   add_1104_n180;
  tri   add_1104_n181;
  tri   add_1104_n166;
  tri   add_1104_n169;
  tri   add_1104_n167;
  tri   add_1104_n168;
  tri   add_1104_n170;
  tri   add_1104_n171;
  tri   add_1104_n172;
  tri   add_1104_n173;
  tri   add_1104_n159;
  tri   add_1104_n158;
  tri   add_1104_n160;
  tri   add_1104_n162;
  tri   add_1104_n161;
  tri   add_1104_n163;
  tri   add_1104_n165;
  tri   add_1104_n164;
  tri   add_1104_n152;
  tri   add_1104_n151;
  tri   add_1104_n153;
  tri   add_1104_n155;
  tri   add_1104_n156;
  tri   add_1104_n154;
  tri   add_1104_n157;
  tri   add_1104_n145;
  tri   add_1104_n146;
  tri   add_1104_n144;
  tri   add_1104_n149;
  tri   add_1104_n150;
  tri   add_1104_n147;
  tri   add_1104_n148;
  tri   add_1104_n139;
  tri   add_1104_n137;
  tri   add_1104_n138;
  tri   add_1104_n140;
  tri   add_1104_n142;
  tri   add_1104_n141;
  tri   add_1104_n143;
  tri   add_1104_n130;
  tri   add_1104_n132;
  tri   add_1104_n131;
  tri   add_1104_n133;
  tri   add_1104_n134;
  tri   add_1104_n135;
  tri   add_1104_n136;
  tri   add_1104_n123;
  tri   add_1104_n125;
  tri   add_1104_n126;
  tri   add_1104_n124;
  tri   add_1104_n127;
  tri   add_1104_n129;
  tri   add_1104_n128;
  tri   add_1104_n115;
  tri   add_1104_n116;
  tri   add_1104_n114;
  tri   add_1104_n119;
  tri   add_1104_n117;
  tri   add_1104_n118;
  tri   add_1104_n120;
  tri   add_1104_n122;
  tri   add_1104_n121;
  tri   add_1104_n109;
  tri   add_1104_n108;
  tri   add_1104_n110;
  tri   add_1104_n112;
  tri   add_1104_n111;
  tri   add_1104_n113;
  tri   add_1104_n102;
  tri   add_1104_n101;
  tri   add_1104_n103;
  tri   add_1104_n104;
  tri   add_1104_n105;
  tri   add_1104_n106;
  tri   add_1104_n107;
  tri   add_1104_n95;
  tri   add_1104_n96;
  tri   add_1104_n94;
  tri   add_1104_n98;
  tri   add_1104_n99;
  tri   add_1104_n100;
  tri   add_1104_n97;
  tri   add_1104_n86;
  tri   add_1104_n89;
  tri   add_1104_n87;
  tri   add_1104_n88;
  tri   add_1104_n90;
  tri   add_1104_n91;
  tri   add_1104_n92;
  tri   add_1104_n93;
  tri   add_1104_n79;
  tri   add_1104_n78;
  tri   add_1104_n80;
  tri   add_1104_n82;
  tri   add_1104_n81;
  tri   add_1104_n83;
  tri   add_1104_n85;
  tri   add_1104_n84;
  tri   add_1104_n72;
  tri   add_1104_n73;
  tri   add_1104_n71;
  tri   add_1104_n74;
  tri   add_1104_n76;
  tri   add_1104_n75;
  tri   add_1104_n77;
  tri   add_1104_n65;
  tri   add_1104_n64;
  tri   add_1104_n66;
  tri   add_1104_n67;
  tri   add_1104_n68;
  tri   add_1104_n69;
  tri   add_1104_n70;
  tri   add_1104_n59;
  tri   add_1104_n58;
  tri   add_1104_n60;
  tri   add_1104_n61;
  tri   add_1104_n62;
  tri   add_1104_n63;
  tri   add_1104_n57;
  tri   add_1104_n49;
  tri   add_1104_n51;
  tri   add_1104_n53;
  tri   add_1104_n50;
  tri   add_1104_n52;
  tri   add_1104_n54;
  tri   add_1104_n55;
  tri   add_1104_n56;
  tri   add_1104_n41;
  tri   add_1104_n40;
  tri   add_1104_n42;
  tri   add_1104_n44;
  tri   add_1104_n45;
  tri   add_1104_n43;
  tri   add_1104_n46;
  tri   add_1104_n48;
  tri   add_1104_n47;
  tri   add_1104_n34;
  tri   add_1104_n33;
  tri   add_1104_n35;
  tri   add_1104_n37;
  tri   add_1104_n39;
  tri   add_1104_n38;
  tri   add_1104_n36;
  tri   add_1104_n24;
  tri   add_1104_n25;
  tri   add_1104_n27;
  tri   add_1104_n26;
  tri   add_1104_n28;
  tri   add_1104_n29;
  tri   add_1104_n30;
  tri   add_1104_n32;
  tri   add_1104_n31;
  tri   add_1104_n16;
  tri   add_1104_n17;
  tri   add_1104_n15;
  tri   add_1104_n18;
  tri   add_1104_n20;
  tri   add_1104_n19;
  tri   add_1104_n21;
  tri   add_1104_n23;
  tri   add_1104_n22;
  tri   add_1104_n9;
  tri   add_1104_n10;
  tri   add_1104_n8;
  tri   add_1104_n11;
  tri   add_1104_n13;
  tri   add_1104_n12;
  tri   add_1104_n14;
  tri   add_1104_n2;
  tri   add_1104_n3;
  tri   add_1104_n1;
  tri   add_1104_n4;
  tri   add_1104_n6;
  tri   add_1104_n5;
  tri   add_1104_n7;
  tri   r794_n26;
  tri   r794_n25;
  tri   r794_n24;
  tri   r794_n23;
  tri   r794_n22;
  tri   r794_n20;
  tri   r794_n19;
  tri   r794_n18;
  tri   r794_n16;
  tri   r794_n15;
  tri   r794_n14;
  tri   r794_n13;
  tri   r794_n12;
  tri   r794_n11;
  tri   r794_n10;
  tri   r794_n9;
  tri   r794_n7;
  tri   r794_n6;
  tri   r794_n5;
  tri   r794_n3;
  tri   r794_n2;
  tri   r794_n100;
  tri   r794_n99;
  tri   r794_n98;
  tri   r794_n97;
  tri   r794_n96;
  tri   r794_n95;
  tri   r794_n94;
  tri   r794_n93;
  tri   r794_n92;
  tri   r794_n91;
  tri   r794_n90;
  tri   r794_n89;
  tri   r794_n88;
  tri   r794_n87;
  tri   r794_n86;
  tri   r794_n85;
  tri   r794_n84;
  tri   r794_n83;
  tri   r794_n82;
  tri   r794_n81;
  tri   r794_n80;
  tri   r794_n79;
  tri   r794_n78;
  tri   r794_n77;
  tri   r794_n76;
  tri   r794_n75;
  tri   r794_n73;
  tri   r794_n72;
  tri   r794_n71;
  tri   r794_n70;
  tri   r794_n69;
  tri   r794_n68;
  tri   r794_n67;
  tri   r794_n66;
  tri   r794_n65;
  tri   r794_n64;
  tri   r794_n63;
  tri   r794_n62;
  tri   r794_n61;
  tri   r794_n60;
  tri   r794_n59;
  tri   r794_n58;
  tri   r794_n57;
  tri   r794_n56;
  tri   r794_n55;
  tri   r794_n54;
  tri   r794_n53;
  tri   r794_n52;
  tri   r794_n51;
  tri   r794_n50;
  tri   r794_n49;
  tri   r794_n48;
  tri   r794_n47;
  tri   r794_n46;
  tri   r794_n45;
  tri   r794_n44;
  tri   r794_n43;
  tri   r794_n42;
  tri   r794_n41;
  tri   r794_n40;
  tri   r794_n39;
  tri   r794_n38;
  tri   r794_n37;
  tri   r794_n36;
  tri   r794_n35;
  tri   r794_n34;
  tri   r794_n33;
  tri   r794_n32;
  tri   r794_n31;
  tri   r794_n30;
  tri   r794_n28;
  tri   r794_n27;
  tri   r794_n29;
  tri   r794_n115;
  tri   r794_n21;
  tri   r794_n114;
  tri   r794_n17;
  tri   r794_n113;
  tri   r794_n8;
  tri   r794_n112;
  tri   r794_n4;
  tri   r794_n111;
  tri   r794_n110;
  tri   r794_n109;
  tri   r794_n108;
  tri   r794_n107;
  tri   r794_n106;
  tri   r794_n105;
  tri   r794_n101;
  tri   r794_n102;
  tri   r794_n104;
  tri   r794_n103;
  tri   P1_add_122_n57;
  tri   P1_add_122_n56;
  tri   P1_add_122_n55;
  tri   P1_add_122_n54;
  tri   P1_add_122_n52;
  tri   P1_add_122_n51;
  tri   P1_add_122_n50;
  tri   P1_add_122_n49;
  tri   P1_add_122_n48;
  tri   P1_add_122_n47;
  tri   P1_add_122_n46;
  tri   P1_add_122_n45;
  tri   P1_add_122_n44;
  tri   P1_add_122_n43;
  tri   P1_add_122_n42;
  tri   P1_add_122_n41;
  tri   P1_add_122_n40;
  tri   P1_add_122_n39;
  tri   P1_add_122_n38;
  tri   P1_add_122_n37;
  tri   P1_add_122_n36;
  tri   P1_add_122_n35;
  tri   P1_add_122_n34;
  tri   P1_add_122_n33;
  tri   P1_add_122_n32;
  tri   P1_add_122_n31;
  tri   P1_add_122_n30;
  tri   P1_add_122_n29;
  tri   P1_add_122_n28;
  tri   P1_add_122_n27;
  tri   P1_add_122_n26;
  tri   P1_add_122_n25;
  tri   P1_add_122_n24;
  tri   P1_add_122_n22;
  tri   P1_add_122_n21;
  tri   P1_add_122_n20;
  tri   P1_add_122_n19;
  tri   P1_add_122_n18;
  tri   P1_add_122_n17;
  tri   P1_add_122_n16;
  tri   P1_add_122_n13;
  tri   P1_add_122_n12;
  tri   P1_add_122_n11;
  tri   P1_add_122_n10;
  tri   P1_add_122_n9;
  tri   P1_add_122_n6;
  tri   P1_add_122_n23;
  tri   P1_add_122_n102;
  tri   P1_add_122_n14;
  tri   P1_add_122_n15;
  tri   P1_add_122_n101;
  tri   P1_add_122_n7;
  tri   P1_add_122_n8;
  tri   P1_add_122_n100;
  tri   P1_add_122_n99;
  tri   P1_add_122_n98;
  tri   P1_add_122_n97;
  tri   P1_add_122_n96;
  tri   P1_add_122_n95;
  tri   P1_add_122_n94;
  tri   P1_add_122_n93;
  tri   P1_add_122_n92;
  tri   P1_add_122_n91;
  tri   P1_add_122_n90;
  tri   P1_add_122_n89;
  tri   P1_add_122_n88;
  tri   P1_add_122_n87;
  tri   P1_add_122_n86;
  tri   P1_add_122_n85;
  tri   P1_add_122_n84;
  tri   P1_add_122_n83;
  tri   P1_add_122_n82;
  tri   P1_add_122_n81;
  tri   P1_add_122_n80;
  tri   P1_add_122_n79;
  tri   P1_add_122_n78;
  tri   P1_add_122_n77;
  tri   P1_add_122_n76;
  tri   P1_add_122_n75;
  tri   P1_add_122_n74;
  tri   P1_add_122_n73;
  tri   P1_add_122_n72;
  tri   P1_add_122_n71;
  tri   P1_add_122_n70;
  tri   P1_add_122_n69;
  tri   P1_add_122_n68;
  tri   P1_add_122_n67;
  tri   P1_add_122_n66;
  tri   P1_add_122_n65;
  tri   P1_add_122_n64;
  tri   P1_add_122_n63;
  tri   P1_add_122_n62;
  tri   P1_add_122_n61;
  tri   P1_add_122_n60;
  tri   P1_add_122_n58;
  tri   P1_add_122_n59;
  tri   P1_add_122_n53;
  tri   P1_add_122_n5;
  tri   P1_add_122_n4;
  tri   r796_n13;
  tri   r796_n12;
  tri   r796_n11;
  tri   r796_n9;
  tri   r796_n8;
  tri   r796_n6;
  tri   r796_n5;
  tri   r796_n4;
  tri   r796_n2;
  tri   r796_n1;
  tri   r796_n102;
  tri   r796_n101;
  tri   r796_n100;
  tri   r796_n99;
  tri   r796_n98;
  tri   r796_n97;
  tri   r796_n96;
  tri   r796_n95;
  tri   r796_n94;
  tri   r796_n92;
  tri   r796_n91;
  tri   r796_n90;
  tri   r796_n89;
  tri   r796_n88;
  tri   r796_n87;
  tri   r796_n86;
  tri   r796_n85;
  tri   r796_n84;
  tri   r796_n82;
  tri   r796_n81;
  tri   r796_n80;
  tri   r796_n79;
  tri   r796_n78;
  tri   r796_n77;
  tri   r796_n76;
  tri   r796_n75;
  tri   r796_n74;
  tri   r796_n72;
  tri   r796_n71;
  tri   r796_n70;
  tri   r796_n69;
  tri   r796_n68;
  tri   r796_n66;
  tri   r796_n65;
  tri   r796_n64;
  tri   r796_n63;
  tri   r796_n62;
  tri   r796_n61;
  tri   r796_n60;
  tri   r796_n59;
  tri   r796_n58;
  tri   r796_n57;
  tri   r796_n55;
  tri   r796_n54;
  tri   r796_n53;
  tri   r796_n51;
  tri   r796_n50;
  tri   r796_n48;
  tri   r796_n47;
  tri   r796_n46;
  tri   r796_n44;
  tri   r796_n43;
  tri   r796_n41;
  tri   r796_n40;
  tri   r796_n39;
  tri   r796_n37;
  tri   r796_n36;
  tri   r796_n34;
  tri   r796_n33;
  tri   r796_n32;
  tri   r796_n30;
  tri   r796_n29;
  tri   r796_n27;
  tri   r796_n26;
  tri   r796_n25;
  tri   r796_n23;
  tri   r796_n22;
  tri   r796_n20;
  tri   r796_n19;
  tri   r796_n15;
  tri   r796_n16;
  tri   r796_n18;
  tri   r796_n189;
  tri   r796_n188;
  tri   r796_n187;
  tri   r796_n186;
  tri   r796_n185;
  tri   r796_n183;
  tri   r796_n182;
  tri   r796_n181;
  tri   r796_n179;
  tri   r796_n178;
  tri   r796_n177;
  tri   r796_n176;
  tri   r796_n175;
  tri   r796_n174;
  tri   r796_n173;
  tri   r796_n172;
  tri   r796_n171;
  tri   r796_n169;
  tri   r796_n168;
  tri   r796_n167;
  tri   r796_n166;
  tri   r796_n165;
  tri   r796_n163;
  tri   r796_n162;
  tri   r796_n160;
  tri   r796_n159;
  tri   r796_n158;
  tri   r796_n157;
  tri   r796_n156;
  tri   r796_n155;
  tri   r796_n154;
  tri   r796_n152;
  tri   r796_n151;
  tri   r796_n150;
  tri   r796_n149;
  tri   r796_n148;
  tri   r796_n147;
  tri   r796_n146;
  tri   r796_n145;
  tri   r796_n144;
  tri   r796_n142;
  tri   r796_n141;
  tri   r796_n140;
  tri   r796_n139;
  tri   r796_n138;
  tri   r796_n137;
  tri   r796_n136;
  tri   r796_n135;
  tri   r796_n134;
  tri   r796_n132;
  tri   r796_n131;
  tri   r796_n130;
  tri   r796_n129;
  tri   r796_n128;
  tri   r796_n127;
  tri   r796_n126;
  tri   r796_n125;
  tri   r796_n124;
  tri   r796_n122;
  tri   r796_n121;
  tri   r796_n120;
  tri   r796_n119;
  tri   r796_n118;
  tri   r796_n117;
  tri   r796_n116;
  tri   r796_n115;
  tri   r796_n114;
  tri   r796_n112;
  tri   r796_n111;
  tri   r796_n110;
  tri   r796_n109;
  tri   r796_n108;
  tri   r796_n104;
  tri   r796_n107;
  tri   r796_n105;
  tri   r796_n106;
  tri   r796_n272;
  tri   r796_n271;
  tri   r796_n270;
  tri   r796_n17;
  tri   r796_n269;
  tri   r796_n268;
  tri   r796_n267;
  tri   r796_n10;
  tri   r796_n266;
  tri   r796_n265;
  tri   r796_n264;
  tri   r796_n3;
  tri   r796_n263;
  tri   r796_n262;
  tri   r796_n261;
  tri   r796_n259;
  tri   r796_n258;
  tri   r796_n257;
  tri   r796_n256;
  tri   r796_n255;
  tri   r796_n254;
  tri   r796_n253;
  tri   r796_n252;
  tri   r796_n251;
  tri   r796_n249;
  tri   r796_n248;
  tri   r796_n247;
  tri   r796_n246;
  tri   r796_n245;
  tri   r796_n244;
  tri   r796_n243;
  tri   r796_n242;
  tri   r796_n241;
  tri   r796_n239;
  tri   r796_n238;
  tri   r796_n237;
  tri   r796_n236;
  tri   r796_n235;
  tri   r796_n234;
  tri   r796_n233;
  tri   r796_n232;
  tri   r796_n231;
  tri   r796_n229;
  tri   r796_n228;
  tri   r796_n227;
  tri   r796_n226;
  tri   r796_n225;
  tri   r796_n224;
  tri   r796_n223;
  tri   r796_n222;
  tri   r796_n221;
  tri   r796_n219;
  tri   r796_n218;
  tri   r796_n217;
  tri   r796_n216;
  tri   r796_n215;
  tri   r796_n214;
  tri   r796_n213;
  tri   r796_n212;
  tri   r796_n211;
  tri   r796_n209;
  tri   r796_n208;
  tri   r796_n207;
  tri   r796_n206;
  tri   r796_n205;
  tri   r796_n204;
  tri   r796_n203;
  tri   r796_n202;
  tri   r796_n201;
  tri   r796_n199;
  tri   r796_n198;
  tri   r796_n197;
  tri   r796_n196;
  tri   r796_n195;
  tri   r796_n194;
  tri   r796_n193;
  tri   r796_n184;
  tri   r796_n192;
  tri   r796_n191;
  tri   r796_n289;
  tri   r796_n288;
  tri   r796_n161;
  tri   r796_n287;
  tri   r796_n286;
  tri   r796_n285;
  tri   r796_n52;
  tri   r796_n284;
  tri   r796_n283;
  tri   r796_n282;
  tri   r796_n45;
  tri   r796_n281;
  tri   r796_n280;
  tri   r796_n279;
  tri   r796_n38;
  tri   r796_n278;
  tri   r796_n277;
  tri   r796_n276;
  tri   r796_n31;
  tri   r796_n275;
  tri   r796_n24;
  tri   r796_n274;
  tri   r796_n273;
  tri   r798_n55;
  tri   r798_n54;
  tri   r798_n53;
  tri   r798_n51;
  tri   r798_n50;
  tri   r798_n48;
  tri   r798_n47;
  tri   r798_n46;
  tri   r798_n44;
  tri   r798_n43;
  tri   r798_n41;
  tri   r798_n40;
  tri   r798_n39;
  tri   r798_n37;
  tri   r798_n36;
  tri   r798_n34;
  tri   r798_n33;
  tri   r798_n32;
  tri   r798_n30;
  tri   r798_n29;
  tri   r798_n27;
  tri   r798_n26;
  tri   r798_n25;
  tri   r798_n23;
  tri   r798_n22;
  tri   r798_n20;
  tri   r798_n19;
  tri   r798_n18;
  tri   r798_n16;
  tri   r798_n15;
  tri   r798_n13;
  tri   r798_n12;
  tri   r798_n11;
  tri   r798_n9;
  tri   r798_n8;
  tri   r798_n6;
  tri   r798_n5;
  tri   r798_n4;
  tri   r798_n2;
  tri   r798_n1;
  tri   r798_n142;
  tri   r798_n140;
  tri   r798_n139;
  tri   r798_n138;
  tri   r798_n136;
  tri   r798_n135;
  tri   r798_n134;
  tri   r798_n132;
  tri   r798_n131;
  tri   r798_n130;
  tri   r798_n129;
  tri   r798_n128;
  tri   r798_n127;
  tri   r798_n126;
  tri   r798_n125;
  tri   r798_n124;
  tri   r798_n122;
  tri   r798_n121;
  tri   r798_n120;
  tri   r798_n119;
  tri   r798_n118;
  tri   r798_n117;
  tri   r798_n116;
  tri   r798_n115;
  tri   r798_n114;
  tri   r798_n112;
  tri   r798_n111;
  tri   r798_n110;
  tri   r798_n109;
  tri   r798_n108;
  tri   r798_n107;
  tri   r798_n106;
  tri   r798_n105;
  tri   r798_n104;
  tri   r798_n102;
  tri   r798_n101;
  tri   r798_n100;
  tri   r798_n99;
  tri   r798_n98;
  tri   r798_n97;
  tri   r798_n96;
  tri   r798_n95;
  tri   r798_n94;
  tri   r798_n92;
  tri   r798_n91;
  tri   r798_n90;
  tri   r798_n89;
  tri   r798_n88;
  tri   r798_n87;
  tri   r798_n86;
  tri   r798_n85;
  tri   r798_n84;
  tri   r798_n82;
  tri   r798_n81;
  tri   r798_n80;
  tri   r798_n79;
  tri   r798_n78;
  tri   r798_n77;
  tri   r798_n76;
  tri   r798_n75;
  tri   r798_n74;
  tri   r798_n72;
  tri   r798_n71;
  tri   r798_n70;
  tri   r798_n69;
  tri   r798_n68;
  tri   r798_n66;
  tri   r798_n65;
  tri   r798_n64;
  tri   r798_n63;
  tri   r798_n62;
  tri   r798_n61;
  tri   r798_n60;
  tri   r798_n59;
  tri   r798_n58;
  tri   r798_n57;
  tri   r798_n227;
  tri   r798_n226;
  tri   r798_n225;
  tri   r798_n223;
  tri   r798_n222;
  tri   r798_n221;
  tri   r798_n219;
  tri   r798_n218;
  tri   r798_n217;
  tri   r798_n216;
  tri   r798_n215;
  tri   r798_n214;
  tri   r798_n213;
  tri   r798_n212;
  tri   r798_n211;
  tri   r798_n209;
  tri   r798_n208;
  tri   r798_n207;
  tri   r798_n206;
  tri   r798_n205;
  tri   r798_n204;
  tri   r798_n203;
  tri   r798_n202;
  tri   r798_n201;
  tri   r798_n199;
  tri   r798_n198;
  tri   r798_n197;
  tri   r798_n196;
  tri   r798_n195;
  tri   r798_n194;
  tri   r798_n193;
  tri   r798_n192;
  tri   r798_n191;
  tri   r798_n189;
  tri   r798_n188;
  tri   r798_n187;
  tri   r798_n186;
  tri   r798_n185;
  tri   r798_n184;
  tri   r798_n183;
  tri   r798_n182;
  tri   r798_n181;
  tri   r798_n179;
  tri   r798_n178;
  tri   r798_n177;
  tri   r798_n176;
  tri   r798_n175;
  tri   r798_n174;
  tri   r798_n173;
  tri   r798_n172;
  tri   r798_n171;
  tri   r798_n169;
  tri   r798_n168;
  tri   r798_n167;
  tri   r798_n166;
  tri   r798_n165;
  tri   r798_n163;
  tri   r798_n162;
  tri   r798_n160;
  tri   r798_n159;
  tri   r798_n158;
  tri   r798_n157;
  tri   r798_n156;
  tri   r798_n155;
  tri   r798_n154;
  tri   r798_n152;
  tri   r798_n151;
  tri   r798_n150;
  tri   r798_n149;
  tri   r798_n148;
  tri   r798_n147;
  tri   r798_n146;
  tri   r798_n137;
  tri   r798_n145;
  tri   r798_n144;
  tri   r798_n141;
  tri   r798_n289;
  tri   r798_n288;
  tri   r798_n161;
  tri   r798_n287;
  tri   r798_n286;
  tri   r798_n285;
  tri   r798_n52;
  tri   r798_n284;
  tri   r798_n283;
  tri   r798_n282;
  tri   r798_n45;
  tri   r798_n281;
  tri   r798_n280;
  tri   r798_n279;
  tri   r798_n38;
  tri   r798_n278;
  tri   r798_n277;
  tri   r798_n276;
  tri   r798_n31;
  tri   r798_n275;
  tri   r798_n274;
  tri   r798_n273;
  tri   r798_n24;
  tri   r798_n272;
  tri   r798_n271;
  tri   r798_n270;
  tri   r798_n17;
  tri   r798_n269;
  tri   r798_n268;
  tri   r798_n267;
  tri   r798_n10;
  tri   r798_n266;
  tri   r798_n265;
  tri   r798_n264;
  tri   r798_n3;
  tri   r798_n263;
  tri   r798_n262;
  tri   r798_n261;
  tri   r798_n259;
  tri   r798_n258;
  tri   r798_n257;
  tri   r798_n256;
  tri   r798_n255;
  tri   r798_n254;
  tri   r798_n253;
  tri   r798_n252;
  tri   r798_n251;
  tri   r798_n249;
  tri   r798_n248;
  tri   r798_n247;
  tri   r798_n246;
  tri   r798_n245;
  tri   r798_n244;
  tri   r798_n243;
  tri   r798_n242;
  tri   r798_n241;
  tri   r798_n239;
  tri   r798_n238;
  tri   r798_n237;
  tri   r798_n236;
  tri   r798_n235;
  tri   r798_n234;
  tri   r798_n233;
  tri   r798_n224;
  tri   r798_n232;
  tri   r798_n231;
  tri   r798_n228;
  tri   r798_n229;
  tri   r798_n314;

  NBUFFX2 CBUFNBUFFX32_G1B2I1 ( .Z(clock_G1B2I1_1), .INP(clock_G1B1I2_1) );
  NBUFFX16 CBUFNBUFFX32_G1B1I1_1 ( .Z(clock_G1B1I1_1), .INP(clock) );
  NBUFFX2 CBUFNBUFFX32_G1B2I38 ( .Z(clock_G1B2I38_1), .INP(clock_G1B1I2_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I37 ( .Z(clock_G1B2I37_1), .INP(clock_G1B1I2_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I34 ( .Z(clock_G1B2I34_1), .INP(clock_G1B1I2_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I33 ( .Z(clock_G1B2I33_1), .INP(clock_G1B1I1_1) );
  NBUFFX4 CBUFNBUFFX32_G1B2I36 ( .Z(clock_G1B2I36_1), .INP(clock_G1B1I3_1) );
  NBUFFX4 CBUFNBUFFX32_G1B2I32 ( .Z(clock_G1B2I32_1), .INP(clock_G1B1I1_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I27 ( .Z(clock_G1B2I27_1), .INP(clock_G1B1I1_1) );
  NBUFFX8 CBUFNBUFFX32_G1B2I35 ( .Z(clock_G1B2I35_1), .INP(clock_G1B1I3_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I15 ( .Z(clock_G1B2I15_1), .INP(clock_G1B1I1_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I31 ( .Z(clock_G1B2I31_1), .INP(clock_G1B1I2_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I9 ( .Z(clock_G1B2I9_1), .INP(clock_G1B1I1_1) );
  NBUFFX4 CBUFNBUFFX32_G1B2I30 ( .Z(clock_G1B2I30_1), .INP(clock_G1B1I3_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I29 ( .Z(clock_G1B2I29_1), .INP(clock_G1B1I2_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I17 ( .Z(clock_G1B2I17_1), .INP(clock_G1B1I3_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I21 ( .Z(clock_G1B2I21_1), .INP(clock_G1B1I2_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I23 ( .Z(clock_G1B2I23_1), .INP(clock_G1B1I2_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I28 ( .Z(clock_G1B2I28_1), .INP(clock_G1B1I2_1) );
  NBUFFX4 CBUFNBUFFX32_G1B2I14 ( .Z(clock_G1B2I14_1), .INP(clock_G1B1I3_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I26 ( .Z(clock_G1B2I26_1), .INP(clock_G1B1I1_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I18 ( .Z(clock_G1B2I18_1), .INP(clock_G1B1I3_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I12 ( .Z(clock_G1B2I12_1), .INP(clock_G1B1I1_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I13 ( .Z(clock_G1B2I13_1), .INP(clock_G1B1I3_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I24 ( .Z(clock_G1B2I24_1), .INP(clock_G1B1I1_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I25 ( .Z(clock_G1B2I25_1), .INP(clock_G1B1I1_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I3 ( .Z(clock_G1B2I3_1), .INP(clock_G1B1I1_1) );
  NBUFFX4 CBUFNBUFFX32_G1B2I22 ( .Z(clock_G1B2I22_1), .INP(clock_G1B1I1_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I20 ( .Z(clock_G1B2I20_1), .INP(clock_G1B1I2_1) );
  NBUFFX8 CBUFNBUFFX32_G1B2I19 ( .Z(clock_G1B2I19_1), .INP(clock_G1B1I3_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I8 ( .Z(clock_G1B2I8_1), .INP(clock_G1B1I2_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I16 ( .Z(clock_G1B2I16_1), .INP(clock_G1B1I1_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I7 ( .Z(clock_G1B2I7_1), .INP(clock_G1B1I3_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I11 ( .Z(clock_G1B2I11_1), .INP(clock_G1B1I2_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I2 ( .Z(clock_G1B2I2_1), .INP(clock_G1B1I2_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I4 ( .Z(clock_G1B2I4_1), .INP(clock_G1B1I2_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I6 ( .Z(clock_G1B2I6_1), .INP(clock_G1B1I1_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I5 ( .Z(clock_G1B2I5_1), .INP(clock_G1B1I1_1) );
  NBUFFX2 CBUFNBUFFX32_G1B2I10 ( .Z(clock_G1B2I10_1), .INP(clock_G1B1I2_1) );
  NBUFFX8 CBUFNBUFFX8_G1B1I3 ( .Z(clock_G1B1I3_1), .INP(clock) );
  NBUFFX16 CBUFNBUFFX16_G1B1I2 ( .Z(clock_G1B1I2_1), .INP(clock) );
  INVX2 U1655 ( .INP(P2_N5470), .ZN(n6729) );
  NBUFFX8 U1857 ( .Z(n6931), .INP(n7460) );
  NBUFFX8 U1893 ( .Z(n6967), .INP(P2_N294) );
  NBUFFX8 U1631 ( .Z(n6705), .INP(n7480) );
  INVX2 U1933 ( .INP(n7462), .ZN(n7007) );
  NBUFFX4 U1619 ( .Z(n6693), .INP(n7479) );
  NBUFFX8 U2088 ( .Z(n7162), .INP(P2_N5077) );
  SDFFARX1 P1_state_reg ( .QN(n4169), .CLK(clock_G1B2I2_1), .RSTB(n7580), 
        .SE(n7582), .SI(n18293), .D(n6580) );
  SDFFARX1 P2_state_reg ( .QN(n2166), .CLK(clock_G1B2I25_1), .RSTB(n7501), 
        .SE(n6573), .SI(n18762), .D(n6589) );
  INVX0 U399 ( .ZN(n6596), .INP(n18345) );
  INVX0 U400 ( .ZN(n6597), .INP(n18343) );
  INVX0 U401 ( .ZN(n6598), .INP(n18341) );
  INVX0 U438 ( .ZN(n6624), .INP(n18695) );
  INVX0 U398 ( .ZN(n6595), .INP(n18347) );
  NBUFFX4 U1641 ( .Z(n6715), .INP(n7480) );
  NBUFFX2 U1625 ( .Z(n6699), .INP(n7479) );
  NBUFFX2 U1611 ( .Z(n6685), .INP(n7479) );
  NBUFFX4 U1629 ( .Z(n6703), .INP(n7480) );
  INVX0 U1642 ( .ZN(n6716), .INP(n6715) );
  INVX0 U1614 ( .ZN(n6688), .INP(n6687) );
  INVX0 U1632 ( .ZN(n6706), .INP(n6705) );
  INVX0 U1630 ( .ZN(n6704), .INP(n6703) );
  INVX0 U1638 ( .ZN(n6712), .INP(n7480) );
  INVX0 U1620 ( .ZN(n6694), .INP(n6693) );
  INVX0 U1616 ( .ZN(n6690), .INP(n19025) );
  INVX0 U1644 ( .ZN(n6718), .INP(n6705) );
  INVX0 U1618 ( .ZN(n6692), .INP(n7479) );
  INVX0 U1634 ( .ZN(n6708), .INP(n19009) );
  INVX0 U1636 ( .ZN(n6710), .INP(n19009) );
  INVX2 U1663 ( .INP(n6736), .ZN(n6737) );
  INVX0 U1665 ( .ZN(n6739), .INP(N5) );
  INVX0 U435 ( .ZN(n6621), .INP(n18465) );
  INVX0 U1607 ( .ZN(n6681), .INP(n18819) );
  NOR2X1 U6803 ( .QN(n4480), .IN1(n4615), .IN2(n4616) );
  NOR2X1 U3937 ( .QN(n2569), .IN1(n2660), .IN2(n2661) );
  INVX0 U436 ( .ZN(n6622), .INP(n18459) );
  INVX0 U1608 ( .ZN(n6682), .INP(n18817) );
  NOR2X1 U8710 ( .QN(P1_N583), .IN1(n4157), .IN2(n4158) );
  NOR2X1 U5620 ( .QN(n2693), .IN1(n2153), .IN2(n2154) );
  NOR2X0 U6790 ( .QN(n4803), .IN1(n4804), .IN2(n4805) );
  NOR2X0 U3924 ( .QN(n2919), .IN1(n2920), .IN2(n2921) );
  INVX2 U1960 ( .INP(n4803), .ZN(n7034) );
  INVX0 U1961 ( .ZN(n7035), .INP(n2919) );
  INVX0 U1609 ( .ZN(n6683), .INP(n18815) );
  INVX0 U437 ( .ZN(n6623), .INP(n18455) );
  INVX0 U2112 ( .ZN(n7186), .INP(P2_N5072) );
  INVX0 U1974 ( .ZN(n7048), .INP(P1_N5150) );
  INVX0 U1977 ( .ZN(n7051), .INP(P1_N5150) );
  INVX0 U2110 ( .ZN(n7184), .INP(P2_N5072) );
  NBUFFX8 U2006 ( .Z(n7080), .INP(P1_N5155) );
  INVX2 U2207 ( .INP(P1_N5147), .ZN(n7281) );
  INVX0 U1971 ( .ZN(n7045), .INP(P1_N5151) );
  INVX0 U1969 ( .ZN(n7043), .INP(P1_N5152) );
  INVX0 U2005 ( .ZN(n7079), .INP(P1_N5155) );
  NBUFFX8 U1992 ( .Z(n7066), .INP(P1_N5159) );
  INVX0 U2002 ( .ZN(n7076), .INP(n7075) );
  INVX0 U2083 ( .ZN(n7157), .INP(P2_N5078) );
  INVX0 U2079 ( .ZN(n7153), .INP(P2_N5079) );
  INVX0 U2145 ( .ZN(n7219), .INP(n7220) );
  INVX0 U2075 ( .ZN(n7149), .INP(P2_N5080) );
  NBUFFX4 U2135 ( .Z(n7209), .INP(P2_N5084) );
  NBUFFX4 U2132 ( .Z(n7206), .INP(P2_N5085) );
  INVX0 U1984 ( .ZN(n7058), .INP(P1_N5161) );
  INVX0 U2137 ( .ZN(n7211), .INP(n7210) );
  INVX0 U2041 ( .ZN(n7115), .INP(P1_N5163) );
  INVX0 U2134 ( .ZN(n7208), .INP(P2_N5084) );
  INVX0 U2131 ( .ZN(n7205), .INP(P2_N5085) );
  INVX0 U2038 ( .ZN(n7112), .INP(P1_N5164) );
  INVX0 U2127 ( .ZN(n7201), .INP(P2_N5086) );
  INVX0 U2123 ( .ZN(n7197), .INP(P2_N5087) );
  INVX0 U2035 ( .ZN(n7109), .INP(P1_N5165) );
  NBUFFX8 U2113 ( .Z(n7187), .INP(P2_N5089) );
  INVX0 U2028 ( .ZN(n7102), .INP(P1_N5167) );
  INVX0 U2031 ( .ZN(n7105), .INP(P1_N5166) );
  NBUFFX8 U2189 ( .Z(n7263), .INP(P2_N5090) );
  INVX0 U2024 ( .ZN(n7098), .INP(n7099) );
  INVX0 U2237 ( .ZN(n7311), .INP(n2205) );
  INVX0 U2021 ( .ZN(n7095), .INP(P1_N5169) );
  INVX2 U1941 ( .INP(P2_N914), .ZN(n7015) );
  INVX0 U2240 ( .ZN(n7314), .INP(n4202) );
  INVX0 U2241 ( .ZN(n7315), .INP(n2199) );
  INVX0 U2239 ( .ZN(n7313), .INP(n2202) );
  INVX0 U2018 ( .ZN(n7092), .INP(P1_N5170) );
  INVX0 U2242 ( .ZN(n7316), .INP(n4199) );
  INVX0 U2243 ( .ZN(n7317), .INP(n2196) );
  INVX0 U2244 ( .ZN(n7318), .INP(n4196) );
  INVX0 U2245 ( .ZN(n7319), .INP(n2193) );
  INVX0 U2248 ( .ZN(n7322), .INP(n4190) );
  INVX0 U2246 ( .ZN(n7320), .INP(n4193) );
  INVX0 U2249 ( .ZN(n7323), .INP(n2187) );
  INVX0 U2247 ( .ZN(n7321), .INP(n2190) );
  INVX0 U2250 ( .ZN(n7324), .INP(n4187) );
  INVX0 U2251 ( .ZN(n7325), .INP(n2184) );
  INVX0 U2253 ( .ZN(n7327), .INP(n2181) );
  INVX0 U2252 ( .ZN(n7326), .INP(n4184) );
  INVX0 U2148 ( .ZN(n7222), .INP(P2_N5099) );
  INVX0 U2043 ( .ZN(n7117), .INP(P1_N5177) );
  INVX0 U2254 ( .ZN(n7328), .INP(n4181) );
  NBUFFX4 U2163 ( .Z(n7237), .INP(P2_N5096) );
  INVX0 U2192 ( .ZN(n7266), .INP(P2_N5100) );
  INVX0 U2072 ( .ZN(n7146), .INP(P1_N5178) );
  INVX0 U395 ( .ZN(n6592), .INP(n18207) );
  INVX0 U434 ( .ZN(n6620), .INP(n18285) );
  INVX0 U433 ( .ZN(n6619), .INP(n18287) );
  INVX0 U396 ( .ZN(n6593), .INP(n18205) );
  INVX0 U2197 ( .ZN(n7271), .INP(P1_N536) );
  INVX0 U2198 ( .ZN(n7272), .INP(P2_N536) );
  NBUFFX4 U1821 ( .Z(n6895), .INP(n7483) );
  INVX0 U1925 ( .ZN(n6999), .INP(P2_N584) );
  NBUFFX4 U1763 ( .Z(n6837), .INP(n7485) );
  INVX0 U1822 ( .ZN(n6896), .INP(n6895) );
  INVX0 U1764 ( .ZN(n6838), .INP(n6837) );
  INVX2 U1836 ( .INP(n7483), .ZN(n6910) );
  NAND2X1 U1855 ( .IN2(n6332), .IN1(n6333), .QN(n7458) );
  INVX0 U1922 ( .ZN(n6996), .INP(P1_N584) );
  NBUFFX4 U1773 ( .Z(n6847), .INP(n7484) );
  NBUFFX4 U1795 ( .Z(n6869), .INP(n7458) );
  NBUFFX4 U1735 ( .Z(n6809), .INP(n7484) );
  NBUFFX4 U1819 ( .Z(n6893), .INP(n7482) );
  NBUFFX4 U1823 ( .Z(n6897), .INP(n7482) );
  NBUFFX4 U1825 ( .Z(n6899), .INP(n7482) );
  INVX0 U1774 ( .ZN(n6848), .INP(n6847) );
  NBUFFX4 U1841 ( .Z(n6915), .INP(n7482) );
  INVX0 U1796 ( .ZN(n6870), .INP(n6869) );
  INVX0 U1734 ( .ZN(n6808), .INP(n6807) );
  INVX0 U1780 ( .ZN(n6854), .INP(n7459) );
  NBUFFX4 U1809 ( .Z(n6883), .INP(n7482) );
  INVX0 U1824 ( .ZN(n6898), .INP(n6897) );
  INVX0 U1826 ( .ZN(n6900), .INP(n6899) );
  INVX0 U1842 ( .ZN(n6916), .INP(n6915) );
  NBUFFX4 U1843 ( .Z(n6917), .INP(n7482) );
  NBUFFX4 U1745 ( .Z(n6819), .INP(n7485) );
  AND2X1 U4028 ( .IN1(n2992), .IN2(n7354), .Q(n2934) );
  NOR2X2 U8377 ( .QN(n5709), .IN1(n7356), .IN2(n7355) );
  NOR2X2 U5855 ( .QN(n4022), .IN1(n7376), .IN2(n7375) );
  NOR2X1 U5624 ( .QN(n3796), .IN1(n7378), .IN2(n7377) );
  NOR2X1 U5330 ( .QN(n3710), .IN1(n7380), .IN2(n7379) );
  NOR2X1 U5179 ( .QN(n3624), .IN1(n7382), .IN2(n7381) );
  NOR2X1 U5001 ( .QN(n3512), .IN1(n7384), .IN2(n7383) );
  NOR2X1 U4826 ( .QN(n3403), .IN1(n7386), .IN2(n7385) );
  NOR2X1 U4656 ( .QN(n3299), .IN1(n7388), .IN2(n7387) );
  NOR2X1 U4505 ( .QN(n3213), .IN1(n7390), .IN2(n7389) );
  NOR2X1 U4331 ( .QN(n3105), .IN1(n7392), .IN2(n7391) );
  NOR2X1 U4180 ( .QN(n3019), .IN1(n7394), .IN2(n7393) );
  NOR2X1 U2875 ( .QN(n2069), .IN1(n7395), .IN2(n7396) );
  NAND2X1 U1514 ( .IN2(P2_N4244), .IN1(n1466), .QN(P2_N5509) );
  OR2X2 U1551 ( .IN2(n1485), .IN1(P1_N3434), .Q(P1_N5581) );
  NBUFFX4 U1817 ( .Z(n6891), .INP(P1_N292) );
  NBUFFX4 U1875 ( .Z(n6949), .INP(P1_N293) );
  NBUFFX4 U1777 ( .Z(n6851), .INP(P2_N292) );
  NBUFFX4 U1761 ( .Z(n6835), .INP(P2_N292) );
  INVX0 U1760 ( .ZN(n6834), .INP(n7484) );
  NBUFFX4 U1741 ( .Z(n6815), .INP(n7486) );
  INVX0 U432 ( .ZN(n6618), .INP(P1_N506) );
  INVX0 U394 ( .ZN(n6591), .INP(P2_N506) );
  INVX0 P1_I_289 ( .ZN(P1_N3062), .INP(P1_N2878) );
  INVX0 P1_I_290 ( .ZN(P1_N3031), .INP(P1_N2880) );
  INVX0 P1_I_324 ( .ZN(P1_N3435), .INP(P1_N3251) );
  INVX0 P1_I_325 ( .ZN(P1_N3404), .INP(P1_N3253) );
  INVX0 P1_I_359 ( .ZN(P1_N3808), .INP(P1_N3624) );
  INVX0 P1_I_360 ( .ZN(P1_N3777), .INP(P1_N3626) );
  INVX0 P1_I_394 ( .ZN(P1_N4181), .INP(P1_N3997) );
  INVX0 P1_I_395 ( .ZN(P1_N4150), .INP(P1_N3999) );
  INVX0 P1_I_429 ( .ZN(P1_N4554), .INP(P1_N4370) );
  INVX0 P1_I_430 ( .ZN(P1_N4523), .INP(P1_N4372) );
  INVX0 P1_I_472 ( .ZN(P1_N6685), .INP(P1_N5137) );
  INVX0 P1_I_473 ( .ZN(P1_N6686), .INP(P1_N5140) );
  INVX0 P1_I_477 ( .ZN(P1_N6688), .INP(P1_N5431) );
  INVX0 P1_I_79 ( .ZN(P1_N969), .INP(P1_N779) );
  INVX0 P1_I_80 ( .ZN(P1_N938), .INP(P1_N781) );
  INVX0 P1_I_114 ( .ZN(P1_N1315), .INP(P1_N1250) );
  INVX0 P1_I_115 ( .ZN(P1_N1284), .INP(P1_N1252) );
  INVX0 P1_I_184 ( .ZN(P1_N1943), .INP(P1_N1759) );
  INVX0 P1_I_185 ( .ZN(P1_N1912), .INP(P1_N1761) );
  INVX0 P1_I_219 ( .ZN(P1_N2316), .INP(P1_N2132) );
  INVX0 P1_I_220 ( .ZN(P1_N2285), .INP(P1_N2134) );
  INVX0 P1_I_254 ( .ZN(P1_N2689), .INP(P1_N2505) );
  INVX0 P1_I_255 ( .ZN(P1_N2658), .INP(P1_N2507) );
  INVX0 P2_I_477 ( .ZN(P2_N6610), .INP(P2_N5353) );
  INVX0 P2_I_184 ( .ZN(P2_N1817), .INP(P2_N1633) );
  INVX0 P2_I_185 ( .ZN(P2_N1786), .INP(P2_N1635) );
  INVX0 P2_I_219 ( .ZN(P2_N2190), .INP(P2_N2006) );
  INVX0 P2_I_220 ( .ZN(P2_N2159), .INP(P2_N2008) );
  INVX0 P2_I_254 ( .ZN(P2_N2563), .INP(P2_N2379) );
  INVX0 P2_I_255 ( .ZN(P2_N2532), .INP(P2_N2381) );
  INVX0 P2_I_289 ( .ZN(P2_N2936), .INP(P2_N2752) );
  INVX0 P2_I_290 ( .ZN(P2_N2905), .INP(P2_N2754) );
  INVX0 P2_I_324 ( .ZN(P2_N3309), .INP(P2_N3125) );
  INVX0 P2_I_325 ( .ZN(P2_N3278), .INP(P2_N3127) );
  INVX0 P2_I_359 ( .ZN(P2_N3682), .INP(P2_N3498) );
  INVX0 P2_I_360 ( .ZN(P2_N3651), .INP(P2_N3500) );
  INVX0 P2_I_394 ( .ZN(P2_N4055), .INP(P2_N3871) );
  INVX0 P2_I_395 ( .ZN(P2_N4024), .INP(P2_N3873) );
  INVX0 P2_I_429 ( .ZN(P2_N4428), .INP(P2_N4244) );
  INVX0 P2_I_472 ( .ZN(P2_N6607), .INP(P2_N5059) );
  INVX0 P2_I_473 ( .ZN(P2_N6608), .INP(P2_N5062) );
  INVX0 U1866 ( .ZN(n6940), .INP(n7460) );
  INVX0 P2_I_79 ( .ZN(P2_N843), .INP(P2_N778) );
  INVX0 P2_I_80 ( .ZN(P2_N812), .INP(P2_N780) );
  INVX0 P2_I_114 ( .ZN(P2_N1189), .INP(P2_N1124) );
  INVX0 P2_I_115 ( .ZN(P2_N1158), .INP(P2_N1126) );
  NBUFFX4 U1905 ( .Z(n6979), .INP(P1_N294) );
  INVX0 U1750 ( .ZN(n6824), .INP(n6823) );
  NBUFFX4 U1769 ( .Z(n6843), .INP(P2_N292) );
  NBUFFX4 U1707 ( .Z(n6781), .INP(P2_N291) );
  NBUFFX2 U1755 ( .Z(n6829), .INP(n7486) );
  NOR2X1 U6486 ( .QN(n4510), .IN1(n7400), .IN2(n7399) );
  INVX0 P1_I_471 ( .ZN(P1_N5282), .INP(P1_N5281) );
  INVX0 P1_I_149 ( .ZN(P1_N1570), .INP(P1_N1505) );
  INVX0 P1_I_150 ( .ZN(P1_N1539), .INP(P1_N1507) );
  INVX0 P2_I_471 ( .ZN(P2_N5204), .INP(P2_N5203) );
  INVX0 P2_I_149 ( .ZN(P2_N1444), .INP(P2_N1379) );
  INVX0 P2_I_150 ( .ZN(P2_N1413), .INP(P2_N1381) );
  INVX2 U1906 ( .INP(n6979), .ZN(n6980) );
  INVX0 U1898 ( .ZN(n6972), .INP(P2_N294) );
  INVX0 U1728 ( .ZN(n6802), .INP(P2_N291) );
  INVX0 U1786 ( .ZN(n6860), .INP(n7458) );
  NBUFFX8 U1781 ( .Z(n6855), .INP(P1_N291) );
  INVX0 U18978 ( .ZN(n14763), .INP(n14523) );
  INVX0 U15651 ( .ZN(n11550), .INP(n11310) );
  INVX0 P1_I_464 ( .ZN(P1_N4817), .INP(P1_N4752) );
  INVX0 P1_I_465 ( .ZN(P1_N4786), .INP(P1_N4754) );
  INVX0 P2_I_464 ( .ZN(P2_N4691), .INP(P2_N4626) );
  INVX0 U1860 ( .ZN(n6934), .INP(n7460) );
  NBUFFX4 U1901 ( .Z(n6975), .INP(P1_N294) );
  INVX0 U1880 ( .ZN(n6954), .INP(n7461) );
  NBUFFX4 U1903 ( .Z(n6977), .INP(P1_N294) );
  INVX0 U1892 ( .ZN(n6966), .INP(P2_N294) );
  INVX0 U1910 ( .ZN(n6984), .INP(P1_N294) );
  INVX0 U386 ( .ZN(n6584), .INP(n6583) );
  NOR2X0 U3280 ( .QN(n2168), .IN1(n6589), .IN2(P2_N499) );
  NOR2X0 U6158 ( .QN(n4164), .IN1(n6583), .IN2(n4356) );
  NBUFFX4 U387 ( .Z(n6585), .INP(n2166) );
  NOR2X0 U6164 ( .QN(n4171), .IN1(n6583), .IN2(P1_N499) );
  INVX0 U384 ( .ZN(n6582), .INP(n4169) );
  INVX0 U388 ( .ZN(n6586), .INP(n6585) );
  NBUFFX2 U2004 ( .Z(n7455), .INP(n7449) );
  NBUFFX4 U1975 ( .Z(n7448), .INP(n7456) );
  NOR2X1 U304 ( .QN(n598), .IN1(n2459), .IN2(n6589) );
  NOR2X1 U306 ( .QN(n599), .IN1(n2452), .IN2(n6589) );
  NOR2X1 U157 ( .QN(n480), .IN1(n4366), .IN2(n6583) );
  NOR2X1 U159 ( .QN(n481), .IN1(n4356), .IN2(n6583) );
  NBUFFX2 U381 ( .Z(n6579), .INP(n7455) );
  NBUFFX2 U371 ( .Z(n6570), .INP(n7448) );
  INVX0 U2211 ( .ZN(n7285), .INP(P2_N5419) );
  INVX2 U1957 ( .INP(P1_N5554), .ZN(n7031) );
  INVX0 U2210 ( .ZN(n7284), .INP(P1_N5497) );
  NBUFFX2 U374 ( .Z(n6572), .INP(n7457) );
  NBUFFX2 U369 ( .Z(n6568), .INP(n7455) );
  NBUFFX2 U379 ( .Z(n6577), .INP(n7540) );
  NBUFFX2 U380 ( .Z(n6578), .INP(n7454) );
  NBUFFX2 U2054 ( .Z(n7478), .INP(n7539) );
  NBUFFX2 U378 ( .Z(n6576), .INP(n7454) );
  NBUFFX2 U375 ( .Z(n6573), .INP(n7457) );
  NBUFFX2 U2161 ( .Z(n7536), .INP(n7454) );
  NBUFFX2 U2159 ( .Z(n7535), .INP(n7455) );
  NBUFFX2 U2181 ( .Z(n7549), .INP(n7540) );
  NBUFFX2 U2182 ( .Z(n7553), .INP(n7540) );
  NBUFFX2 U2183 ( .Z(n7554), .INP(n7540) );
  NBUFFX2 U2184 ( .Z(n7555), .INP(n7540) );
  NBUFFX2 U370 ( .Z(n6569), .INP(n7454) );
  NBUFFX2 U376 ( .Z(n6574), .INP(n7457) );
  NBUFFX2 U2233 ( .Z(n7584), .INP(n7539) );
  NBUFFX2 U2230 ( .Z(n7581), .INP(n7539) );
  NBUFFX2 U2231 ( .Z(n7582), .INP(n7539) );
  NBUFFX2 U2234 ( .Z(n7585), .INP(n7454) );
  NBUFFX2 U2256 ( .Z(n7586), .INP(n7454) );
  NBUFFX2 U2232 ( .Z(n7583), .INP(n7539) );
  NBUFFX2 U2098 ( .Z(n7505), .INP(n7457) );
  NBUFFX2 U2097 ( .Z(n7504), .INP(n7457) );
  NBUFFX2 U2101 ( .Z(n7506), .INP(n7457) );
  NBUFFX4 U2057 ( .Z(n7480), .INP(n19009) );
  NBUFFX4 U1639 ( .Z(n6713), .INP(n7480) );
  NBUFFX8 U1713 ( .Z(n6787), .INP(n7487) );
  NBUFFX4 U1869 ( .Z(n6943), .INP(n7460) );
  INVX0 U1858 ( .ZN(n6932), .INP(n6931) );
  NBUFFX8 U1863 ( .Z(n6937), .INP(P2_N293) );
  INVX2 U1872 ( .INP(P2_N293), .ZN(n6946) );
  NBUFFX4 U2003 ( .Z(n7454), .INP(Scan_Enable) );
  INVX0 U2276 ( .ZN(n7606), .INP(reset) );
  INVX0 U2275 ( .ZN(n7605), .INP(reset) );
  INVX0 U2274 ( .ZN(n7604), .INP(reset) );
  INVX0 U2273 ( .ZN(n7603), .INP(reset) );
  INVX0 U2272 ( .ZN(n7602), .INP(reset) );
  INVX0 U2271 ( .ZN(n7601), .INP(reset) );
  NBUFFX2 U2270 ( .Z(n7600), .INP(n6577) );
  NBUFFX2 U2269 ( .Z(n7599), .INP(n6577) );
  NBUFFX2 U2268 ( .Z(n7598), .INP(n6577) );
  NBUFFX2 U2267 ( .Z(n7597), .INP(n6577) );
  NBUFFX2 U2266 ( .Z(n7596), .INP(n6577) );
  NBUFFX2 U2265 ( .Z(n7595), .INP(n6577) );
  INVX0 U2264 ( .ZN(n7594), .INP(reset) );
  INVX0 U2263 ( .ZN(n7593), .INP(reset) );
  INVX0 U2262 ( .ZN(n7592), .INP(reset) );
  INVX0 U2261 ( .ZN(n7591), .INP(reset) );
  INVX0 U2260 ( .ZN(n7590), .INP(reset) );
  INVX0 U2259 ( .ZN(n7589), .INP(reset) );
  INVX0 U2258 ( .ZN(n7588), .INP(reset) );
  NBUFFX4 U2257 ( .Z(n7587), .INP(n7539) );
  INVX0 U2228 ( .ZN(n7580), .INP(reset) );
  INVX0 U2227 ( .ZN(n7579), .INP(reset) );
  INVX0 U2226 ( .ZN(n7578), .INP(reset) );
  INVX0 U2224 ( .ZN(n7577), .INP(reset) );
  INVX0 U2223 ( .ZN(n7576), .INP(reset) );
  INVX0 U2222 ( .ZN(n7575), .INP(reset) );
  INVX0 U2220 ( .ZN(n7574), .INP(reset) );
  NBUFFX2 U2219 ( .Z(n7573), .INP(n6571) );
  NBUFFX2 U2218 ( .Z(n7572), .INP(n6571) );
  NBUFFX2 U2216 ( .Z(n7571), .INP(n7453) );
  NBUFFX2 U2215 ( .Z(n7570), .INP(n7453) );
  NBUFFX2 U2214 ( .Z(n7569), .INP(n6571) );
  NBUFFX2 U2212 ( .Z(n7568), .INP(n6571) );
  NBUFFX2 U2209 ( .Z(n7567), .INP(n6571) );
  NBUFFX2 U2208 ( .Z(n7566), .INP(n7453) );
  NBUFFX2 U2206 ( .Z(n7565), .INP(n6571) );
  INVX0 U2204 ( .ZN(n7564), .INP(reset) );
  INVX0 U2203 ( .ZN(n7563), .INP(reset) );
  INVX0 U2202 ( .ZN(n7562), .INP(reset) );
  INVX0 U2195 ( .ZN(n7561), .INP(reset) );
  INVX0 U2194 ( .ZN(n7560), .INP(reset) );
  INVX0 U2193 ( .ZN(n7559), .INP(reset) );
  INVX0 U2188 ( .ZN(n7558), .INP(reset) );
  INVX0 U2187 ( .ZN(n7557), .INP(reset) );
  INVX0 U2180 ( .ZN(n7548), .INP(reset) );
  INVX0 U2177 ( .ZN(n7547), .INP(reset) );
  INVX0 U2176 ( .ZN(n7546), .INP(reset) );
  INVX0 U2175 ( .ZN(n7545), .INP(reset) );
  INVX0 U2172 ( .ZN(n7544), .INP(reset) );
  INVX0 U2171 ( .ZN(n7543), .INP(reset) );
  INVX0 U2170 ( .ZN(n7542), .INP(reset) );
  INVX0 U2167 ( .ZN(n7541), .INP(reset) );
  NBUFFX2 U2166 ( .Z(n7538), .INP(n6560) );
  NBUFFX2 U2162 ( .Z(n7537), .INP(n6560) );
  INVX0 U2158 ( .ZN(n7534), .INP(reset) );
  INVX0 U2156 ( .ZN(n7533), .INP(reset) );
  INVX0 U2154 ( .ZN(n7532), .INP(reset) );
  INVX0 U2152 ( .ZN(n7531), .INP(reset) );
  NBUFFX4 U2151 ( .Z(n7530), .INP(n6568) );
  NBUFFX2 U2149 ( .Z(n7529), .INP(n6568) );
  NBUFFX2 U2147 ( .Z(n7528), .INP(n6568) );
  NBUFFX2 U2144 ( .Z(n7527), .INP(n6568) );
  NBUFFX2 U2143 ( .Z(n7526), .INP(n6568) );
  NBUFFX2 U2141 ( .Z(n7525), .INP(n6568) );
  NBUFFX4 U2139 ( .Z(n7524), .INP(n6556) );
  NBUFFX2 U2138 ( .Z(n7523), .INP(n6556) );
  NBUFFX2 U2133 ( .Z(n7522), .INP(n6556) );
  NBUFFX2 U2130 ( .Z(n7521), .INP(n6556) );
  NBUFFX2 U2129 ( .Z(n7520), .INP(n6556) );
  NBUFFX2 U2126 ( .Z(n7519), .INP(n6556) );
  NBUFFX2 U2125 ( .Z(n7518), .INP(n6579) );
  NBUFFX2 U2122 ( .Z(n7517), .INP(n6579) );
  NBUFFX2 U2119 ( .Z(n7516), .INP(n6579) );
  NBUFFX2 U2118 ( .Z(n7515), .INP(n6579) );
  NBUFFX2 U2117 ( .Z(n7514), .INP(n6579) );
  NBUFFX2 U2116 ( .Z(n7513), .INP(n6579) );
  NBUFFX4 U2115 ( .Z(n7512), .INP(n6567) );
  NBUFFX2 U2111 ( .Z(n7511), .INP(n6567) );
  NBUFFX2 U2109 ( .Z(n7510), .INP(n6567) );
  NBUFFX2 U2106 ( .Z(n7509), .INP(n6567) );
  NBUFFX2 U2105 ( .Z(n7508), .INP(n6567) );
  NBUFFX2 U2102 ( .Z(n7507), .INP(n6567) );
  NBUFFX4 U2096 ( .Z(n7502), .INP(n6561) );
  NBUFFX2 U2095 ( .Z(n7501), .INP(n6561) );
  NBUFFX2 U2094 ( .Z(n7500), .INP(n6561) );
  NBUFFX2 U2093 ( .Z(n7499), .INP(n6561) );
  NBUFFX2 U2089 ( .Z(n7498), .INP(n6561) );
  NBUFFX2 U2087 ( .Z(n7497), .INP(n6561) );
  NBUFFX2 U2086 ( .Z(n7496), .INP(n6570) );
  NBUFFX2 U2085 ( .Z(n7495), .INP(n6570) );
  NBUFFX2 U2082 ( .Z(n7494), .INP(n7448) );
  NBUFFX2 U2081 ( .Z(n7493), .INP(n7448) );
  NBUFFX2 U2078 ( .Z(n7492), .INP(n6570) );
  NBUFFX2 U2076 ( .Z(n7491), .INP(n6570) );
  NBUFFX2 U2074 ( .Z(n7490), .INP(n6570) );
  NBUFFX2 U2069 ( .Z(n7489), .INP(n6570) );
  NAND2X1 U2068 ( .IN2(n6382), .IN1(n6383), .QN(n7488) );
  NAND2X1 U2066 ( .IN2(n6382), .IN1(n6383), .QN(n7487) );
  NAND2X1 U2065 ( .IN2(n6384), .IN1(n6385), .QN(n7486) );
  NAND2X1 U2063 ( .IN2(n6384), .IN1(n6385), .QN(n7485) );
  NAND2X1 U2061 ( .IN2(n6384), .IN1(n6385), .QN(n7484) );
  NAND2X1 U2060 ( .IN2(n6334), .IN1(n6335), .QN(n7483) );
  NAND2X1 U2059 ( .IN2(n6334), .IN1(n6335), .QN(n7482) );
  NAND2X1 U2058 ( .IN2(n6334), .IN1(n6335), .QN(n7481) );
  NBUFFX2 U2053 ( .Z(n7477), .INP(n6566) );
  NBUFFX2 U2052 ( .Z(n7476), .INP(n6566) );
  NBUFFX4 U2049 ( .Z(n7475), .INP(n6575) );
  NBUFFX2 U2047 ( .Z(n7474), .INP(n6575) );
  NBUFFX2 U2046 ( .Z(n7473), .INP(n6575) );
  NBUFFX2 U2044 ( .Z(n7472), .INP(n6575) );
  NBUFFX4 U2040 ( .Z(n7471), .INP(n6563) );
  NBUFFX2 U2037 ( .Z(n7470), .INP(n6563) );
  NBUFFX2 U2034 ( .Z(n7469), .INP(n6563) );
  NBUFFX2 U2033 ( .Z(n7468), .INP(n6563) );
  NBUFFX2 U2030 ( .Z(n7467), .INP(n6572) );
  NBUFFX2 U2027 ( .Z(n7466), .INP(n6572) );
  NBUFFX2 U2026 ( .Z(n7465), .INP(n6572) );
  NBUFFX2 U2023 ( .Z(n7464), .INP(n6572) );
  NAND2X1 U2020 ( .IN2(P1_N584), .IN1(n1502), .QN(n7463) );
  NAND2X1 U2017 ( .IN2(P2_N584), .IN1(n1481), .QN(n7462) );
  NAND2X1 U2014 ( .IN2(n6338), .IN1(n6339), .QN(n7461) );
  NAND2X1 U2013 ( .IN2(n6388), .IN1(n6389), .QN(n7460) );
  NAND2X1 U2012 ( .IN2(n6332), .IN1(n6333), .QN(n7459) );
  NBUFFX2 U2011 ( .Z(n7540), .INP(Scan_Enable) );
  NBUFFX4 U2010 ( .Z(n7457), .INP(n7449) );
  NBUFFX4 U2009 ( .Z(n7539), .INP(n7449) );
  NBUFFX2 U2000 ( .Z(n7550), .INP(n7540) );
  NBUFFX2 U1995 ( .Z(n7452), .INP(n7550) );
  NBUFFX2 U1994 ( .Z(n7451), .INP(n7518) );
  NBUFFX2 U1991 ( .Z(n7450), .INP(n7492) );
  NBUFFX2 U1990 ( .Z(n7556), .INP(n7456) );
  NBUFFX2 U1987 ( .Z(n7503), .INP(n7456) );
  NBUFFX2 U1986 ( .Z(n7453), .INP(n7456) );
  NBUFFX4 U1983 ( .Z(n7449), .INP(Scan_Enable) );
  NBUFFX2 U1980 ( .Z(n7456), .INP(n7449) );
  NBUFFX2 U1979 ( .Z(n7552), .INP(n7448) );
  NBUFFX2 U1976 ( .Z(n7551), .INP(n7448) );
  AND2X1 U1973 ( .IN1(n2586), .IN2(n2587), .Q(n7447) );
  AND2X1 U1970 ( .IN1(n2579), .IN2(n2580), .Q(n7446) );
  NAND2X1 U1968 ( .IN2(n4499), .IN1(n4498), .QN(n7445) );
  NAND2X1 U1966 ( .IN2(n4491), .IN1(n4490), .QN(n7444) );
  AND2X1 U1965 ( .IN1(P1_N5433), .IN2(n4367), .Q(n7443) );
  AND2X1 U1964 ( .IN1(P2_N5355), .IN2(n2460), .Q(n7442) );
  AND2X1 U1959 ( .IN1(n4171), .IN2(P1_N663), .Q(n7441) );
  AND2X1 U1958 ( .IN1(n4171), .IN2(P1_N664), .Q(n7440) );
  AND2X1 U1956 ( .IN1(n4171), .IN2(P1_N666), .Q(n7439) );
  AND2X1 U1951 ( .IN1(n4171), .IN2(P1_N668), .Q(n7438) );
  AND2X1 U1946 ( .IN1(n4171), .IN2(P1_N669), .Q(n7437) );
  AND2X1 U1944 ( .IN1(n4171), .IN2(P1_N670), .Q(n7436) );
  AND2X1 U1943 ( .IN1(n4171), .IN2(P1_N671), .Q(n7435) );
  AND2X1 U1940 ( .IN1(n4171), .IN2(P1_N672), .Q(n7434) );
  AND2X1 U1931 ( .IN1(n4171), .IN2(P1_N673), .Q(n7433) );
  AND2X1 U1930 ( .IN1(n4171), .IN2(P1_N674), .Q(n7432) );
  AND2X1 U1929 ( .IN1(n4171), .IN2(P1_N675), .Q(n7431) );
  AND2X1 U1928 ( .IN1(n4171), .IN2(P1_N676), .Q(n7430) );
  AND2X1 U1927 ( .IN1(n4171), .IN2(P1_N677), .Q(n7429) );
  AND2X1 U1926 ( .IN1(n4171), .IN2(P1_N678), .Q(n7428) );
  AND2X1 U1924 ( .IN1(n4171), .IN2(P1_N679), .Q(n7427) );
  AND2X1 U1923 ( .IN1(n4171), .IN2(P1_N680), .Q(n7426) );
  AND2X1 U1921 ( .IN1(n4171), .IN2(P1_N681), .Q(n7425) );
  AND2X1 U1920 ( .IN1(n4171), .IN2(P1_N682), .Q(n7424) );
  AND2X1 U1917 ( .IN1(n7422), .IN2(n7409), .Q(n7423) );
  NOR2X0 U1916 ( .QN(n7422), .IN1(n6837), .IN2(n6784) );
  NAND2X1 U1915 ( .IN2(n7412), .IN1(n7411), .QN(n7421) );
  AND2X1 U1914 ( .IN1(n7413), .IN2(n7409), .Q(n7420) );
  NAND2X1 U1913 ( .IN2(n7408), .IN1(n7407), .QN(n7419) );
  AND2X1 U1911 ( .IN1(n7410), .IN2(n7409), .Q(n7418) );
  AND2X1 U1909 ( .IN1(n7406), .IN2(n7405), .Q(n7417) );
  AND2X1 U1904 ( .IN1(n7404), .IN2(n7405), .Q(n7416) );
  NAND2X1 U1897 ( .IN2(P2_N245), .IN1(n6381), .QN(n7415) );
  NAND2X1 U1894 ( .IN2(P1_N245), .IN1(n6331), .QN(n7414) );
  NOR2X0 U1891 ( .QN(n7413), .IN1(n6838), .IN2(n6784) );
  NOR2X0 U1890 ( .QN(n7412), .IN1(n6837), .IN2(n6793) );
  NOR2X0 U1879 ( .QN(n7411), .IN1(n6972), .IN2(n6940) );
  NOR2X0 U1877 ( .QN(n7410), .IN1(n6838), .IN2(n6793) );
  NOR2X0 U1876 ( .QN(n7409), .IN1(n6963), .IN2(n6931) );
  NOR2X0 U1873 ( .QN(n7408), .IN1(n6883), .IN2(n6857) );
  NOR2X0 U1871 ( .QN(n7407), .IN1(n6980), .IN2(n6956) );
  NOR2X0 U1862 ( .QN(n7406), .IN1(n6896), .IN2(n6870) );
  NOR2X0 U1861 ( .QN(n7405), .IN1(n6979), .IN2(n6949) );
  NOR2X0 U1859 ( .QN(n7404), .IN1(n6896), .IN2(n6869) );
  NOR2X0 U1856 ( .QN(n7403), .IN1(P1_N5755), .IN2(P1_N5756) );
  AND2X1 U1851 ( .IN1(n7398), .IN2(P2_N4561), .Q(n7402) );
  NOR2X0 U1850 ( .QN(n7401), .IN1(P2_N5677), .IN2(P2_N5678) );
  NOR2X0 U1844 ( .QN(n7400), .IN1(P1_N6683), .IN2(P1_N6684) );
  NOR2X0 U1840 ( .QN(n7399), .IN1(P1_N6681), .IN2(P1_N6682) );
  NOR2X0 U1839 ( .QN(n7398), .IN1(P2_N6605), .IN2(P2_N6606) );
  AND2X1 U1838 ( .IN1(n7354), .IN2(P2_N4178), .Q(n7397) );
  NOR2X0 U1837 ( .QN(n7396), .IN1(P2_N5899), .IN2(P2_N5900) );
  NOR2X0 U1835 ( .QN(n7395), .IN1(P2_N5901), .IN2(P2_N5902) );
  NOR2X0 U1834 ( .QN(n7394), .IN1(P2_N6477), .IN2(P2_N6478) );
  NOR2X0 U1831 ( .QN(n7393), .IN1(P2_N6475), .IN2(P2_N6476) );
  NOR2X0 U1829 ( .QN(n7392), .IN1(P2_N6413), .IN2(P2_N6414) );
  NOR2X0 U1828 ( .QN(n7391), .IN1(P2_N6411), .IN2(P2_N6412) );
  NOR2X0 U1815 ( .QN(n7390), .IN1(P2_N6349), .IN2(P2_N6350) );
  NOR2X0 U1811 ( .QN(n7389), .IN1(P2_N6347), .IN2(P2_N6348) );
  NOR2X0 U1806 ( .QN(n7388), .IN1(P2_N6285), .IN2(P2_N6286) );
  NOR2X0 U1805 ( .QN(n7387), .IN1(P2_N6283), .IN2(P2_N6284) );
  NOR2X0 U1803 ( .QN(n7386), .IN1(P2_N6221), .IN2(P2_N6222) );
  NOR2X0 U1802 ( .QN(n7385), .IN1(P2_N6219), .IN2(P2_N6220) );
  NOR2X0 U1801 ( .QN(n7384), .IN1(P2_N6157), .IN2(P2_N6158) );
  NOR2X0 U1799 ( .QN(n7383), .IN1(P2_N6155), .IN2(P2_N6156) );
  NOR2X0 U1789 ( .QN(n7382), .IN1(P2_N6093), .IN2(P2_N6094) );
  NOR2X0 U1785 ( .QN(n7381), .IN1(P2_N6091), .IN2(P2_N6092) );
  NOR2X0 U1784 ( .QN(n7380), .IN1(P2_N6029), .IN2(P2_N6030) );
  NOR2X0 U1779 ( .QN(n7379), .IN1(P2_N6027), .IN2(P2_N6028) );
  NOR2X0 U1776 ( .QN(n7378), .IN1(P2_N5965), .IN2(P2_N5966) );
  NOR2X0 U1775 ( .QN(n7377), .IN1(P2_N5963), .IN2(P2_N5964) );
  NOR2X0 U1772 ( .QN(n7376), .IN1(P1_N5979), .IN2(P1_N5980) );
  NOR2X0 U1771 ( .QN(n7375), .IN1(P1_N5977), .IN2(P1_N5978) );
  NOR2X0 U1770 ( .QN(n7374), .IN1(P1_N6619), .IN2(P1_N6620) );
  NOR2X0 U1767 ( .QN(n7373), .IN1(P1_N6617), .IN2(P1_N6618) );
  NOR2X0 U1766 ( .QN(n7372), .IN1(P1_N6555), .IN2(P1_N6556) );
  NOR2X0 U1765 ( .QN(n7371), .IN1(P1_N6553), .IN2(P1_N6554) );
  NOR2X0 U1759 ( .QN(n7370), .IN1(P1_N6491), .IN2(P1_N6492) );
  NOR2X0 U1752 ( .QN(n7369), .IN1(P1_N6489), .IN2(P1_N6490) );
  NOR2X0 U1747 ( .QN(n7368), .IN1(P1_N6427), .IN2(P1_N6428) );
  NOR2X0 U1743 ( .QN(n7367), .IN1(P1_N6425), .IN2(P1_N6426) );
  NOR2X0 U1740 ( .QN(n7366), .IN1(P1_N6363), .IN2(P1_N6364) );
  NOR2X0 U1737 ( .QN(n7365), .IN1(P1_N6361), .IN2(P1_N6362) );
  NOR2X0 U1732 ( .QN(n7364), .IN1(P1_N6299), .IN2(P1_N6300) );
  NOR2X0 U1731 ( .QN(n7363), .IN1(P1_N6297), .IN2(P1_N6298) );
  NOR2X0 U1727 ( .QN(n7362), .IN1(P1_N6235), .IN2(P1_N6236) );
  NOR2X0 U1726 ( .QN(n7361), .IN1(P1_N6233), .IN2(P1_N6234) );
  NOR2X0 U1725 ( .QN(n7360), .IN1(P1_N6171), .IN2(P1_N6172) );
  NOR2X0 U1723 ( .QN(n7359), .IN1(P1_N6169), .IN2(P1_N6170) );
  NOR2X0 U1722 ( .QN(n7358), .IN1(P1_N6107), .IN2(P1_N6108) );
  NOR2X0 U1721 ( .QN(n7357), .IN1(P1_N6105), .IN2(P1_N6106) );
  NOR2X0 U1714 ( .QN(n7356), .IN1(P1_N6043), .IN2(P1_N6044) );
  NOR2X0 U1711 ( .QN(n7355), .IN1(P1_N6041), .IN2(P1_N6042) );
  NOR2X0 U1709 ( .QN(n7354), .IN1(P2_N6541), .IN2(P2_N6542) );
  NOR2X0 U1704 ( .QN(n7353), .IN1(P2_N5631), .IN2(P2_N5632) );
  NOR2X0 U1703 ( .QN(n7352), .IN1(P1_N5709), .IN2(P1_N5710) );
  NOR2X0 U1664 ( .QN(n7351), .IN1(P1_N5653), .IN2(P1_N5654) );
  NOR2X0 U1654 ( .QN(n7350), .IN1(P2_N5575), .IN2(P2_N5576) );
  AND2X1 U1653 ( .IN1(n9310), .IN2(n4480), .Q(n7349) );
  AND2X1 U1652 ( .IN1(n9314), .IN2(n4480), .Q(n7348) );
  AND2X1 U1650 ( .IN1(n4615), .IN2(n4616), .Q(n7347) );
  AND2X1 U1649 ( .IN1(n2660), .IN2(n2661), .Q(n7346) );
  AND2X1 U1648 ( .IN1(n7336), .IN2(n4616), .Q(n7345) );
  AND2X1 U1635 ( .IN1(n7335), .IN2(n4615), .Q(n7344) );
  AND2X1 U1633 ( .IN1(n7339), .IN2(n2661), .Q(n7343) );
  AND2X1 U1627 ( .IN1(n7338), .IN2(n2660), .Q(n7342) );
  AND2X1 U1623 ( .IN1(n2153), .IN2(n2154), .Q(n7341) );
  AND2X1 U1621 ( .IN1(n4157), .IN2(n4158), .Q(n7340) );
  AND2X1 U1617 ( .IN1(n6415), .IN2(n6414), .Q(n7339) );
  AND2X1 U1615 ( .IN1(n6418), .IN2(n6417), .Q(n7338) );
  AND2X1 U1573 ( .IN1(n7331), .IN2(n4158), .Q(n7337) );
  AND2X1 U1569 ( .IN1(n6365), .IN2(n6364), .Q(n7336) );
  AND2X1 U1542 ( .IN1(n6368), .IN2(n6367), .Q(n7335) );
  AND2X1 U1538 ( .IN1(n7333), .IN2(n2154), .Q(n7334) );
  AND2X1 U389 ( .IN1(n6401), .IN2(n6400), .Q(n7333) );
  AND2X1 U383 ( .IN1(n6404), .IN2(n6403), .Q(n7332) );
  AND2X1 U350 ( .IN1(n6351), .IN2(n6350), .Q(n7331) );
  AND2X1 U346 ( .IN1(n6354), .IN2(n6353), .Q(n7330) );
  NBUFFX8 U12 ( .Z(n7479), .INP(n19025) );
  NOR2X2 U19984 ( .QN(P1_N5147), .IN1(n7052), .IN2(n7145) );
  NBUFFX4 U2042 ( .Z(n7116), .INP(P1_N5163) );
  NBUFFX4 U2039 ( .Z(n7113), .INP(P1_N5164) );
  NOR2X2 U19982 ( .QN(P2_N5069), .IN1(n7147), .IN2(n7265) );
  NBUFFX4 U2036 ( .Z(n7110), .INP(P1_N5165) );
  NBUFFX4 U2029 ( .Z(n7103), .INP(P1_N5167) );
  NBUFFX4 U2022 ( .Z(n7096), .INP(P1_N5169) );
  NBUFFX8 U2084 ( .Z(n7158), .INP(P2_N5078) );
  NBUFFX4 U2019 ( .Z(n7093), .INP(P1_N5170) );
  NBUFFX8 U2080 ( .Z(n7154), .INP(P2_N5079) );
  NBUFFX4 U1996 ( .Z(n7070), .INP(P1_N5158) );
  NBUFFX4 U2146 ( .Z(n7220), .INP(P2_N5081) );
  NBUFFX4 U1988 ( .Z(n7062), .INP(P1_N5160) );
  NBUFFX4 U1981 ( .Z(n7055), .INP(P1_N5162) );
  NBUFFX4 U2128 ( .Z(n7202), .INP(P2_N5086) );
  NBUFFX8 U2032 ( .Z(n7106), .INP(P1_N5166) );
  NBUFFX4 U2124 ( .Z(n7198), .INP(P2_N5087) );
  NBUFFX8 U2025 ( .Z(n7099), .INP(P1_N5168) );
  NBUFFX4 U1945 ( .Z(n7019), .INP(P1_N662) );
  NBUFFX4 U2099 ( .Z(n7173), .INP(P2_N5075) );
  NBUFFX4 U2048 ( .Z(n7122), .INP(P1_N5176) );
  NBUFFX4 U2050 ( .Z(n7124), .INP(P1_N5175) );
  NBUFFX8 U2067 ( .Z(n7141), .INP(P1_N5172) );
  NBUFFX4 U2153 ( .Z(n7227), .INP(P2_N5098) );
  NBUFFX4 U2157 ( .Z(n7231), .INP(P2_N5097) );
  INVX0 U1939 ( .ZN(n7013), .INP(n7012) );
  INVX0 U20011 ( .ZN(n2992), .INP(P2_N4178) );
  INVX0 U1736 ( .ZN(n6810), .INP(n6809) );
  INVX0 U19972 ( .ZN(n17734), .INP(P2_N5065) );
  INVX0 U20012 ( .ZN(n2657), .INP(P2_N4561) );
  INVX0 U16645 ( .ZN(n14521), .INP(P1_N5143) );
  NBUFFX4 U1705 ( .Z(n6779), .INP(P2_N291) );
  INVX0 U1708 ( .ZN(n6782), .INP(n6781) );
  NBUFFX4 U1739 ( .Z(n6813), .INP(n7485) );
  INVX0 U1768 ( .ZN(n6842), .INP(n6827) );
  NBUFFX4 U1833 ( .Z(n6907), .INP(n7483) );
  NBUFFX4 U1849 ( .Z(n6923), .INP(n7481) );
  INVX0 U1848 ( .ZN(n6922), .INP(n6921) );
  INVX0 U1800 ( .ZN(n6874), .INP(n7458) );
  INVX0 U1804 ( .ZN(n6878), .INP(P1_N291) );
  NBUFFX4 U1867 ( .Z(n6941), .INP(P2_N293) );
  NBUFFX4 U1895 ( .Z(n6969), .INP(P2_N294) );
  NAND2X1 U3056 ( .IN2(n6586), .IN1(n19025), .QN(P2_N5470) );
  INVX2 U2235 ( .INP(P2_N5485), .ZN(n7309) );
  NBUFFX2 U373 ( .Z(n6571), .INP(n7456) );
  NAND2X1 U8734 ( .IN2(n6332), .IN1(n6333), .QN(P1_N291) );
  NAND2X1 U1543 ( .IN2(P2_N584), .IN1(n1481), .QN(P2_N914) );
  NAND2X1 U1583 ( .IN2(P1_N584), .IN1(n1502), .QN(P1_N662) );
  INVX0 U364 ( .ZN(n6563), .INP(reset) );
  NBUFFX4 U377 ( .Z(n6575), .INP(n7455) );
  INVX0 U367 ( .ZN(n6566), .INP(reset) );
  NAND2X1 U8738 ( .IN2(n6334), .IN1(n6335), .QN(P1_N292) );
  NAND2X1 U8806 ( .IN2(n6384), .IN1(n6385), .QN(P2_N292) );
  NAND2X1 U8802 ( .IN2(n6382), .IN1(n6383), .QN(P2_N291) );
  INVX0 U362 ( .ZN(n6561), .INP(reset) );
  INVX0 U368 ( .ZN(n6567), .INP(reset) );
  INVX0 U1 ( .ZN(n6556), .INP(reset) );
  INVX0 U365 ( .ZN(n6564), .INP(reset) );
  INVX0 U8 ( .ZN(n6560), .INP(reset) );
  INVX0 U363 ( .ZN(n6562), .INP(reset) );
  INVX0 U5 ( .ZN(n6559), .INP(reset) );
  INVX0 U2 ( .ZN(n6557), .INP(reset) );
  INVX0 U366 ( .ZN(n6565), .INP(reset) );
  INVX0 U4 ( .ZN(n6558), .INP(reset) );
  INVX0 U2255 ( .ZN(n7329), .INP(n2178) );
  INVX0 U2238 ( .ZN(n7312), .INP(n4205) );
  INVX0 U2236 ( .ZN(n7310), .INP(n4208) );
  INVX1 U2229 ( .INP(P2_N5486), .ZN(n7303) );
  INVX1 U2225 ( .INP(P1_N5563), .ZN(n7299) );
  INVX1 U2221 ( .INP(P1_N5564), .ZN(n7295) );
  INVX1 U2217 ( .INP(P2_N5484), .ZN(n7291) );
  INVX1 U2213 ( .INP(P1_N5562), .ZN(n7287) );
  INVX1 U2205 ( .INP(P2_N5069), .ZN(n7279) );
  INVX0 U2201 ( .ZN(n7275), .INP(P2_N5015) );
  INVX0 U2200 ( .ZN(n7274), .INP(P1_N630) );
  INVX0 U2199 ( .ZN(n7273), .INP(P1_N5093) );
  INVX1 U2196 ( .INP(P2_N5476), .ZN(n7270) );
  INVX0 U2191 ( .ZN(n7265), .INP(P2_N497) );
  INVX0 U2190 ( .ZN(n7264), .INP(n7263) );
  INVX0 U2186 ( .ZN(n7260), .INP(n7259) );
  NBUFFX8 U2185 ( .Z(n7259), .INP(P2_N5091) );
  INVX0 U2179 ( .ZN(n7253), .INP(n7252) );
  NBUFFX8 U2178 ( .Z(n7252), .INP(P2_N5092) );
  INVX0 U2174 ( .ZN(n7248), .INP(n7247) );
  NBUFFX8 U2173 ( .Z(n7247), .INP(P2_N5093) );
  INVX0 U2169 ( .ZN(n7243), .INP(n7242) );
  NBUFFX8 U2168 ( .Z(n7242), .INP(P2_N5094) );
  INVX0 U2165 ( .ZN(n7239), .INP(n7238) );
  NBUFFX8 U2164 ( .Z(n7238), .INP(P2_N5095) );
  INVX0 U2160 ( .ZN(n7234), .INP(P2_N5096) );
  INVX0 U2155 ( .ZN(n7229), .INP(P2_N5097) );
  INVX0 U2150 ( .ZN(n7224), .INP(P2_N5098) );
  NBUFFX8 U2142 ( .Z(n7216), .INP(P2_N5082) );
  INVX0 U2140 ( .ZN(n7214), .INP(P2_N5082) );
  NBUFFX8 U2136 ( .Z(n7210), .INP(P2_N5083) );
  INVX0 U2121 ( .ZN(n7195), .INP(n7194) );
  NBUFFX8 U2120 ( .Z(n7194), .INP(P2_N5088) );
  INVX0 U2114 ( .ZN(n7188), .INP(n7187) );
  INVX0 U2108 ( .ZN(n7182), .INP(n7181) );
  NBUFFX8 U2107 ( .Z(n7181), .INP(P2_N5073) );
  INVX0 U2104 ( .ZN(n7178), .INP(n7177) );
  NBUFFX8 U2103 ( .Z(n7177), .INP(P2_N5074) );
  INVX0 U2100 ( .ZN(n7174), .INP(n7173) );
  INVX0 U2092 ( .ZN(n7166), .INP(n7165) );
  NBUFFX8 U2091 ( .Z(n7165), .INP(P2_N5076) );
  INVX0 U2090 ( .ZN(n7164), .INP(P2_N5077) );
  NBUFFX8 U2077 ( .Z(n7151), .INP(P2_N5080) );
  INVX0 U2073 ( .ZN(n7147), .INP(n2562) );
  INVX0 U2071 ( .ZN(n7145), .INP(P1_N497) );
  INVX0 U2070 ( .ZN(n7144), .INP(n7141) );
  NBUFFX8 U2064 ( .Z(n7138), .INP(P1_N5173) );
  INVX0 U2062 ( .ZN(n7136), .INP(n7138) );
  INVX0 U2056 ( .ZN(n7130), .INP(n7129) );
  NBUFFX8 U2055 ( .Z(n7129), .INP(P1_N5174) );
  INVX0 U2051 ( .ZN(n7125), .INP(n7124) );
  INVX0 U2045 ( .ZN(n7119), .INP(P1_N5176) );
  INVX0 U2016 ( .ZN(n7090), .INP(n7089) );
  NBUFFX8 U2015 ( .Z(n7089), .INP(P1_N5171) );
  INVX0 U2008 ( .ZN(n7082), .INP(n7081) );
  NBUFFX8 U2007 ( .Z(n7081), .INP(P1_N5154) );
  NBUFFX8 U2001 ( .Z(n7075), .INP(P1_N5156) );
  INVX0 U1999 ( .ZN(n7073), .INP(n7072) );
  NBUFFX8 U1998 ( .Z(n7072), .INP(P1_N5157) );
  INVX0 U1997 ( .ZN(n7071), .INP(n7070) );
  INVX0 U1993 ( .ZN(n7067), .INP(n7066) );
  INVX0 U1989 ( .ZN(n7063), .INP(n7062) );
  NBUFFX8 U1985 ( .Z(n7059), .INP(P1_N5161) );
  INVX0 U1982 ( .ZN(n7056), .INP(n7055) );
  INVX0 U1978 ( .ZN(n7052), .INP(n4469) );
  NBUFFX8 U1972 ( .Z(n7046), .INP(P1_N5151) );
  NBUFFX8 U1967 ( .Z(n7041), .INP(P1_N5152) );
  INVX0 U1963 ( .ZN(n7037), .INP(n7036) );
  NBUFFX8 U1962 ( .Z(n7036), .INP(P1_N5153) );
  INVX2 U1955 ( .INP(P1_N662), .ZN(n7029) );
  NBUFFX8 U1954 ( .Z(n7028), .INP(P1_N662) );
  INVX2 U1953 ( .INP(P1_N662), .ZN(n7027) );
  NBUFFX8 U1952 ( .Z(n7026), .INP(P1_N662) );
  NBUFFX8 U1950 ( .Z(n7024), .INP(P1_N662) );
  INVX1 U1949 ( .INP(n7022), .ZN(n7023) );
  NBUFFX8 U1948 ( .Z(n7022), .INP(P1_N662) );
  INVX2 U1947 ( .INP(P1_N662), .ZN(n7021) );
  NBUFFX8 U1942 ( .Z(n7016), .INP(n7462) );
  NBUFFX8 U1938 ( .Z(n7012), .INP(P2_N914) );
  INVX2 U1937 ( .INP(P2_N914), .ZN(n7011) );
  NBUFFX8 U1936 ( .Z(n7010), .INP(P2_N914) );
  NBUFFX8 U1935 ( .Z(n7009), .INP(P2_N914) );
  NBUFFX8 U1932 ( .Z(n7006), .INP(n7462) );
  INVX0 U1919 ( .ZN(n6993), .INP(n2693) );
  INVX1 U1918 ( .INP(n11309), .ZN(n6992) );
  INVX1 U1912 ( .INP(n14522), .ZN(n6986) );
  INVX2 U1908 ( .INP(n6981), .ZN(n6982) );
  NBUFFX8 U1907 ( .Z(n6981), .INP(P1_N294) );
  INVX1 U1902 ( .INP(n6975), .ZN(n6976) );
  INVX1 U1900 ( .INP(n6963), .ZN(n6974) );
  INVX1 U1896 ( .INP(n6969), .ZN(n6970) );
  NBUFFX8 U1889 ( .Z(n6963), .INP(P2_N294) );
  INVX1 U1888 ( .INP(n6961), .ZN(n6962) );
  NBUFFX8 U1887 ( .Z(n6961), .INP(P1_N293) );
  NBUFFX8 U1885 ( .Z(n6959), .INP(P1_N293) );
  INVX1 U1884 ( .INP(n6957), .ZN(n6958) );
  NBUFFX8 U1883 ( .Z(n6957), .INP(P1_N293) );
  INVX1 U1882 ( .INP(n6955), .ZN(n6956) );
  NBUFFX8 U1881 ( .Z(n6955), .INP(P1_N293) );
  INVX1 U1878 ( .INP(P1_N293), .ZN(n6952) );
  INVX0 U1874 ( .ZN(n6948), .INP(P2_N293) );
  INVX0 U1868 ( .ZN(n6942), .INP(n6941) );
  INVX0 U1854 ( .ZN(n6928), .INP(n2168) );
  INVX0 U1853 ( .ZN(n6927), .INP(n4171) );
  INVX0 U1852 ( .ZN(n6926), .INP(n6901) );
  NBUFFX8 U1847 ( .Z(n6921), .INP(n7481) );
  INVX1 U1846 ( .INP(n6919), .ZN(n6920) );
  NBUFFX8 U1845 ( .Z(n6919), .INP(P1_N292) );
  INVX0 U1832 ( .ZN(n6906), .INP(n7481) );
  INVX1 U1830 ( .INP(n7483), .ZN(n6904) );
  NBUFFX8 U1827 ( .Z(n6901), .INP(P1_N292) );
  INVX0 U1820 ( .ZN(n6894), .INP(n6893) );
  INVX0 U1818 ( .ZN(n6892), .INP(n6891) );
  INVX1 U1816 ( .INP(P1_N292), .ZN(n6890) );
  INVX1 U1814 ( .INP(n6887), .ZN(n6888) );
  NBUFFX8 U1813 ( .Z(n6887), .INP(n7483) );
  INVX1 U1812 ( .INP(n7481), .ZN(n6886) );
  INVX1 U1810 ( .INP(n6883), .ZN(n6884) );
  INVX1 U1808 ( .INP(n6881), .ZN(n6882) );
  NBUFFX8 U1807 ( .Z(n6881), .INP(n7481) );
  INVX1 U1798 ( .INP(n6871), .ZN(n6872) );
  NBUFFX8 U1797 ( .Z(n6871), .INP(n7458) );
  NBUFFX8 U1793 ( .Z(n6867), .INP(P1_N291) );
  INVX1 U1792 ( .INP(n6865), .ZN(n6866) );
  NBUFFX16 U1791 ( .Z(n6865), .INP(n7458) );
  INVX1 U1790 ( .INP(n6867), .ZN(n6864) );
  INVX2 U1788 ( .INP(n6861), .ZN(n6862) );
  NBUFFX8 U1787 ( .Z(n6861), .INP(P1_N291) );
  NBUFFX8 U1783 ( .Z(n6857), .INP(P1_N291) );
  INVX1 U1782 ( .INP(n6855), .ZN(n6856) );
  INVX1 U1778 ( .INP(n6851), .ZN(n6852) );
  INVX0 U1762 ( .ZN(n6836), .INP(n6835) );
  INVX1 U1758 ( .INP(n6831), .ZN(n6832) );
  NBUFFX8 U1757 ( .Z(n6831), .INP(n7484) );
  INVX0 U1756 ( .ZN(n6830), .INP(n6829) );
  INVX1 U1754 ( .INP(n6827), .ZN(n6828) );
  NBUFFX8 U1753 ( .Z(n6827), .INP(n7485) );
  NBUFFX8 U1751 ( .Z(n6825), .INP(n7486) );
  NBUFFX8 U1749 ( .Z(n6823), .INP(P2_N292) );
  INVX1 U1748 ( .INP(n7486), .ZN(n6822) );
  INVX1 U1746 ( .INP(n6819), .ZN(n6820) );
  INVX1 U1744 ( .INP(n6823), .ZN(n6818) );
  INVX1 U1742 ( .INP(n6815), .ZN(n6816) );
  INVX1 U1738 ( .INP(n7486), .ZN(n6812) );
  NBUFFX8 U1733 ( .Z(n6807), .INP(n7484) );
  INVX1 U1730 ( .INP(n6803), .ZN(n6804) );
  NBUFFX8 U1729 ( .Z(n6803), .INP(P2_N291) );
  INVX0 U1720 ( .ZN(n6794), .INP(n6793) );
  NBUFFX8 U1719 ( .Z(n6793), .INP(n7488) );
  INVX0 U1718 ( .ZN(n6792), .INP(n6787) );
  INVX1 U1716 ( .INP(n6789), .ZN(n6790) );
  NBUFFX8 U1715 ( .Z(n6789), .INP(n7487) );
  INVX1 U1712 ( .INP(n6775), .ZN(n6786) );
  INVX1 U1710 ( .INP(n6793), .ZN(n6784) );
  INVX1 U1706 ( .INP(n6779), .ZN(n6780) );
  INVX1 U1702 ( .INP(n6775), .ZN(n6776) );
  NBUFFX8 U1701 ( .Z(n6775), .INP(n7487) );
  INVX0 U1700 ( .ZN(n6774), .INP(P2_N345) );
  INVX0 U1699 ( .ZN(n6773), .INP(P1_N345) );
  INVX0 U1698 ( .ZN(n6772), .INP(P2_N346) );
  INVX0 U1697 ( .ZN(n6771), .INP(P2_N344) );
  INVX0 U1696 ( .ZN(n6770), .INP(P1_N346) );
  INVX0 U1695 ( .ZN(n6769), .INP(P2_N349) );
  INVX0 U1694 ( .ZN(n6768), .INP(P2_N347) );
  INVX0 U1693 ( .ZN(n6767), .INP(P1_N349) );
  INVX0 U1692 ( .ZN(n6766), .INP(P1_N347) );
  INVX0 U1691 ( .ZN(n6765), .INP(P2_N350) );
  INVX0 U1690 ( .ZN(n6764), .INP(P2_N348) );
  INVX0 U1689 ( .ZN(n6763), .INP(P1_N350) );
  INVX0 U1688 ( .ZN(n6762), .INP(P1_N348) );
  INVX0 U1687 ( .ZN(n6761), .INP(P2_N351) );
  INVX0 U1686 ( .ZN(n6760), .INP(P2_N353) );
  INVX0 U1685 ( .ZN(n6759), .INP(P1_N353) );
  INVX0 U1684 ( .ZN(n6758), .INP(P1_N351) );
  INVX0 U1683 ( .ZN(n6757), .INP(P2_N354) );
  INVX0 U1682 ( .ZN(n6756), .INP(P2_N352) );
  INVX0 U1681 ( .ZN(n6755), .INP(P1_N354) );
  INVX0 U1680 ( .ZN(n6754), .INP(P1_N352) );
  INVX0 U1679 ( .ZN(n6753), .INP(P2_N357) );
  INVX0 U1678 ( .ZN(n6752), .INP(P2_N355) );
  INVX0 U1677 ( .ZN(n6751), .INP(P1_N357) );
  INVX0 U1676 ( .ZN(n6750), .INP(P1_N355) );
  INVX0 U1675 ( .ZN(n6749), .INP(P2_N358) );
  INVX0 U1674 ( .ZN(n6748), .INP(P2_N356) );
  INVX0 U1673 ( .ZN(n6747), .INP(P1_N358) );
  INVX0 U1672 ( .ZN(n6746), .INP(P1_N356) );
  INVX0 U1671 ( .ZN(n6745), .INP(P2_N359) );
  INVX0 U1670 ( .ZN(n6744), .INP(P1_N359) );
  INVX0 U1669 ( .ZN(n6743), .INP(P2_N360) );
  INVX0 U1668 ( .ZN(n6742), .INP(P1_N360) );
  NBUFFX8 U1662 ( .Z(n6736), .INP(N5) );
  INVX0 U1661 ( .ZN(n6735), .INP(P2_N361) );
  INVX0 U1660 ( .ZN(n6734), .INP(P1_N361) );
  INVX0 U1659 ( .ZN(n6733), .INP(P2_N362) );
  INVX0 U1658 ( .ZN(n6732), .INP(P1_N362) );
  INVX0 U1657 ( .ZN(n6731), .INP(P2_N363) );
  INVX0 U1656 ( .ZN(n6730), .INP(P1_N363) );
  INVX0 U1651 ( .ZN(n6725), .INP(P1_N5548) );
  INVX0 U1647 ( .ZN(n6721), .INP(n18995) );
  INVX0 U1646 ( .ZN(n6720), .INP(n18997) );
  INVX0 U1645 ( .ZN(n6719), .INP(n19001) );
  INVX0 U1640 ( .ZN(n6714), .INP(n6713) );
  INVX0 U1628 ( .ZN(n6702), .INP(n6687) );
  INVX0 U1626 ( .ZN(n6700), .INP(n6699) );
  INVX0 U1624 ( .ZN(n6698), .INP(n7479) );
  INVX0 U1622 ( .ZN(n6696), .INP(n6687) );
  NBUFFX8 U1613 ( .Z(n6687), .INP(n19025) );
  INVX0 U1612 ( .ZN(n6686), .INP(n6685) );
  INVX0 U1610 ( .ZN(n6684), .INP(n18813) );
  INVX0 U1606 ( .ZN(n6680), .INP(n18907) );
  INVX0 U1605 ( .ZN(n6679), .INP(n18909) );
  INVX0 U1604 ( .ZN(n6678), .INP(n18911) );
  INVX0 U1603 ( .ZN(n6677), .INP(n18913) );
  INVX0 U1602 ( .ZN(n6676), .INP(n18915) );
  INVX0 U1601 ( .ZN(n6675), .INP(n18917) );
  INVX0 U1600 ( .ZN(n6674), .INP(n18919) );
  INVX0 U1599 ( .ZN(n6673), .INP(n18921) );
  INVX0 U1598 ( .ZN(n6672), .INP(n18923) );
  INVX0 U1597 ( .ZN(n6671), .INP(n18925) );
  INVX0 U1596 ( .ZN(n6670), .INP(n18927) );
  INVX0 U1595 ( .ZN(n6669), .INP(n18929) );
  INVX0 U1594 ( .ZN(n6668), .INP(n18931) );
  INVX0 U1593 ( .ZN(n6667), .INP(n18933) );
  INVX0 U1592 ( .ZN(n6666), .INP(n18935) );
  INVX0 U1591 ( .ZN(n6665), .INP(n18937) );
  INVX0 U1590 ( .ZN(n6664), .INP(n18939) );
  INVX0 U1589 ( .ZN(n6663), .INP(n18963) );
  INVX0 U1588 ( .ZN(n6662), .INP(n18965) );
  INVX0 U1587 ( .ZN(n6661), .INP(n18967) );
  INVX0 U1586 ( .ZN(n6660), .INP(n18969) );
  INVX0 U1585 ( .ZN(n6659), .INP(n18971) );
  INVX0 U1580 ( .ZN(n6658), .INP(n18973) );
  INVX0 U1512 ( .ZN(n6657), .INP(n18975) );
  INVX0 U1425 ( .ZN(n6656), .INP(n18977) );
  INVX0 U1334 ( .ZN(n6655), .INP(n18979) );
  INVX0 U1243 ( .ZN(n6654), .INP(n18981) );
  INVX0 U1145 ( .ZN(n6653), .INP(n18983) );
  INVX0 U1081 ( .ZN(n6652), .INP(n18985) );
  INVX0 U973 ( .ZN(n6651), .INP(n18987) );
  INVX0 U877 ( .ZN(n6650), .INP(n18989) );
  INVX0 U786 ( .ZN(n6649), .INP(n18991) );
  INVX0 U695 ( .ZN(n6648), .INP(n18993) );
  INVX0 U603 ( .ZN(n6647), .INP(n18643) );
  INVX0 U542 ( .ZN(n6646), .INP(n18645) );
  INVX0 U470 ( .ZN(n6645), .INP(n18647) );
  INVX0 U469 ( .ZN(n6644), .INP(n18649) );
  INVX0 U468 ( .ZN(n6643), .INP(n18651) );
  INVX0 U463 ( .ZN(n6642), .INP(n18653) );
  INVX0 U462 ( .ZN(n6641), .INP(n18655) );
  INVX0 U455 ( .ZN(n6640), .INP(n18657) );
  INVX0 U454 ( .ZN(n6639), .INP(n18659) );
  INVX0 U453 ( .ZN(n6638), .INP(n18661) );
  INVX0 U452 ( .ZN(n6637), .INP(n18663) );
  INVX0 U451 ( .ZN(n6636), .INP(n18671) );
  INVX0 U450 ( .ZN(n6635), .INP(n18673) );
  INVX0 U449 ( .ZN(n6634), .INP(n18675) );
  INVX0 U447 ( .ZN(n6633), .INP(n18677) );
  INVX0 U446 ( .ZN(n6632), .INP(n18679) );
  INVX0 U445 ( .ZN(n6631), .INP(n18681) );
  INVX0 U444 ( .ZN(n6630), .INP(n18683) );
  INVX0 U443 ( .ZN(n6629), .INP(n18685) );
  INVX0 U442 ( .ZN(n6628), .INP(n18687) );
  INVX0 U441 ( .ZN(n6627), .INP(n18689) );
  INVX0 U440 ( .ZN(n6626), .INP(n18691) );
  INVX0 U439 ( .ZN(n6625), .INP(n18693) );
  INVX0 U427 ( .ZN(n6617), .INP(n18297) );
  INVX0 U426 ( .ZN(n6616), .INP(n18299) );
  INVX0 U419 ( .ZN(n6615), .INP(n18301) );
  INVX0 U417 ( .ZN(n6614), .INP(n18303) );
  INVX0 U416 ( .ZN(n6613), .INP(n18305) );
  INVX0 U415 ( .ZN(n6612), .INP(n18307) );
  INVX0 U414 ( .ZN(n6611), .INP(n18309) );
  INVX0 U413 ( .ZN(n6610), .INP(n18311) );
  INVX0 U412 ( .ZN(n6609), .INP(n18313) );
  INVX0 U411 ( .ZN(n6608), .INP(n18315) );
  INVX0 U410 ( .ZN(n6607), .INP(n18323) );
  INVX0 U409 ( .ZN(n6606), .INP(n18325) );
  INVX0 U408 ( .ZN(n6605), .INP(n18327) );
  INVX0 U407 ( .ZN(n6604), .INP(n18329) );
  INVX0 U406 ( .ZN(n6603), .INP(n18331) );
  INVX0 U405 ( .ZN(n6602), .INP(n18333) );
  INVX0 U404 ( .ZN(n6601), .INP(n18335) );
  INVX0 U403 ( .ZN(n6600), .INP(n18337) );
  INVX0 U402 ( .ZN(n6599), .INP(n18339) );
  INVX0 U397 ( .ZN(n6594), .INP(n18451) );
  INVX0 U393 ( .ZN(n6590), .INP(n6589) );
  NBUFFX8 U392 ( .Z(n6589), .INP(n2166) );
  INVX0 U390 ( .ZN(n6588), .INP(n2166) );
  NBUFFX8 U385 ( .Z(n6583), .INP(n4169) );
  NBUFFX8 U382 ( .Z(n6580), .INP(n4169) );
  NAND2X1 U8693 ( .IN2(n5946), .IN1(n5945), .QN(n4150) );
  NAND2X1 U8699 ( .IN2(n5949), .IN1(n5948), .QN(n4153) );
  NAND2X1 U8705 ( .IN2(n5952), .IN1(n5951), .QN(n4156) );
  NAND2X1 U8687 ( .IN2(n5943), .IN1(n5942), .QN(n4147) );
  NAND2X1 U8681 ( .IN2(n5940), .IN1(n5939), .QN(n4144) );
  NAND2X1 U8675 ( .IN2(n5937), .IN1(n5936), .QN(n4141) );
  NAND2X1 U8669 ( .IN2(n5934), .IN1(n5933), .QN(n4138) );
  NAND2X1 U5553 ( .IN2(n3887), .IN1(n3886), .QN(n2044) );
  NAND2X1 U8750 ( .IN2(n6347), .IN1(n6348), .QN(P1_N294) );
  NAND2X1 U5544 ( .IN2(n3882), .IN1(n3881), .QN(n2041) );
  NAND2X1 U5680 ( .IN2(n3964), .IN1(n3963), .QN(P2_N925) );
  NAND2X1 U5508 ( .IN2(n3862), .IN1(n3861), .QN(n2029) );
  NAND2X1 U5499 ( .IN2(n3857), .IN1(n3856), .QN(n2026) );
  NAND2X1 U5665 ( .IN2(n3952), .IN1(n3951), .QN(P2_N928) );
  NAND2X1 U5490 ( .IN2(n3852), .IN1(n3851), .QN(n2023) );
  NAND2X1 U5660 ( .IN2(n3948), .IN1(n3947), .QN(P2_N929) );
  NAND2X1 U5481 ( .IN2(n3847), .IN1(n3846), .QN(n2020) );
  NAND2X1 U5472 ( .IN2(n3842), .IN1(n3841), .QN(n2017) );
  NAND2X1 U5463 ( .IN2(n3837), .IN1(n3836), .QN(n2014) );
  NAND2X1 U8591 ( .IN2(n5895), .IN1(n5894), .QN(n4099) );
  NAND2X1 U5445 ( .IN2(n3827), .IN1(n3826), .QN(n2008) );
  NAND2X1 U8812 ( .IN2(n6388), .IN1(n6389), .QN(P2_N293) );
  NAND2X1 U8744 ( .IN2(n6338), .IN1(n6339), .QN(P1_N293) );
  NAND2X1 U8818 ( .IN2(n6397), .IN1(n6398), .QN(P2_N294) );
  NAND2X1 U8651 ( .IN2(n5925), .IN1(n5924), .QN(n4129) );
  NAND2X1 U8624 ( .IN2(P1_N349), .IN1(P1_N583), .QN(n4112) );
  NAND2X1 U8630 ( .IN2(P1_N350), .IN1(P1_N583), .QN(n4115) );
  NAND2X1 U8636 ( .IN2(P1_N351), .IN1(P1_N583), .QN(n4118) );
  NAND2X1 U8642 ( .IN2(P1_N352), .IN1(P1_N583), .QN(n4121) );
  NAND2X1 U8648 ( .IN2(P1_N353), .IN1(P1_N583), .QN(n4124) );
  NAND2X1 U8654 ( .IN2(P1_N354), .IN1(P1_N583), .QN(n4127) );
  NAND2X1 U8672 ( .IN2(P1_N357), .IN1(P1_N583), .QN(n4136) );
  NAND2X1 U5502 ( .IN2(n2693), .IN1(P2_N350), .QN(n2024) );
  NAND2X1 U5511 ( .IN2(n2693), .IN1(P2_N351), .QN(n2027) );
  NAND2X1 U5520 ( .IN2(n2693), .IN1(P2_N352), .QN(n2030) );
  NAND2X1 U8645 ( .IN2(n5922), .IN1(n5921), .QN(n4126) );
  NAND2X1 U8639 ( .IN2(n5919), .IN1(n5918), .QN(n4123) );
  NAND2X1 U6188 ( .IN2(n4376), .IN1(n4375), .QN(P1_N536) );
  NAND2X1 U3302 ( .IN2(n2469), .IN1(n2468), .QN(P2_N536) );
  NAND2X1 U8633 ( .IN2(n5916), .IN1(n5915), .QN(n4120) );
  NAND2X1 U8627 ( .IN2(n5913), .IN1(n5912), .QN(n4117) );
  NOR2X2 U8226 ( .QN(n5623), .IN1(n7358), .IN2(n7357) );
  NOR2X2 U8048 ( .QN(n5511), .IN1(n7360), .IN2(n7359) );
  NOR2X2 U7897 ( .QN(n5425), .IN1(n7362), .IN2(n7361) );
  NOR2X2 U7722 ( .QN(n5316), .IN1(n7364), .IN2(n7363) );
  NOR2X2 U7552 ( .QN(n5212), .IN1(n7366), .IN2(n7365) );
  NOR2X2 U7401 ( .QN(n5104), .IN1(n7368), .IN2(n7367) );
  NOR2X2 U7227 ( .QN(n5018), .IN1(n7370), .IN2(n7369) );
  NOR2X2 U7076 ( .QN(n4932), .IN1(n7372), .IN2(n7371) );
  NOR2X2 U6925 ( .QN(n4818), .IN1(n7374), .IN2(n7373) );
  NAND2X1 U8621 ( .IN2(n5910), .IN1(n5909), .QN(n4114) );
  NAND2X1 U1530 ( .IN2(P2_N4626), .IN1(n1474), .QN(P2_N5497) );
  NAND2X1 U8615 ( .IN2(n5907), .IN1(n5906), .QN(n4111) );
  NAND2X1 U8609 ( .IN2(n5904), .IN1(n5903), .QN(n4108) );
  NAND2X1 U5454 ( .IN2(n3832), .IN1(n3831), .QN(n2011) );
  INVX0 U12460 ( .ZN(n18952), .INP(n18953) );
  INVX0 U12463 ( .ZN(n18954), .INP(n18955) );
  INVX0 U12466 ( .ZN(n18956), .INP(n18957) );
  INVX0 U12469 ( .ZN(n18958), .INP(n18959) );
  INVX0 U12472 ( .ZN(n18960), .INP(n18961) );
  INVX0 U12529 ( .ZN(n18998), .INP(n18999) );
  INVX0 U12535 ( .ZN(n19002), .INP(n19003) );
  INVX0 U12538 ( .ZN(n19004), .INP(n19005) );
  INVX0 U12541 ( .ZN(n19006), .INP(n19007) );
  INVX0 U12547 ( .ZN(n19010), .INP(n19011) );
  INVX0 U12550 ( .ZN(n19012), .INP(n19013) );
  INVX0 U12553 ( .ZN(n19014), .INP(n19015) );
  INVX0 U12556 ( .ZN(n19016), .INP(n19017) );
  INVX0 U12559 ( .ZN(n19018), .INP(n19019) );
  INVX0 U12562 ( .ZN(n19020), .INP(n19021) );
  INVX0 U12565 ( .ZN(n19022), .INP(n19023) );
  INVX0 U12155 ( .ZN(n18766), .INP(n18767) );
  INVX0 U12158 ( .ZN(n18768), .INP(n18769) );
  INVX0 U12161 ( .ZN(n18770), .INP(n18771) );
  INVX0 U12164 ( .ZN(n18772), .INP(n18773) );
  INVX0 U12167 ( .ZN(n18774), .INP(n18775) );
  INVX0 U12170 ( .ZN(n18776), .INP(n18777) );
  INVX0 U12173 ( .ZN(n18778), .INP(n18779) );
  INVX0 U12176 ( .ZN(n18780), .INP(n18781) );
  INVX0 U12179 ( .ZN(n18782), .INP(n18783) );
  INVX0 U12182 ( .ZN(n18784), .INP(n18785) );
  INVX0 U12185 ( .ZN(n18786), .INP(n18787) );
  INVX0 U12188 ( .ZN(n18788), .INP(n18789) );
  INVX0 U12191 ( .ZN(n18790), .INP(n18791) );
  INVX0 U12194 ( .ZN(n18792), .INP(n18793) );
  INVX0 U12197 ( .ZN(n18794), .INP(n18795) );
  INVX0 U12200 ( .ZN(n18796), .INP(n18797) );
  INVX0 U12203 ( .ZN(n18798), .INP(n18799) );
  INVX0 U12206 ( .ZN(n18800), .INP(n18801) );
  INVX0 U12209 ( .ZN(n18802), .INP(n18803) );
  INVX0 U12212 ( .ZN(n18804), .INP(n18805) );
  INVX0 U12215 ( .ZN(n18806), .INP(n18807) );
  INVX0 U12218 ( .ZN(n18808), .INP(n18809) );
  INVX0 U12221 ( .ZN(n18810), .INP(n18811) );
  INVX0 U12230 ( .ZN(n18820), .INP(n18821) );
  INVX0 U12234 ( .ZN(n18822), .INP(n18823) );
  INVX0 U12235 ( .ZN(n18824), .INP(n18825) );
  INVX0 U12238 ( .ZN(n18826), .INP(n18827) );
  INVX0 U12241 ( .ZN(n18828), .INP(n18829) );
  INVX0 U12244 ( .ZN(n18830), .INP(n18831) );
  INVX0 U12247 ( .ZN(n18832), .INP(n18833) );
  INVX0 U12250 ( .ZN(n18834), .INP(n18835) );
  INVX0 U12253 ( .ZN(n18836), .INP(n18837) );
  INVX0 U12256 ( .ZN(n18838), .INP(n18839) );
  INVX0 U12259 ( .ZN(n18840), .INP(n18841) );
  INVX0 U12262 ( .ZN(n18842), .INP(n18843) );
  INVX0 U12265 ( .ZN(n18844), .INP(n18845) );
  INVX0 U12268 ( .ZN(n18846), .INP(n18847) );
  INVX0 U12271 ( .ZN(n18848), .INP(n18849) );
  INVX0 U12274 ( .ZN(n18850), .INP(n18851) );
  INVX0 U12277 ( .ZN(n18852), .INP(n18853) );
  INVX0 U12281 ( .ZN(n18854), .INP(n18855) );
  INVX0 U12285 ( .ZN(n18856), .INP(n18857) );
  INVX0 U12288 ( .ZN(n18858), .INP(n18859) );
  INVX0 U12291 ( .ZN(n18860), .INP(n18861) );
  INVX0 U12294 ( .ZN(n18862), .INP(n18863) );
  INVX0 U12297 ( .ZN(n18864), .INP(n18865) );
  INVX0 U12301 ( .ZN(n18866), .INP(n18867) );
  INVX0 U12305 ( .ZN(n18868), .INP(n18869) );
  INVX0 U12309 ( .ZN(n18870), .INP(n18871) );
  INVX0 U12313 ( .ZN(n18872), .INP(n18873) );
  INVX0 U12317 ( .ZN(n18874), .INP(n18875) );
  INVX0 U12321 ( .ZN(n18876), .INP(n18877) );
  INVX0 U12325 ( .ZN(n18878), .INP(n18879) );
  INVX0 U12329 ( .ZN(n18880), .INP(n18881) );
  INVX0 U12333 ( .ZN(n18882), .INP(n18883) );
  INVX0 U12337 ( .ZN(n18884), .INP(n18885) );
  INVX0 U12338 ( .ZN(n18886), .INP(n18887) );
  INVX0 U12341 ( .ZN(n18888), .INP(n18889) );
  INVX0 U12345 ( .ZN(n18890), .INP(n18891) );
  INVX0 U12349 ( .ZN(n18892), .INP(n18893) );
  INVX0 U12353 ( .ZN(n18894), .INP(n18895) );
  INVX0 U12357 ( .ZN(n18896), .INP(n18897) );
  INVX0 U12361 ( .ZN(n18898), .INP(n18899) );
  INVX0 U12365 ( .ZN(n18900), .INP(n18901) );
  INVX0 U12369 ( .ZN(n18902), .INP(n18903) );
  INVX0 U12373 ( .ZN(n18904), .INP(n18905) );
  INVX0 U12442 ( .ZN(n18940), .INP(n18941) );
  INVX0 U12445 ( .ZN(n18942), .INP(n18943) );
  INVX0 U12448 ( .ZN(n18944), .INP(n18945) );
  INVX0 U12451 ( .ZN(n18946), .INP(n18947) );
  INVX0 U12454 ( .ZN(n18948), .INP(n18949) );
  INVX0 U12457 ( .ZN(n18950), .INP(n18951) );
  INVX0 U11877 ( .ZN(n18580), .INP(n18581) );
  INVX0 U11880 ( .ZN(n18582), .INP(n18583) );
  INVX0 U11883 ( .ZN(n18584), .INP(n18585) );
  INVX0 U11886 ( .ZN(n18586), .INP(n18587) );
  INVX0 U11889 ( .ZN(n18588), .INP(n18589) );
  INVX0 U11892 ( .ZN(n18590), .INP(n18591) );
  INVX0 U11895 ( .ZN(n18592), .INP(n18593) );
  INVX0 U11898 ( .ZN(n18594), .INP(n18595) );
  INVX0 U11901 ( .ZN(n18596), .INP(n18597) );
  INVX0 U11904 ( .ZN(n18598), .INP(n18599) );
  INVX0 U11907 ( .ZN(n18600), .INP(n18601) );
  INVX0 U11910 ( .ZN(n18602), .INP(n18603) );
  INVX0 U11913 ( .ZN(n18604), .INP(n18605) );
  INVX0 U11916 ( .ZN(n18606), .INP(n18607) );
  INVX0 U11919 ( .ZN(n18608), .INP(n18609) );
  INVX0 U11922 ( .ZN(n18610), .INP(n18611) );
  INVX0 U11925 ( .ZN(n18612), .INP(n18613) );
  INVX0 U11928 ( .ZN(n18614), .INP(n18615) );
  INVX0 U11931 ( .ZN(n18616), .INP(n18617) );
  INVX0 U11934 ( .ZN(n18618), .INP(n18619) );
  INVX0 U11937 ( .ZN(n18620), .INP(n18621) );
  INVX0 U11940 ( .ZN(n18622), .INP(n18623) );
  INVX0 U11943 ( .ZN(n18624), .INP(n18625) );
  INVX0 U11946 ( .ZN(n18626), .INP(n18627) );
  INVX0 U11947 ( .ZN(n18628), .INP(n18629) );
  INVX0 U11949 ( .ZN(n18630), .INP(n18631) );
  INVX0 U11952 ( .ZN(n18632), .INP(n18633) );
  INVX0 U11955 ( .ZN(n18634), .INP(n18635) );
  INVX0 U11958 ( .ZN(n18636), .INP(n18637) );
  INVX0 U11961 ( .ZN(n18638), .INP(n18639) );
  INVX0 U11964 ( .ZN(n18640), .INP(n18641) );
  INVX0 U12000 ( .ZN(n18664), .INP(n18665) );
  INVX0 U12003 ( .ZN(n18666), .INP(n18667) );
  INVX0 U12006 ( .ZN(n18668), .INP(n18669) );
  INVX0 U12050 ( .ZN(n18696), .INP(n18697) );
  INVX0 U12053 ( .ZN(n18698), .INP(n18699) );
  INVX0 U12056 ( .ZN(n18700), .INP(n18701) );
  INVX0 U12059 ( .ZN(n18702), .INP(n18703) );
  INVX0 U12062 ( .ZN(n18704), .INP(n18705) );
  INVX0 U12065 ( .ZN(n18706), .INP(n18707) );
  INVX0 U12068 ( .ZN(n18708), .INP(n18709) );
  INVX0 U12071 ( .ZN(n18710), .INP(n18711) );
  INVX0 U12074 ( .ZN(n18712), .INP(n18713) );
  INVX0 U12077 ( .ZN(n18714), .INP(n18715) );
  INVX0 U12080 ( .ZN(n18716), .INP(n18717) );
  INVX0 U12083 ( .ZN(n18718), .INP(n18719) );
  INVX0 U12086 ( .ZN(n18720), .INP(n18721) );
  INVX0 U12089 ( .ZN(n18722), .INP(n18723) );
  INVX0 U12092 ( .ZN(n18724), .INP(n18725) );
  INVX0 U12095 ( .ZN(n18726), .INP(n18727) );
  INVX0 U12098 ( .ZN(n18728), .INP(n18729) );
  INVX0 U12101 ( .ZN(n18730), .INP(n18731) );
  INVX0 U12104 ( .ZN(n18732), .INP(n18733) );
  INVX0 U12107 ( .ZN(n18734), .INP(n18735) );
  INVX0 U12110 ( .ZN(n18736), .INP(n18737) );
  INVX0 U12113 ( .ZN(n18738), .INP(n18739) );
  INVX0 U12116 ( .ZN(n18740), .INP(n18741) );
  INVX0 U12119 ( .ZN(n18742), .INP(n18743) );
  INVX0 U12122 ( .ZN(n18744), .INP(n18745) );
  INVX0 U12125 ( .ZN(n18746), .INP(n18747) );
  INVX0 U12128 ( .ZN(n18748), .INP(n18749) );
  INVX0 U12131 ( .ZN(n18750), .INP(n18751) );
  INVX0 U12134 ( .ZN(n18752), .INP(n18753) );
  INVX0 U12137 ( .ZN(n18754), .INP(n18755) );
  INVX0 U12140 ( .ZN(n18756), .INP(n18757) );
  INVX0 U12143 ( .ZN(n18758), .INP(n18759) );
  INVX0 U12146 ( .ZN(n18760), .INP(n18761) );
  INVX0 U12149 ( .ZN(n18762), .INP(n18763) );
  INVX0 U12152 ( .ZN(n18764), .INP(n18765) );
  INVX0 U11603 ( .ZN(n18394), .INP(n18395) );
  INVX0 U11606 ( .ZN(n18396), .INP(n18397) );
  INVX0 U11609 ( .ZN(n18398), .INP(n18399) );
  INVX0 U11612 ( .ZN(n18400), .INP(n18401) );
  INVX0 U11615 ( .ZN(n18402), .INP(n18403) );
  INVX0 U11618 ( .ZN(n18404), .INP(n18405) );
  INVX0 U11621 ( .ZN(n18406), .INP(n18407) );
  INVX0 U11624 ( .ZN(n18408), .INP(n18409) );
  INVX0 U11627 ( .ZN(n18410), .INP(n18411) );
  INVX0 U11630 ( .ZN(n18412), .INP(n18413) );
  INVX0 U11633 ( .ZN(n18414), .INP(n18415) );
  INVX0 U11636 ( .ZN(n18416), .INP(n18417) );
  INVX0 U11639 ( .ZN(n18418), .INP(n18419) );
  INVX0 U11642 ( .ZN(n18420), .INP(n18421) );
  INVX0 U11645 ( .ZN(n18422), .INP(n18423) );
  INVX0 U11648 ( .ZN(n18424), .INP(n18425) );
  INVX0 U11651 ( .ZN(n18426), .INP(n18427) );
  INVX0 U11654 ( .ZN(n18428), .INP(n18429) );
  INVX0 U11657 ( .ZN(n18430), .INP(n18431) );
  INVX0 U11660 ( .ZN(n18432), .INP(n18433) );
  INVX0 U11663 ( .ZN(n18434), .INP(n18435) );
  INVX0 U11666 ( .ZN(n18436), .INP(n18437) );
  INVX0 U11669 ( .ZN(n18438), .INP(n18439) );
  INVX0 U11672 ( .ZN(n18440), .INP(n18441) );
  INVX0 U11675 ( .ZN(n18442), .INP(n18443) );
  INVX0 U11678 ( .ZN(n18444), .INP(n18445) );
  INVX0 U11681 ( .ZN(n18446), .INP(n18447) );
  INVX0 U11684 ( .ZN(n18448), .INP(n18449) );
  INVX0 U11690 ( .ZN(n18452), .INP(n18453) );
  INVX0 U11696 ( .ZN(n18456), .INP(n18457) );
  INVX0 U11702 ( .ZN(n18460), .INP(n18461) );
  INVX0 U11705 ( .ZN(n18462), .INP(n18463) );
  INVX0 U11711 ( .ZN(n18466), .INP(n18467) );
  INVX0 U11714 ( .ZN(n18468), .INP(n18469) );
  INVX0 U11717 ( .ZN(n18470), .INP(n18471) );
  INVX0 U11720 ( .ZN(n18472), .INP(n18473) );
  INVX0 U11723 ( .ZN(n18474), .INP(n18475) );
  INVX0 U11726 ( .ZN(n18476), .INP(n18477) );
  INVX0 U11729 ( .ZN(n18478), .INP(n18479) );
  INVX0 U11732 ( .ZN(n18480), .INP(n18481) );
  INVX0 U11735 ( .ZN(n18482), .INP(n18483) );
  INVX0 U11736 ( .ZN(n18484), .INP(n18485) );
  INVX0 U11738 ( .ZN(n18486), .INP(n18487) );
  INVX0 U11741 ( .ZN(n18488), .INP(n18489) );
  INVX0 U11744 ( .ZN(n18490), .INP(n18491) );
  INVX0 U11747 ( .ZN(n18492), .INP(n18493) );
  INVX0 U11750 ( .ZN(n18494), .INP(n18495) );
  INVX0 U11753 ( .ZN(n18496), .INP(n18497) );
  INVX0 U11756 ( .ZN(n18498), .INP(n18499) );
  INVX0 U11759 ( .ZN(n18500), .INP(n18501) );
  INVX0 U11762 ( .ZN(n18502), .INP(n18503) );
  INVX0 U11765 ( .ZN(n18504), .INP(n18505) );
  INVX0 U11768 ( .ZN(n18506), .INP(n18507) );
  INVX0 U11769 ( .ZN(n18508), .INP(n18509) );
  INVX0 U11771 ( .ZN(n18510), .INP(n18511) );
  INVX0 U11774 ( .ZN(n18512), .INP(n18513) );
  INVX0 U11777 ( .ZN(n18514), .INP(n18515) );
  INVX0 U11780 ( .ZN(n18516), .INP(n18517) );
  INVX0 U11783 ( .ZN(n18518), .INP(n18519) );
  INVX0 U11786 ( .ZN(n18520), .INP(n18521) );
  INVX0 U11789 ( .ZN(n18522), .INP(n18523) );
  INVX0 U11792 ( .ZN(n18524), .INP(n18525) );
  INVX0 U11795 ( .ZN(n18526), .INP(n18527) );
  INVX0 U11798 ( .ZN(n18528), .INP(n18529) );
  INVX0 U11801 ( .ZN(n18530), .INP(n18531) );
  INVX0 U11804 ( .ZN(n18532), .INP(n18533) );
  INVX0 U11807 ( .ZN(n18534), .INP(n18535) );
  INVX0 U11810 ( .ZN(n18536), .INP(n18537) );
  INVX0 U11813 ( .ZN(n18538), .INP(n18539) );
  INVX0 U11816 ( .ZN(n18540), .INP(n18541) );
  INVX0 U11823 ( .ZN(n18542), .INP(n18543) );
  INVX0 U11826 ( .ZN(n18544), .INP(n18545) );
  INVX0 U11829 ( .ZN(n18546), .INP(n18547) );
  INVX0 U11832 ( .ZN(n18548), .INP(n18549) );
  INVX0 U11835 ( .ZN(n18550), .INP(n18551) );
  INVX0 U11838 ( .ZN(n18552), .INP(n18553) );
  INVX0 U11841 ( .ZN(n18554), .INP(n18555) );
  INVX0 U11844 ( .ZN(n18556), .INP(n18557) );
  INVX0 U11847 ( .ZN(n18558), .INP(n18559) );
  INVX0 U11848 ( .ZN(n18560), .INP(n18561) );
  INVX0 U11850 ( .ZN(n18562), .INP(n18563) );
  INVX0 U11853 ( .ZN(n18564), .INP(n18565) );
  INVX0 U11856 ( .ZN(n18566), .INP(n18567) );
  INVX0 U11859 ( .ZN(n18568), .INP(n18569) );
  INVX0 U11862 ( .ZN(n18570), .INP(n18571) );
  INVX0 U11865 ( .ZN(n18572), .INP(n18573) );
  INVX0 U11868 ( .ZN(n18574), .INP(n18575) );
  INVX0 U11871 ( .ZN(n18576), .INP(n18577) );
  INVX0 U11874 ( .ZN(n18578), .INP(n18579) );
  INVX0 U11324 ( .ZN(n18211), .INP(n18212) );
  INVX0 U11327 ( .ZN(n18213), .INP(n18214) );
  INVX0 U11330 ( .ZN(n18215), .INP(n18216) );
  INVX0 U11333 ( .ZN(n18217), .INP(n18218) );
  INVX0 U11336 ( .ZN(n18219), .INP(n18220) );
  INVX0 U11339 ( .ZN(n18221), .INP(n18222) );
  INVX0 U11342 ( .ZN(n18223), .INP(n18224) );
  INVX0 U11345 ( .ZN(n18225), .INP(n18226) );
  INVX0 U11348 ( .ZN(n18227), .INP(n18228) );
  INVX0 U11351 ( .ZN(n18229), .INP(n18230) );
  INVX0 U11354 ( .ZN(n18231), .INP(n18232) );
  INVX0 U11357 ( .ZN(n18233), .INP(n18234) );
  INVX0 U11360 ( .ZN(n18235), .INP(n18236) );
  INVX0 U11363 ( .ZN(n18237), .INP(n18238) );
  INVX0 U11366 ( .ZN(n18239), .INP(n18240) );
  INVX0 U11369 ( .ZN(n18241), .INP(n18242) );
  INVX0 U11372 ( .ZN(n18243), .INP(n18244) );
  INVX0 U11375 ( .ZN(n18245), .INP(n18246) );
  INVX0 U11378 ( .ZN(n18247), .INP(n18248) );
  INVX0 U11381 ( .ZN(n18249), .INP(n18250) );
  INVX0 U11384 ( .ZN(n18251), .INP(n18252) );
  INVX0 U11387 ( .ZN(n18253), .INP(n18254) );
  INVX0 U11390 ( .ZN(n18255), .INP(n18256) );
  INVX0 U11393 ( .ZN(n18257), .INP(n18258) );
  INVX0 U11396 ( .ZN(n18259), .INP(n18260) );
  INVX0 U11399 ( .ZN(n18261), .INP(n18262) );
  INVX0 U11402 ( .ZN(n18263), .INP(n18264) );
  INVX0 U11405 ( .ZN(n18265), .INP(n18266) );
  INVX0 U11408 ( .ZN(n18267), .INP(n18268) );
  INVX0 U11411 ( .ZN(n18269), .INP(n18270) );
  INVX0 U11414 ( .ZN(n18271), .INP(n18272) );
  INVX0 U11417 ( .ZN(n18273), .INP(n18274) );
  INVX0 U11420 ( .ZN(n18275), .INP(n18276) );
  INVX0 U11423 ( .ZN(n18277), .INP(n18278) );
  INVX0 U11426 ( .ZN(n18279), .INP(n18280) );
  INVX0 U11429 ( .ZN(n18281), .INP(n18282) );
  INVX0 U11432 ( .ZN(n18283), .INP(N74) );
  INVX0 U11444 ( .ZN(n18289), .INP(n18290) );
  INVX0 U11447 ( .ZN(n18291), .INP(n18292) );
  INVX0 U11450 ( .ZN(n18293), .INP(n18294) );
  INVX0 U11453 ( .ZN(n18295), .INP(N71) );
  INVX0 U11486 ( .ZN(n18316), .INP(n18317) );
  INVX0 U11489 ( .ZN(n18318), .INP(n18319) );
  INVX0 U11492 ( .ZN(n18320), .INP(n18321) );
  INVX0 U11534 ( .ZN(n18348), .INP(n18349) );
  INVX0 U11537 ( .ZN(n18350), .INP(n18351) );
  INVX0 U11540 ( .ZN(n18352), .INP(n18353) );
  INVX0 U11543 ( .ZN(n18354), .INP(n18355) );
  INVX0 U11546 ( .ZN(n18356), .INP(n18357) );
  INVX0 U11549 ( .ZN(n18358), .INP(n18359) );
  INVX0 U11552 ( .ZN(n18360), .INP(n18361) );
  INVX0 U11555 ( .ZN(n18362), .INP(n18363) );
  INVX0 U11558 ( .ZN(n18364), .INP(n18365) );
  INVX0 U11561 ( .ZN(n18366), .INP(n18367) );
  INVX0 U11564 ( .ZN(n18368), .INP(n18369) );
  INVX0 U11567 ( .ZN(n18370), .INP(n18371) );
  INVX0 U11570 ( .ZN(n18372), .INP(n18373) );
  INVX0 U11573 ( .ZN(n18374), .INP(n18375) );
  INVX0 U11576 ( .ZN(n18376), .INP(n18377) );
  INVX0 U11579 ( .ZN(n18378), .INP(n18379) );
  INVX0 U11582 ( .ZN(n18380), .INP(n18381) );
  INVX0 U11585 ( .ZN(n18382), .INP(n18383) );
  INVX0 U11588 ( .ZN(n18384), .INP(n18385) );
  INVX0 U11591 ( .ZN(n18386), .INP(n18387) );
  INVX0 U11594 ( .ZN(n18388), .INP(n18389) );
  INVX0 U11597 ( .ZN(n18390), .INP(n18391) );
  INVX0 U11600 ( .ZN(n18392), .INP(n18393) );
  OR2X1 U19932 ( .IN2(n17624), .IN1(n17623), .Q(n17628) );
  OR2X1 U19933 ( .IN2(n17626), .IN1(n17625), .Q(n17630) );
  OR2X1 U19934 ( .IN2(n17629), .IN1(n17627), .Q(n17634) );
  OR2X1 U19935 ( .IN2(n17633), .IN1(n17631), .Q(n17643) );
  OR2X1 U19936 ( .IN2(n17636), .IN1(n17635), .Q(n17640) );
  OR2X1 U19937 ( .IN2(n17638), .IN1(n17637), .Q(n17642) );
  OR2X1 U19938 ( .IN2(n17641), .IN1(n17639), .Q(n17644) );
  OR2X1 U19939 ( .IN2(n17646), .IN1(n17645), .Q(n17650) );
  OR2X1 U19940 ( .IN2(n17648), .IN1(n17647), .Q(n17652) );
  OR2X1 U19941 ( .IN2(n17651), .IN1(n17649), .Q(n17662) );
  OR2X1 U19942 ( .IN2(n17654), .IN1(n17653), .Q(n17658) );
  OR2X1 U19943 ( .IN2(n17656), .IN1(n17655), .Q(n17660) );
  OR2X1 U19944 ( .IN2(n17659), .IN1(n17657), .Q(n17664) );
  OR2X1 U19945 ( .IN2(n17663), .IN1(n17661), .Q(n17673) );
  OR2X1 U19946 ( .IN2(n17666), .IN1(n17665), .Q(n17670) );
  OR2X1 U19947 ( .IN2(n17668), .IN1(n17667), .Q(n17672) );
  OR2X1 U19948 ( .IN2(n17671), .IN1(n17669), .Q(n17674) );
  OR2X1 U19949 ( .IN2(n17676), .IN1(n17675), .Q(n17680) );
  OR2X1 U19950 ( .IN2(n17678), .IN1(n17677), .Q(n17682) );
  OR2X1 U19951 ( .IN2(n17681), .IN1(n17679), .Q(n17692) );
  OR2X1 U19952 ( .IN2(n17684), .IN1(n17683), .Q(n17688) );
  OR2X1 U19953 ( .IN2(n17686), .IN1(n17685), .Q(n17690) );
  OR2X1 U19954 ( .IN2(n17689), .IN1(n17687), .Q(n17694) );
  OR2X1 U19955 ( .IN2(n17693), .IN1(n17691), .Q(n17703) );
  OR2X1 U19956 ( .IN2(n17696), .IN1(n17695), .Q(n17700) );
  OR2X1 U19957 ( .IN2(n17698), .IN1(n17697), .Q(n17702) );
  OR2X1 U19958 ( .IN2(n17701), .IN1(n17699), .Q(n17704) );
  OR2X1 U19959 ( .IN2(n17706), .IN1(n17705), .Q(n17710) );
  OR2X1 U19960 ( .IN2(n17708), .IN1(n17707), .Q(n17712) );
  OR2X1 U19961 ( .IN2(n17711), .IN1(n17709), .Q(n17722) );
  OR2X1 U19962 ( .IN2(n17714), .IN1(n17713), .Q(n17718) );
  OR2X1 U19963 ( .IN2(n17716), .IN1(n17715), .Q(n17720) );
  OR2X1 U19964 ( .IN2(n17719), .IN1(n17717), .Q(n17724) );
  OR2X1 U19965 ( .IN2(n17723), .IN1(n17721), .Q(n17733) );
  OR2X1 U19966 ( .IN2(n7012), .IN1(n6837), .Q(n17727) );
  OR2X1 U19967 ( .IN2(n6842), .IN1(n7012), .Q(n17726) );
  OR2X1 U19968 ( .IN2(n7012), .IN1(n6813), .Q(n17730) );
  OR2X1 U19969 ( .IN2(n6842), .IN1(n7012), .Q(n17729) );
  OR2X1 U19970 ( .IN2(n17725), .IN1(n6793), .Q(n17732) );
  OR2X1 U19971 ( .IN2(n17728), .IN1(n6784), .Q(n17731) );
  AND2X1 U19974 ( .IN1(n7145), .IN2(n7052), .Q(n17736) );
  NOR2X0 U19975 ( .QN(n17735), .IN1(n7052), .IN2(n7145) );
  NOR2X0 U19976 ( .QN(P1_N5180), .IN1(n17736), .IN2(n17735) );
  AND2X1 U19978 ( .IN1(n7265), .IN2(n7147), .Q(n17738) );
  NOR2X0 U19979 ( .QN(n17737), .IN1(n7147), .IN2(n7265) );
  NOR2X0 U19980 ( .QN(P2_N5102), .IN1(n17738), .IN2(n17737) );
  INVX0 U11295 ( .ZN(n18194), .INP(n1503) );
  INVX0 U11296 ( .ZN(n18195), .INP(n1504) );
  INVX0 U11303 ( .ZN(n18198), .INP(n18199) );
  INVX0 U11306 ( .ZN(n18200), .INP(n18201) );
  INVX0 U11309 ( .ZN(n18202), .INP(n18203) );
  INVX0 U11321 ( .ZN(n18209), .INP(n18210) );
  OR2X1 U19839 ( .IN2(n17346), .IN1(n17345), .Q(n17350) );
  OR2X1 U19840 ( .IN2(n17348), .IN1(n17347), .Q(n17352) );
  OR2X1 U19841 ( .IN2(n17351), .IN1(n17349), .Q(n17362) );
  OR2X1 U19842 ( .IN2(n17354), .IN1(n17353), .Q(n17358) );
  OR2X1 U19843 ( .IN2(n17356), .IN1(n17355), .Q(n17360) );
  OR2X1 U19844 ( .IN2(n17359), .IN1(n17357), .Q(n17364) );
  OR2X1 U19845 ( .IN2(n17363), .IN1(n17361), .Q(n17373) );
  OR2X1 U19846 ( .IN2(n17366), .IN1(n17365), .Q(n17370) );
  OR2X1 U19847 ( .IN2(n17368), .IN1(n17367), .Q(n17372) );
  OR2X1 U19848 ( .IN2(n17371), .IN1(n17369), .Q(n17374) );
  OR2X1 U19849 ( .IN2(n17376), .IN1(n17375), .Q(n17380) );
  OR2X1 U19850 ( .IN2(n17378), .IN1(n17377), .Q(n17382) );
  OR2X1 U19851 ( .IN2(n17381), .IN1(n17379), .Q(n17392) );
  OR2X1 U19852 ( .IN2(n17384), .IN1(n17383), .Q(n17388) );
  OR2X1 U19853 ( .IN2(n17386), .IN1(n17385), .Q(n17390) );
  OR2X1 U19854 ( .IN2(n17389), .IN1(n17387), .Q(n17394) );
  OR2X1 U19855 ( .IN2(n17393), .IN1(n17391), .Q(n17403) );
  OR2X1 U19856 ( .IN2(n17396), .IN1(n17395), .Q(n17400) );
  OR2X1 U19857 ( .IN2(n17398), .IN1(n17397), .Q(n17402) );
  OR2X1 U19858 ( .IN2(n17401), .IN1(n17399), .Q(n17404) );
  OR2X1 U19859 ( .IN2(n17406), .IN1(n17405), .Q(n17410) );
  OR2X1 U19860 ( .IN2(n17408), .IN1(n17407), .Q(n17412) );
  OR2X1 U19861 ( .IN2(n17411), .IN1(n17409), .Q(n17422) );
  OR2X1 U19862 ( .IN2(n17414), .IN1(n17413), .Q(n17418) );
  OR2X1 U19863 ( .IN2(n17416), .IN1(n17415), .Q(n17420) );
  OR2X1 U19864 ( .IN2(n17419), .IN1(n17417), .Q(n17424) );
  OR2X1 U19865 ( .IN2(n17423), .IN1(n17421), .Q(n17433) );
  OR2X1 U19866 ( .IN2(n17426), .IN1(n17425), .Q(n17430) );
  OR2X1 U19867 ( .IN2(n17428), .IN1(n17427), .Q(n17432) );
  OR2X1 U19868 ( .IN2(n17431), .IN1(n17429), .Q(n17434) );
  OR2X1 U19869 ( .IN2(n17436), .IN1(n17435), .Q(n17440) );
  OR2X1 U19870 ( .IN2(n17438), .IN1(n17437), .Q(n17442) );
  OR2X1 U19871 ( .IN2(n17441), .IN1(n17439), .Q(n17452) );
  OR2X1 U19872 ( .IN2(n17444), .IN1(n17443), .Q(n17448) );
  OR2X1 U19873 ( .IN2(n17446), .IN1(n17445), .Q(n17450) );
  OR2X1 U19874 ( .IN2(n17449), .IN1(n17447), .Q(n17454) );
  OR2X1 U19875 ( .IN2(n17453), .IN1(n17451), .Q(n17463) );
  OR2X1 U19876 ( .IN2(n17456), .IN1(n17455), .Q(n17460) );
  OR2X1 U19877 ( .IN2(n17458), .IN1(n17457), .Q(n17462) );
  OR2X1 U19878 ( .IN2(n17461), .IN1(n17459), .Q(n17464) );
  OR2X1 U19879 ( .IN2(n17466), .IN1(n17465), .Q(n17470) );
  OR2X1 U19880 ( .IN2(n17468), .IN1(n17467), .Q(n17472) );
  OR2X1 U19881 ( .IN2(n17471), .IN1(n17469), .Q(n17482) );
  OR2X1 U19882 ( .IN2(n17474), .IN1(n17473), .Q(n17478) );
  OR2X1 U19883 ( .IN2(n17476), .IN1(n17475), .Q(n17480) );
  OR2X1 U19884 ( .IN2(n17479), .IN1(n17477), .Q(n17484) );
  OR2X1 U19885 ( .IN2(n17483), .IN1(n17481), .Q(n17493) );
  OR2X1 U19886 ( .IN2(n17486), .IN1(n17485), .Q(n17490) );
  OR2X1 U19887 ( .IN2(n17488), .IN1(n17487), .Q(n17492) );
  OR2X1 U19888 ( .IN2(n17491), .IN1(n17489), .Q(n17494) );
  OR2X1 U19889 ( .IN2(n17496), .IN1(n17495), .Q(n17500) );
  OR2X1 U19890 ( .IN2(n17498), .IN1(n17497), .Q(n17502) );
  OR2X1 U19891 ( .IN2(n17501), .IN1(n17499), .Q(n17512) );
  OR2X1 U19892 ( .IN2(n17504), .IN1(n17503), .Q(n17508) );
  OR2X1 U19893 ( .IN2(n17506), .IN1(n17505), .Q(n17510) );
  OR2X1 U19894 ( .IN2(n17509), .IN1(n17507), .Q(n17514) );
  OR2X1 U19895 ( .IN2(n17513), .IN1(n17511), .Q(n17523) );
  OR2X1 U19896 ( .IN2(n17516), .IN1(n17515), .Q(n17520) );
  OR2X1 U19897 ( .IN2(n17518), .IN1(n17517), .Q(n17522) );
  OR2X1 U19898 ( .IN2(n17521), .IN1(n17519), .Q(n17524) );
  OR2X1 U19899 ( .IN2(n17526), .IN1(n17525), .Q(n17530) );
  OR2X1 U19900 ( .IN2(n17528), .IN1(n17527), .Q(n17532) );
  OR2X1 U19901 ( .IN2(n17531), .IN1(n17529), .Q(n17542) );
  OR2X1 U19902 ( .IN2(n17534), .IN1(n17533), .Q(n17538) );
  OR2X1 U19903 ( .IN2(n17536), .IN1(n17535), .Q(n17540) );
  OR2X1 U19904 ( .IN2(n17539), .IN1(n17537), .Q(n17544) );
  OR2X1 U19905 ( .IN2(n17543), .IN1(n17541), .Q(n17553) );
  OR2X1 U19906 ( .IN2(n17546), .IN1(n17545), .Q(n17550) );
  OR2X1 U19907 ( .IN2(n17548), .IN1(n17547), .Q(n17552) );
  OR2X1 U19908 ( .IN2(n17551), .IN1(n17549), .Q(n17554) );
  OR2X1 U19909 ( .IN2(n17556), .IN1(n17555), .Q(n17560) );
  OR2X1 U19910 ( .IN2(n17558), .IN1(n17557), .Q(n17562) );
  OR2X1 U19911 ( .IN2(n17561), .IN1(n17559), .Q(n17572) );
  OR2X1 U19912 ( .IN2(n17564), .IN1(n17563), .Q(n17568) );
  OR2X1 U19913 ( .IN2(n17566), .IN1(n17565), .Q(n17570) );
  OR2X1 U19914 ( .IN2(n17569), .IN1(n17567), .Q(n17574) );
  OR2X1 U19915 ( .IN2(n17573), .IN1(n17571), .Q(n17583) );
  OR2X1 U19916 ( .IN2(n17576), .IN1(n17575), .Q(n17580) );
  OR2X1 U19917 ( .IN2(n17578), .IN1(n17577), .Q(n17582) );
  OR2X1 U19918 ( .IN2(n17581), .IN1(n17579), .Q(n17584) );
  OR2X1 U19919 ( .IN2(n17586), .IN1(n17585), .Q(n17590) );
  OR2X1 U19920 ( .IN2(n17588), .IN1(n17587), .Q(n17592) );
  OR2X1 U19921 ( .IN2(n17591), .IN1(n17589), .Q(n17602) );
  OR2X1 U19922 ( .IN2(n17594), .IN1(n17593), .Q(n17598) );
  OR2X1 U19923 ( .IN2(n17596), .IN1(n17595), .Q(n17600) );
  OR2X1 U19924 ( .IN2(n17599), .IN1(n17597), .Q(n17604) );
  OR2X1 U19925 ( .IN2(n17603), .IN1(n17601), .Q(n17613) );
  OR2X1 U19926 ( .IN2(n17606), .IN1(n17605), .Q(n17610) );
  OR2X1 U19927 ( .IN2(n17608), .IN1(n17607), .Q(n17612) );
  OR2X1 U19928 ( .IN2(n17611), .IN1(n17609), .Q(n17614) );
  OR2X1 U19929 ( .IN2(n17616), .IN1(n17615), .Q(n17620) );
  OR2X1 U19930 ( .IN2(n17618), .IN1(n17617), .Q(n17622) );
  OR2X1 U19931 ( .IN2(n17621), .IN1(n17619), .Q(n17632) );
  OR2X1 U19746 ( .IN2(n17065), .IN1(n17064), .Q(n17069) );
  OR2X1 U19747 ( .IN2(n17068), .IN1(n17066), .Q(n17071) );
  OR2X1 U19748 ( .IN2(n17072), .IN1(n17070), .Q(n17074) );
  OR2X1 U19749 ( .IN2(n17076), .IN1(n17075), .Q(n17078) );
  OR2X1 U19750 ( .IN2(n17079), .IN1(n17077), .Q(n17089) );
  OR2X1 U19751 ( .IN2(n17081), .IN1(n17080), .Q(n17085) );
  OR2X1 U19752 ( .IN2(n17083), .IN1(n17082), .Q(n17087) );
  OR2X1 U19753 ( .IN2(n17086), .IN1(n17084), .Q(n17091) );
  OR2X1 U19754 ( .IN2(n17090), .IN1(n17088), .Q(n17103) );
  OR2X1 U19755 ( .IN2(n17093), .IN1(n17092), .Q(n17097) );
  OR2X1 U19756 ( .IN2(n17095), .IN1(n17094), .Q(n17099) );
  OR2X1 U19757 ( .IN2(n17098), .IN1(n17096), .Q(n17101) );
  OR2X1 U19758 ( .IN2(n17102), .IN1(n17100), .Q(n17104) );
  OR2X1 U19759 ( .IN2(n17106), .IN1(n17105), .Q(n17110) );
  OR2X1 U19760 ( .IN2(n17108), .IN1(n17107), .Q(n17112) );
  OR2X1 U19761 ( .IN2(n17111), .IN1(n17109), .Q(n17122) );
  OR2X1 U19762 ( .IN2(n17114), .IN1(n17113), .Q(n17118) );
  OR2X1 U19763 ( .IN2(n17116), .IN1(n17115), .Q(n17120) );
  OR2X1 U19764 ( .IN2(n17119), .IN1(n17117), .Q(n17124) );
  OR2X1 U19765 ( .IN2(n17123), .IN1(n17121), .Q(n17133) );
  OR2X1 U19766 ( .IN2(n17126), .IN1(n17125), .Q(n17130) );
  OR2X1 U19767 ( .IN2(n17128), .IN1(n17127), .Q(n17132) );
  OR2X1 U19768 ( .IN2(n17131), .IN1(n17129), .Q(n17134) );
  OR2X1 U19769 ( .IN2(n17136), .IN1(n17135), .Q(n17140) );
  OR2X1 U19770 ( .IN2(n17138), .IN1(n17137), .Q(n17142) );
  OR2X1 U19771 ( .IN2(n17141), .IN1(n17139), .Q(n17152) );
  OR2X1 U19772 ( .IN2(n17144), .IN1(n17143), .Q(n17148) );
  OR2X1 U19773 ( .IN2(n17146), .IN1(n17145), .Q(n17150) );
  OR2X1 U19774 ( .IN2(n17149), .IN1(n17147), .Q(n17154) );
  OR2X1 U19775 ( .IN2(n17153), .IN1(n17151), .Q(n17163) );
  OR2X1 U19776 ( .IN2(n17156), .IN1(n17155), .Q(n17160) );
  OR2X1 U19777 ( .IN2(n17158), .IN1(n17157), .Q(n17162) );
  OR2X1 U19778 ( .IN2(n17161), .IN1(n17159), .Q(n17164) );
  OR2X1 U19779 ( .IN2(n17166), .IN1(n17165), .Q(n17170) );
  OR2X1 U19780 ( .IN2(n17168), .IN1(n17167), .Q(n17172) );
  OR2X1 U19781 ( .IN2(n17171), .IN1(n17169), .Q(n17182) );
  OR2X1 U19782 ( .IN2(n17174), .IN1(n17173), .Q(n17178) );
  OR2X1 U19783 ( .IN2(n17176), .IN1(n17175), .Q(n17180) );
  OR2X1 U19784 ( .IN2(n17179), .IN1(n17177), .Q(n17184) );
  OR2X1 U19785 ( .IN2(n17183), .IN1(n17181), .Q(n17193) );
  OR2X1 U19786 ( .IN2(n17186), .IN1(n17185), .Q(n17190) );
  OR2X1 U19787 ( .IN2(n17188), .IN1(n17187), .Q(n17192) );
  OR2X1 U19788 ( .IN2(n17191), .IN1(n17189), .Q(n17194) );
  OR2X1 U19789 ( .IN2(n17196), .IN1(n17195), .Q(n17200) );
  OR2X1 U19790 ( .IN2(n17198), .IN1(n17197), .Q(n17202) );
  OR2X1 U19791 ( .IN2(n17201), .IN1(n17199), .Q(n17212) );
  OR2X1 U19792 ( .IN2(n17204), .IN1(n17203), .Q(n17208) );
  OR2X1 U19793 ( .IN2(n17206), .IN1(n17205), .Q(n17210) );
  OR2X1 U19794 ( .IN2(n17209), .IN1(n17207), .Q(n17214) );
  OR2X1 U19795 ( .IN2(n17213), .IN1(n17211), .Q(n17223) );
  OR2X1 U19796 ( .IN2(n17216), .IN1(n17215), .Q(n17220) );
  OR2X1 U19797 ( .IN2(n17218), .IN1(n17217), .Q(n17222) );
  OR2X1 U19798 ( .IN2(n17221), .IN1(n17219), .Q(n17224) );
  OR2X1 U19799 ( .IN2(n17226), .IN1(n17225), .Q(n17230) );
  OR2X1 U19800 ( .IN2(n17228), .IN1(n17227), .Q(n17232) );
  OR2X1 U19801 ( .IN2(n17231), .IN1(n17229), .Q(n17242) );
  OR2X1 U19802 ( .IN2(n17234), .IN1(n17233), .Q(n17238) );
  OR2X1 U19803 ( .IN2(n17236), .IN1(n17235), .Q(n17240) );
  OR2X1 U19804 ( .IN2(n17239), .IN1(n17237), .Q(n17244) );
  OR2X1 U19805 ( .IN2(n17243), .IN1(n17241), .Q(n17253) );
  OR2X1 U19806 ( .IN2(n17246), .IN1(n17245), .Q(n17250) );
  OR2X1 U19807 ( .IN2(n17248), .IN1(n17247), .Q(n17252) );
  OR2X1 U19808 ( .IN2(n17251), .IN1(n17249), .Q(n17254) );
  OR2X1 U19809 ( .IN2(n17256), .IN1(n17255), .Q(n17260) );
  OR2X1 U19810 ( .IN2(n17258), .IN1(n17257), .Q(n17262) );
  OR2X1 U19811 ( .IN2(n17261), .IN1(n17259), .Q(n17272) );
  OR2X1 U19812 ( .IN2(n17264), .IN1(n17263), .Q(n17268) );
  OR2X1 U19813 ( .IN2(n17266), .IN1(n17265), .Q(n17270) );
  OR2X1 U19814 ( .IN2(n17269), .IN1(n17267), .Q(n17274) );
  OR2X1 U19815 ( .IN2(n17273), .IN1(n17271), .Q(n17283) );
  OR2X1 U19816 ( .IN2(n17276), .IN1(n17275), .Q(n17280) );
  OR2X1 U19817 ( .IN2(n17278), .IN1(n17277), .Q(n17282) );
  OR2X1 U19818 ( .IN2(n17281), .IN1(n17279), .Q(n17284) );
  OR2X1 U19819 ( .IN2(n17286), .IN1(n17285), .Q(n17290) );
  OR2X1 U19820 ( .IN2(n17288), .IN1(n17287), .Q(n17292) );
  OR2X1 U19821 ( .IN2(n17291), .IN1(n17289), .Q(n17302) );
  OR2X1 U19822 ( .IN2(n17294), .IN1(n17293), .Q(n17298) );
  OR2X1 U19823 ( .IN2(n17296), .IN1(n17295), .Q(n17300) );
  OR2X1 U19824 ( .IN2(n17299), .IN1(n17297), .Q(n17304) );
  OR2X1 U19825 ( .IN2(n17303), .IN1(n17301), .Q(n17313) );
  OR2X1 U19826 ( .IN2(n17306), .IN1(n17305), .Q(n17310) );
  OR2X1 U19827 ( .IN2(n17308), .IN1(n17307), .Q(n17312) );
  OR2X1 U19828 ( .IN2(n17311), .IN1(n17309), .Q(n17314) );
  OR2X1 U19829 ( .IN2(n17316), .IN1(n17315), .Q(n17320) );
  OR2X1 U19830 ( .IN2(n17318), .IN1(n17317), .Q(n17322) );
  OR2X1 U19831 ( .IN2(n17321), .IN1(n17319), .Q(n17332) );
  OR2X1 U19832 ( .IN2(n17324), .IN1(n17323), .Q(n17328) );
  OR2X1 U19833 ( .IN2(n17326), .IN1(n17325), .Q(n17330) );
  OR2X1 U19834 ( .IN2(n17329), .IN1(n17327), .Q(n17334) );
  OR2X1 U19835 ( .IN2(n17333), .IN1(n17331), .Q(n17343) );
  OR2X1 U19836 ( .IN2(n17336), .IN1(n17335), .Q(n17340) );
  OR2X1 U19837 ( .IN2(n17338), .IN1(n17337), .Q(n17342) );
  OR2X1 U19838 ( .IN2(n17341), .IN1(n17339), .Q(n17344) );
  OR2X1 U19653 ( .IN2(n16786), .IN1(n16784), .Q(n16799) );
  OR2X1 U19654 ( .IN2(n16789), .IN1(n16788), .Q(n16793) );
  OR2X1 U19655 ( .IN2(n16791), .IN1(n16790), .Q(n16795) );
  OR2X1 U19656 ( .IN2(n16794), .IN1(n16792), .Q(n16798) );
  OR2X1 U19657 ( .IN2(n16797), .IN1(n16796), .Q(n16800) );
  OR2X1 U19658 ( .IN2(n16802), .IN1(n16801), .Q(n16806) );
  OR2X1 U19659 ( .IN2(n16804), .IN1(n16803), .Q(n16808) );
  OR2X1 U19660 ( .IN2(n16807), .IN1(n16805), .Q(n16818) );
  OR2X1 U19661 ( .IN2(n16810), .IN1(n16809), .Q(n16814) );
  OR2X1 U19662 ( .IN2(n16812), .IN1(n16811), .Q(n16816) );
  OR2X1 U19663 ( .IN2(n16815), .IN1(n16813), .Q(n16820) );
  OR2X1 U19664 ( .IN2(n16819), .IN1(n16817), .Q(n16832) );
  OR2X1 U19665 ( .IN2(n16822), .IN1(n16821), .Q(n16826) );
  OR2X1 U19666 ( .IN2(n16824), .IN1(n16823), .Q(n16828) );
  OR2X1 U19667 ( .IN2(n16827), .IN1(n16825), .Q(n16831) );
  OR2X1 U19668 ( .IN2(n16830), .IN1(n16829), .Q(n16833) );
  OR2X1 U19669 ( .IN2(n16835), .IN1(n16834), .Q(n16838) );
  OR2X1 U19670 ( .IN2(n16837), .IN1(n16836), .Q(n16839) );
  OR2X1 U19671 ( .IN2(n16841), .IN1(n16840), .Q(n16844) );
  OR2X1 U19672 ( .IN2(n16843), .IN1(n16842), .Q(n16845) );
  OR2X1 U19673 ( .IN2(n16847), .IN1(n16846), .Q(n16850) );
  OR2X1 U19674 ( .IN2(n16849), .IN1(n16848), .Q(n16851) );
  OR2X1 U19675 ( .IN2(n16853), .IN1(n16852), .Q(n16856) );
  OR2X1 U19676 ( .IN2(n16855), .IN1(n16854), .Q(n16857) );
  OR2X1 U19677 ( .IN2(n16859), .IN1(n16858), .Q(n16862) );
  OR2X1 U19678 ( .IN2(n16861), .IN1(n16860), .Q(n16863) );
  OR2X1 U19679 ( .IN2(n16865), .IN1(n16864), .Q(n16868) );
  OR2X1 U19680 ( .IN2(n16867), .IN1(n16866), .Q(n16869) );
  OR2X1 U19681 ( .IN2(n16871), .IN1(n16870), .Q(n16874) );
  OR2X1 U19682 ( .IN2(n16873), .IN1(n16872), .Q(n16875) );
  OR2X1 U19683 ( .IN2(n16877), .IN1(n16876), .Q(n16880) );
  OR2X1 U19684 ( .IN2(n16879), .IN1(n16878), .Q(n16881) );
  OR2X1 U19685 ( .IN2(n16883), .IN1(n16882), .Q(n16886) );
  OR2X1 U19686 ( .IN2(n16885), .IN1(n16884), .Q(n16887) );
  OR2X1 U19687 ( .IN2(n16889), .IN1(n16888), .Q(n16892) );
  OR2X1 U19688 ( .IN2(n16891), .IN1(n16890), .Q(n16893) );
  OR2X1 U19689 ( .IN2(n16895), .IN1(n16894), .Q(n16898) );
  OR2X1 U19690 ( .IN2(n16897), .IN1(n16896), .Q(n16899) );
  OR2X1 U19691 ( .IN2(n16901), .IN1(n16900), .Q(n16904) );
  OR2X1 U19692 ( .IN2(n16903), .IN1(n16902), .Q(n16905) );
  OR2X1 U19693 ( .IN2(n16907), .IN1(n16906), .Q(n16910) );
  OR2X1 U19694 ( .IN2(n16909), .IN1(n16908), .Q(n16911) );
  OR2X1 U19695 ( .IN2(n16913), .IN1(n16912), .Q(n16916) );
  OR2X1 U19696 ( .IN2(n16915), .IN1(n16914), .Q(n16917) );
  OR2X1 U19697 ( .IN2(n16919), .IN1(n16918), .Q(n16922) );
  OR2X1 U19698 ( .IN2(n16921), .IN1(n16920), .Q(n16923) );
  OR2X1 U19699 ( .IN2(n16925), .IN1(n16924), .Q(n16928) );
  OR2X1 U19700 ( .IN2(n16927), .IN1(n16926), .Q(n16929) );
  OR2X1 U19701 ( .IN2(n16931), .IN1(n16930), .Q(n16934) );
  OR2X1 U19702 ( .IN2(n16933), .IN1(n16932), .Q(n16935) );
  OR2X1 U19703 ( .IN2(n16937), .IN1(n16936), .Q(n16940) );
  OR2X1 U19704 ( .IN2(n16939), .IN1(n16938), .Q(n16941) );
  OR2X1 U19705 ( .IN2(n16943), .IN1(n16942), .Q(n16946) );
  OR2X1 U19706 ( .IN2(n16945), .IN1(n16944), .Q(n16947) );
  OR2X1 U19707 ( .IN2(n16949), .IN1(n16948), .Q(n16952) );
  OR2X1 U19708 ( .IN2(n16951), .IN1(n16950), .Q(n16953) );
  OR2X1 U19709 ( .IN2(n16955), .IN1(n16954), .Q(n16958) );
  OR2X1 U19710 ( .IN2(n16957), .IN1(n16956), .Q(n16959) );
  OR2X1 U19711 ( .IN2(n16961), .IN1(n16960), .Q(n16964) );
  OR2X1 U19712 ( .IN2(n16963), .IN1(n16962), .Q(n16965) );
  OR2X1 U19713 ( .IN2(n16967), .IN1(n16966), .Q(n16970) );
  OR2X1 U19714 ( .IN2(n16969), .IN1(n16968), .Q(n16971) );
  OR2X1 U19715 ( .IN2(n16973), .IN1(n16972), .Q(n16976) );
  OR2X1 U19716 ( .IN2(n16975), .IN1(n16974), .Q(n16977) );
  OR2X1 U19717 ( .IN2(n16979), .IN1(n16978), .Q(n16982) );
  OR2X1 U19718 ( .IN2(n16981), .IN1(n16980), .Q(n16983) );
  OR2X1 U19719 ( .IN2(n16985), .IN1(n16984), .Q(n16988) );
  OR2X1 U19720 ( .IN2(n16987), .IN1(n16986), .Q(n16989) );
  OR2X1 U19721 ( .IN2(n16991), .IN1(n16990), .Q(n16994) );
  OR2X1 U19722 ( .IN2(n16993), .IN1(n16992), .Q(n16995) );
  OR2X1 U19723 ( .IN2(n16997), .IN1(n16996), .Q(n17000) );
  OR2X1 U19724 ( .IN2(n16999), .IN1(n16998), .Q(n17001) );
  OR2X1 U19725 ( .IN2(n17003), .IN1(n17002), .Q(n17006) );
  OR2X1 U19726 ( .IN2(n17005), .IN1(n17004), .Q(n17007) );
  OR2X1 U19727 ( .IN2(n17009), .IN1(n17008), .Q(n17012) );
  OR2X1 U19728 ( .IN2(n17011), .IN1(n17010), .Q(n17013) );
  OR2X1 U19729 ( .IN2(n17015), .IN1(n17014), .Q(n17017) );
  OR2X1 U19730 ( .IN2(n17018), .IN1(n17016), .Q(n17029) );
  OR2X1 U19731 ( .IN2(n17021), .IN1(n17020), .Q(n17025) );
  OR2X1 U19732 ( .IN2(n17023), .IN1(n17022), .Q(n17027) );
  OR2X1 U19733 ( .IN2(n17026), .IN1(n17024), .Q(n17031) );
  OR2X1 U19734 ( .IN2(n17030), .IN1(n17028), .Q(n17043) );
  OR2X1 U19735 ( .IN2(n17033), .IN1(n17032), .Q(n17037) );
  OR2X1 U19736 ( .IN2(n17035), .IN1(n17034), .Q(n17039) );
  OR2X1 U19737 ( .IN2(n17038), .IN1(n17036), .Q(n17041) );
  OR2X1 U19738 ( .IN2(n17042), .IN1(n17040), .Q(n17044) );
  OR2X1 U19739 ( .IN2(n17046), .IN1(n17045), .Q(n17048) );
  OR2X1 U19740 ( .IN2(n17049), .IN1(n17047), .Q(n17059) );
  OR2X1 U19741 ( .IN2(n17051), .IN1(n17050), .Q(n17055) );
  OR2X1 U19742 ( .IN2(n17053), .IN1(n17052), .Q(n17057) );
  OR2X1 U19743 ( .IN2(n17056), .IN1(n17054), .Q(n17061) );
  OR2X1 U19744 ( .IN2(n17060), .IN1(n17058), .Q(n17073) );
  OR2X1 U19745 ( .IN2(n17063), .IN1(n17062), .Q(n17067) );
  OR2X1 U19560 ( .IN2(n16507), .IN1(n16506), .Q(n16511) );
  OR2X1 U19561 ( .IN2(n16510), .IN1(n16508), .Q(n16521) );
  OR2X1 U19562 ( .IN2(n16513), .IN1(n16512), .Q(n16517) );
  OR2X1 U19563 ( .IN2(n16515), .IN1(n16514), .Q(n16519) );
  OR2X1 U19564 ( .IN2(n16518), .IN1(n16516), .Q(n16523) );
  OR2X1 U19565 ( .IN2(n16522), .IN1(n16520), .Q(n16535) );
  OR2X1 U19566 ( .IN2(n16525), .IN1(n16524), .Q(n16529) );
  OR2X1 U19567 ( .IN2(n16527), .IN1(n16526), .Q(n16531) );
  OR2X1 U19568 ( .IN2(n16530), .IN1(n16528), .Q(n16534) );
  OR2X1 U19569 ( .IN2(n16533), .IN1(n16532), .Q(n16536) );
  OR2X1 U19570 ( .IN2(n16538), .IN1(n16537), .Q(n16542) );
  OR2X1 U19571 ( .IN2(n16540), .IN1(n16539), .Q(n16544) );
  OR2X1 U19572 ( .IN2(n16543), .IN1(n16541), .Q(n16554) );
  OR2X1 U19573 ( .IN2(n16546), .IN1(n16545), .Q(n16550) );
  OR2X1 U19574 ( .IN2(n16548), .IN1(n16547), .Q(n16552) );
  OR2X1 U19575 ( .IN2(n16551), .IN1(n16549), .Q(n16556) );
  OR2X1 U19576 ( .IN2(n16555), .IN1(n16553), .Q(n16568) );
  OR2X1 U19577 ( .IN2(n16558), .IN1(n16557), .Q(n16562) );
  OR2X1 U19578 ( .IN2(n16560), .IN1(n16559), .Q(n16564) );
  OR2X1 U19579 ( .IN2(n16563), .IN1(n16561), .Q(n16567) );
  OR2X1 U19580 ( .IN2(n16566), .IN1(n16565), .Q(n16569) );
  OR2X1 U19581 ( .IN2(n16571), .IN1(n16570), .Q(n16575) );
  OR2X1 U19582 ( .IN2(n16573), .IN1(n16572), .Q(n16577) );
  OR2X1 U19583 ( .IN2(n16576), .IN1(n16574), .Q(n16587) );
  OR2X1 U19584 ( .IN2(n16579), .IN1(n16578), .Q(n16583) );
  OR2X1 U19585 ( .IN2(n16581), .IN1(n16580), .Q(n16585) );
  OR2X1 U19586 ( .IN2(n16584), .IN1(n16582), .Q(n16589) );
  OR2X1 U19587 ( .IN2(n16588), .IN1(n16586), .Q(n16601) );
  OR2X1 U19588 ( .IN2(n16591), .IN1(n16590), .Q(n16595) );
  OR2X1 U19589 ( .IN2(n16593), .IN1(n16592), .Q(n16597) );
  OR2X1 U19590 ( .IN2(n16596), .IN1(n16594), .Q(n16600) );
  OR2X1 U19591 ( .IN2(n16599), .IN1(n16598), .Q(n16602) );
  OR2X1 U19592 ( .IN2(n16604), .IN1(n16603), .Q(n16608) );
  OR2X1 U19593 ( .IN2(n16606), .IN1(n16605), .Q(n16610) );
  OR2X1 U19594 ( .IN2(n16609), .IN1(n16607), .Q(n16620) );
  OR2X1 U19595 ( .IN2(n16612), .IN1(n16611), .Q(n16616) );
  OR2X1 U19596 ( .IN2(n16614), .IN1(n16613), .Q(n16618) );
  OR2X1 U19597 ( .IN2(n16617), .IN1(n16615), .Q(n16622) );
  OR2X1 U19598 ( .IN2(n16621), .IN1(n16619), .Q(n16634) );
  OR2X1 U19599 ( .IN2(n16624), .IN1(n16623), .Q(n16628) );
  OR2X1 U19600 ( .IN2(n16626), .IN1(n16625), .Q(n16630) );
  OR2X1 U19601 ( .IN2(n16629), .IN1(n16627), .Q(n16633) );
  OR2X1 U19602 ( .IN2(n16632), .IN1(n16631), .Q(n16635) );
  OR2X1 U19603 ( .IN2(n16637), .IN1(n16636), .Q(n16641) );
  OR2X1 U19604 ( .IN2(n16639), .IN1(n16638), .Q(n16643) );
  OR2X1 U19605 ( .IN2(n16642), .IN1(n16640), .Q(n16653) );
  OR2X1 U19606 ( .IN2(n16645), .IN1(n16644), .Q(n16649) );
  OR2X1 U19607 ( .IN2(n16647), .IN1(n16646), .Q(n16651) );
  OR2X1 U19608 ( .IN2(n16650), .IN1(n16648), .Q(n16655) );
  OR2X1 U19609 ( .IN2(n16654), .IN1(n16652), .Q(n16667) );
  OR2X1 U19610 ( .IN2(n16657), .IN1(n16656), .Q(n16661) );
  OR2X1 U19611 ( .IN2(n16659), .IN1(n16658), .Q(n16663) );
  OR2X1 U19612 ( .IN2(n16662), .IN1(n16660), .Q(n16666) );
  OR2X1 U19613 ( .IN2(n16665), .IN1(n16664), .Q(n16668) );
  OR2X1 U19614 ( .IN2(n16670), .IN1(n16669), .Q(n16674) );
  OR2X1 U19615 ( .IN2(n16672), .IN1(n16671), .Q(n16676) );
  OR2X1 U19616 ( .IN2(n16675), .IN1(n16673), .Q(n16686) );
  OR2X1 U19617 ( .IN2(n16678), .IN1(n16677), .Q(n16682) );
  OR2X1 U19618 ( .IN2(n16680), .IN1(n16679), .Q(n16684) );
  OR2X1 U19619 ( .IN2(n16683), .IN1(n16681), .Q(n16688) );
  OR2X1 U19620 ( .IN2(n16687), .IN1(n16685), .Q(n16700) );
  OR2X1 U19621 ( .IN2(n16690), .IN1(n16689), .Q(n16694) );
  OR2X1 U19622 ( .IN2(n16692), .IN1(n16691), .Q(n16696) );
  OR2X1 U19623 ( .IN2(n16695), .IN1(n16693), .Q(n16699) );
  OR2X1 U19624 ( .IN2(n16698), .IN1(n16697), .Q(n16701) );
  OR2X1 U19625 ( .IN2(n16703), .IN1(n16702), .Q(n16707) );
  OR2X1 U19626 ( .IN2(n16705), .IN1(n16704), .Q(n16709) );
  OR2X1 U19627 ( .IN2(n16708), .IN1(n16706), .Q(n16719) );
  OR2X1 U19628 ( .IN2(n16711), .IN1(n16710), .Q(n16715) );
  OR2X1 U19629 ( .IN2(n16713), .IN1(n16712), .Q(n16717) );
  OR2X1 U19630 ( .IN2(n16716), .IN1(n16714), .Q(n16721) );
  OR2X1 U19631 ( .IN2(n16720), .IN1(n16718), .Q(n16733) );
  OR2X1 U19632 ( .IN2(n16723), .IN1(n16722), .Q(n16727) );
  OR2X1 U19633 ( .IN2(n16725), .IN1(n16724), .Q(n16729) );
  OR2X1 U19634 ( .IN2(n16728), .IN1(n16726), .Q(n16732) );
  OR2X1 U19635 ( .IN2(n16731), .IN1(n16730), .Q(n16734) );
  OR2X1 U19636 ( .IN2(n16736), .IN1(n16735), .Q(n16740) );
  OR2X1 U19637 ( .IN2(n16738), .IN1(n16737), .Q(n16742) );
  OR2X1 U19638 ( .IN2(n16741), .IN1(n16739), .Q(n16752) );
  OR2X1 U19639 ( .IN2(n16744), .IN1(n16743), .Q(n16748) );
  OR2X1 U19640 ( .IN2(n16746), .IN1(n16745), .Q(n16750) );
  OR2X1 U19641 ( .IN2(n16749), .IN1(n16747), .Q(n16754) );
  OR2X1 U19642 ( .IN2(n16753), .IN1(n16751), .Q(n16766) );
  OR2X1 U19643 ( .IN2(n16756), .IN1(n16755), .Q(n16760) );
  OR2X1 U19644 ( .IN2(n16758), .IN1(n16757), .Q(n16762) );
  OR2X1 U19645 ( .IN2(n16761), .IN1(n16759), .Q(n16765) );
  OR2X1 U19646 ( .IN2(n16764), .IN1(n16763), .Q(n16767) );
  OR2X1 U19647 ( .IN2(n16769), .IN1(n16768), .Q(n16773) );
  OR2X1 U19648 ( .IN2(n16771), .IN1(n16770), .Q(n16775) );
  OR2X1 U19649 ( .IN2(n16774), .IN1(n16772), .Q(n16785) );
  OR2X1 U19650 ( .IN2(n16777), .IN1(n16776), .Q(n16781) );
  OR2X1 U19651 ( .IN2(n16779), .IN1(n16778), .Q(n16783) );
  OR2X1 U19652 ( .IN2(n16782), .IN1(n16780), .Q(n16787) );
  OR2X1 U19467 ( .IN2(n16228), .IN1(n16227), .Q(n16232) );
  OR2X1 U19468 ( .IN2(n16230), .IN1(n16229), .Q(n16234) );
  OR2X1 U19469 ( .IN2(n16233), .IN1(n16231), .Q(n16237) );
  OR2X1 U19470 ( .IN2(n16236), .IN1(n16235), .Q(n16239) );
  OR2X1 U19471 ( .IN2(n16241), .IN1(n16240), .Q(n16245) );
  OR2X1 U19472 ( .IN2(n16243), .IN1(n16242), .Q(n16247) );
  OR2X1 U19473 ( .IN2(n16246), .IN1(n16244), .Q(n16257) );
  OR2X1 U19474 ( .IN2(n16249), .IN1(n16248), .Q(n16253) );
  OR2X1 U19475 ( .IN2(n16251), .IN1(n16250), .Q(n16255) );
  OR2X1 U19476 ( .IN2(n16254), .IN1(n16252), .Q(n16259) );
  OR2X1 U19477 ( .IN2(n16258), .IN1(n16256), .Q(n16271) );
  OR2X1 U19478 ( .IN2(n16261), .IN1(n16260), .Q(n16265) );
  OR2X1 U19479 ( .IN2(n16263), .IN1(n16262), .Q(n16267) );
  OR2X1 U19480 ( .IN2(n16266), .IN1(n16264), .Q(n16270) );
  OR2X1 U19481 ( .IN2(n16269), .IN1(n16268), .Q(n16272) );
  OR2X1 U19482 ( .IN2(n16274), .IN1(n16273), .Q(n16278) );
  OR2X1 U19483 ( .IN2(n16276), .IN1(n16275), .Q(n16280) );
  OR2X1 U19484 ( .IN2(n16279), .IN1(n16277), .Q(n16290) );
  OR2X1 U19485 ( .IN2(n16282), .IN1(n16281), .Q(n16286) );
  OR2X1 U19486 ( .IN2(n16284), .IN1(n16283), .Q(n16288) );
  OR2X1 U19487 ( .IN2(n16287), .IN1(n16285), .Q(n16292) );
  OR2X1 U19488 ( .IN2(n16291), .IN1(n16289), .Q(n16304) );
  OR2X1 U19489 ( .IN2(n16294), .IN1(n16293), .Q(n16298) );
  OR2X1 U19490 ( .IN2(n16296), .IN1(n16295), .Q(n16300) );
  OR2X1 U19491 ( .IN2(n16299), .IN1(n16297), .Q(n16303) );
  OR2X1 U19492 ( .IN2(n16302), .IN1(n16301), .Q(n16305) );
  OR2X1 U19493 ( .IN2(n16307), .IN1(n16306), .Q(n16311) );
  OR2X1 U19494 ( .IN2(n16309), .IN1(n16308), .Q(n16313) );
  OR2X1 U19495 ( .IN2(n16312), .IN1(n16310), .Q(n16323) );
  OR2X1 U19496 ( .IN2(n16315), .IN1(n16314), .Q(n16319) );
  OR2X1 U19497 ( .IN2(n16317), .IN1(n16316), .Q(n16321) );
  OR2X1 U19498 ( .IN2(n16320), .IN1(n16318), .Q(n16325) );
  OR2X1 U19499 ( .IN2(n16324), .IN1(n16322), .Q(n16337) );
  OR2X1 U19500 ( .IN2(n16327), .IN1(n16326), .Q(n16331) );
  OR2X1 U19501 ( .IN2(n16329), .IN1(n16328), .Q(n16333) );
  OR2X1 U19502 ( .IN2(n16332), .IN1(n16330), .Q(n16336) );
  OR2X1 U19503 ( .IN2(n16335), .IN1(n16334), .Q(n16338) );
  OR2X1 U19504 ( .IN2(n16340), .IN1(n16339), .Q(n16344) );
  OR2X1 U19505 ( .IN2(n16342), .IN1(n16341), .Q(n16346) );
  OR2X1 U19506 ( .IN2(n16345), .IN1(n16343), .Q(n16356) );
  OR2X1 U19507 ( .IN2(n16348), .IN1(n16347), .Q(n16352) );
  OR2X1 U19508 ( .IN2(n16350), .IN1(n16349), .Q(n16354) );
  OR2X1 U19509 ( .IN2(n16353), .IN1(n16351), .Q(n16358) );
  OR2X1 U19510 ( .IN2(n16357), .IN1(n16355), .Q(n16370) );
  OR2X1 U19511 ( .IN2(n16360), .IN1(n16359), .Q(n16364) );
  OR2X1 U19512 ( .IN2(n16362), .IN1(n16361), .Q(n16366) );
  OR2X1 U19513 ( .IN2(n16365), .IN1(n16363), .Q(n16369) );
  OR2X1 U19514 ( .IN2(n16368), .IN1(n16367), .Q(n16371) );
  OR2X1 U19515 ( .IN2(n16373), .IN1(n16372), .Q(n16377) );
  OR2X1 U19516 ( .IN2(n16375), .IN1(n16374), .Q(n16379) );
  OR2X1 U19517 ( .IN2(n16378), .IN1(n16376), .Q(n16389) );
  OR2X1 U19518 ( .IN2(n16381), .IN1(n16380), .Q(n16385) );
  OR2X1 U19519 ( .IN2(n16383), .IN1(n16382), .Q(n16387) );
  OR2X1 U19520 ( .IN2(n16386), .IN1(n16384), .Q(n16391) );
  OR2X1 U19521 ( .IN2(n16390), .IN1(n16388), .Q(n16403) );
  OR2X1 U19522 ( .IN2(n16393), .IN1(n16392), .Q(n16397) );
  OR2X1 U19523 ( .IN2(n16395), .IN1(n16394), .Q(n16399) );
  OR2X1 U19524 ( .IN2(n16398), .IN1(n16396), .Q(n16402) );
  OR2X1 U19525 ( .IN2(n16401), .IN1(n16400), .Q(n16404) );
  OR2X1 U19526 ( .IN2(n16406), .IN1(n16405), .Q(n16410) );
  OR2X1 U19527 ( .IN2(n16408), .IN1(n16407), .Q(n16412) );
  OR2X1 U19528 ( .IN2(n16411), .IN1(n16409), .Q(n16422) );
  OR2X1 U19529 ( .IN2(n16414), .IN1(n16413), .Q(n16418) );
  OR2X1 U19530 ( .IN2(n16416), .IN1(n16415), .Q(n16420) );
  OR2X1 U19531 ( .IN2(n16419), .IN1(n16417), .Q(n16424) );
  OR2X1 U19532 ( .IN2(n16423), .IN1(n16421), .Q(n16436) );
  OR2X1 U19533 ( .IN2(n16426), .IN1(n16425), .Q(n16430) );
  OR2X1 U19534 ( .IN2(n16428), .IN1(n16427), .Q(n16432) );
  OR2X1 U19535 ( .IN2(n16431), .IN1(n16429), .Q(n16435) );
  OR2X1 U19536 ( .IN2(n16434), .IN1(n16433), .Q(n16437) );
  OR2X1 U19537 ( .IN2(n16439), .IN1(n16438), .Q(n16443) );
  OR2X1 U19538 ( .IN2(n16441), .IN1(n16440), .Q(n16445) );
  OR2X1 U19539 ( .IN2(n16444), .IN1(n16442), .Q(n16455) );
  OR2X1 U19540 ( .IN2(n16447), .IN1(n16446), .Q(n16451) );
  OR2X1 U19541 ( .IN2(n16449), .IN1(n16448), .Q(n16453) );
  OR2X1 U19542 ( .IN2(n16452), .IN1(n16450), .Q(n16457) );
  OR2X1 U19543 ( .IN2(n16456), .IN1(n16454), .Q(n16469) );
  OR2X1 U19544 ( .IN2(n16459), .IN1(n16458), .Q(n16463) );
  OR2X1 U19545 ( .IN2(n16461), .IN1(n16460), .Q(n16465) );
  OR2X1 U19546 ( .IN2(n16464), .IN1(n16462), .Q(n16468) );
  OR2X1 U19547 ( .IN2(n16467), .IN1(n16466), .Q(n16470) );
  OR2X1 U19548 ( .IN2(n16472), .IN1(n16471), .Q(n16476) );
  OR2X1 U19549 ( .IN2(n16474), .IN1(n16473), .Q(n16478) );
  OR2X1 U19550 ( .IN2(n16477), .IN1(n16475), .Q(n16488) );
  OR2X1 U19551 ( .IN2(n16480), .IN1(n16479), .Q(n16484) );
  OR2X1 U19552 ( .IN2(n16482), .IN1(n16481), .Q(n16486) );
  OR2X1 U19553 ( .IN2(n16485), .IN1(n16483), .Q(n16490) );
  OR2X1 U19554 ( .IN2(n16489), .IN1(n16487), .Q(n16502) );
  OR2X1 U19555 ( .IN2(n16492), .IN1(n16491), .Q(n16496) );
  OR2X1 U19556 ( .IN2(n16494), .IN1(n16493), .Q(n16498) );
  OR2X1 U19557 ( .IN2(n16497), .IN1(n16495), .Q(n16501) );
  OR2X1 U19558 ( .IN2(n16500), .IN1(n16499), .Q(n16503) );
  OR2X1 U19559 ( .IN2(n16505), .IN1(n16504), .Q(n16509) );
  OR2X1 U19374 ( .IN2(n15949), .IN1(n15947), .Q(n15960) );
  OR2X1 U19375 ( .IN2(n15952), .IN1(n15951), .Q(n15956) );
  OR2X1 U19376 ( .IN2(n15954), .IN1(n15953), .Q(n15958) );
  OR2X1 U19377 ( .IN2(n15957), .IN1(n15955), .Q(n15962) );
  OR2X1 U19378 ( .IN2(n15961), .IN1(n15959), .Q(n15974) );
  OR2X1 U19379 ( .IN2(n15964), .IN1(n15963), .Q(n15968) );
  OR2X1 U19380 ( .IN2(n15966), .IN1(n15965), .Q(n15970) );
  OR2X1 U19381 ( .IN2(n15969), .IN1(n15967), .Q(n15973) );
  OR2X1 U19382 ( .IN2(n15972), .IN1(n15971), .Q(n15975) );
  OR2X1 U19383 ( .IN2(n15977), .IN1(n15976), .Q(n15981) );
  OR2X1 U19384 ( .IN2(n15979), .IN1(n15978), .Q(n15983) );
  OR2X1 U19385 ( .IN2(n15982), .IN1(n15980), .Q(n15993) );
  OR2X1 U19386 ( .IN2(n15985), .IN1(n15984), .Q(n15989) );
  OR2X1 U19387 ( .IN2(n15987), .IN1(n15986), .Q(n15991) );
  OR2X1 U19388 ( .IN2(n15990), .IN1(n15988), .Q(n15995) );
  OR2X1 U19389 ( .IN2(n15994), .IN1(n15992), .Q(n16007) );
  OR2X1 U19390 ( .IN2(n15997), .IN1(n15996), .Q(n16001) );
  OR2X1 U19391 ( .IN2(n15999), .IN1(n15998), .Q(n16003) );
  OR2X1 U19392 ( .IN2(n16002), .IN1(n16000), .Q(n16006) );
  OR2X1 U19393 ( .IN2(n16005), .IN1(n16004), .Q(n16008) );
  OR2X1 U19394 ( .IN2(n16010), .IN1(n16009), .Q(n16014) );
  OR2X1 U19395 ( .IN2(n16012), .IN1(n16011), .Q(n16016) );
  OR2X1 U19396 ( .IN2(n16015), .IN1(n16013), .Q(n16026) );
  OR2X1 U19397 ( .IN2(n16018), .IN1(n16017), .Q(n16022) );
  OR2X1 U19398 ( .IN2(n16020), .IN1(n16019), .Q(n16024) );
  OR2X1 U19399 ( .IN2(n16023), .IN1(n16021), .Q(n16028) );
  OR2X1 U19400 ( .IN2(n16027), .IN1(n16025), .Q(n16040) );
  OR2X1 U19401 ( .IN2(n16030), .IN1(n16029), .Q(n16034) );
  OR2X1 U19402 ( .IN2(n16032), .IN1(n16031), .Q(n16036) );
  OR2X1 U19403 ( .IN2(n16035), .IN1(n16033), .Q(n16039) );
  OR2X1 U19404 ( .IN2(n16038), .IN1(n16037), .Q(n16041) );
  OR2X1 U19405 ( .IN2(n16043), .IN1(n16042), .Q(n16047) );
  OR2X1 U19406 ( .IN2(n16045), .IN1(n16044), .Q(n16049) );
  OR2X1 U19407 ( .IN2(n16048), .IN1(n16046), .Q(n16059) );
  OR2X1 U19408 ( .IN2(n16051), .IN1(n16050), .Q(n16055) );
  OR2X1 U19409 ( .IN2(n16053), .IN1(n16052), .Q(n16057) );
  OR2X1 U19410 ( .IN2(n16056), .IN1(n16054), .Q(n16061) );
  OR2X1 U19411 ( .IN2(n16060), .IN1(n16058), .Q(n16073) );
  OR2X1 U19412 ( .IN2(n16063), .IN1(n16062), .Q(n16067) );
  OR2X1 U19413 ( .IN2(n16065), .IN1(n16064), .Q(n16069) );
  OR2X1 U19414 ( .IN2(n16068), .IN1(n16066), .Q(n16072) );
  OR2X1 U19415 ( .IN2(n16071), .IN1(n16070), .Q(n16074) );
  OR2X1 U19416 ( .IN2(n16076), .IN1(n16075), .Q(n16080) );
  OR2X1 U19417 ( .IN2(n16078), .IN1(n16077), .Q(n16082) );
  OR2X1 U19418 ( .IN2(n16081), .IN1(n16079), .Q(n16092) );
  OR2X1 U19419 ( .IN2(n16084), .IN1(n16083), .Q(n16088) );
  OR2X1 U19420 ( .IN2(n16086), .IN1(n16085), .Q(n16090) );
  OR2X1 U19421 ( .IN2(n16089), .IN1(n16087), .Q(n16094) );
  OR2X1 U19422 ( .IN2(n16093), .IN1(n16091), .Q(n16106) );
  OR2X1 U19423 ( .IN2(n16096), .IN1(n16095), .Q(n16100) );
  OR2X1 U19424 ( .IN2(n16098), .IN1(n16097), .Q(n16102) );
  OR2X1 U19425 ( .IN2(n16101), .IN1(n16099), .Q(n16105) );
  OR2X1 U19426 ( .IN2(n16104), .IN1(n16103), .Q(n16107) );
  OR2X1 U19427 ( .IN2(n16109), .IN1(n16108), .Q(n16113) );
  OR2X1 U19428 ( .IN2(n16111), .IN1(n16110), .Q(n16115) );
  OR2X1 U19429 ( .IN2(n16114), .IN1(n16112), .Q(n16125) );
  OR2X1 U19430 ( .IN2(n16117), .IN1(n16116), .Q(n16121) );
  OR2X1 U19431 ( .IN2(n16119), .IN1(n16118), .Q(n16123) );
  OR2X1 U19432 ( .IN2(n16122), .IN1(n16120), .Q(n16127) );
  OR2X1 U19433 ( .IN2(n16126), .IN1(n16124), .Q(n16139) );
  OR2X1 U19434 ( .IN2(n16129), .IN1(n16128), .Q(n16133) );
  OR2X1 U19435 ( .IN2(n16131), .IN1(n16130), .Q(n16135) );
  OR2X1 U19436 ( .IN2(n16134), .IN1(n16132), .Q(n16138) );
  OR2X1 U19437 ( .IN2(n16137), .IN1(n16136), .Q(n16140) );
  OR2X1 U19438 ( .IN2(n16142), .IN1(n16141), .Q(n16146) );
  OR2X1 U19439 ( .IN2(n16144), .IN1(n16143), .Q(n16148) );
  OR2X1 U19440 ( .IN2(n16147), .IN1(n16145), .Q(n16158) );
  OR2X1 U19441 ( .IN2(n16150), .IN1(n16149), .Q(n16154) );
  OR2X1 U19442 ( .IN2(n16152), .IN1(n16151), .Q(n16156) );
  OR2X1 U19443 ( .IN2(n16155), .IN1(n16153), .Q(n16160) );
  OR2X1 U19444 ( .IN2(n16159), .IN1(n16157), .Q(n16172) );
  OR2X1 U19445 ( .IN2(n16162), .IN1(n16161), .Q(n16166) );
  OR2X1 U19446 ( .IN2(n16164), .IN1(n16163), .Q(n16168) );
  OR2X1 U19447 ( .IN2(n16167), .IN1(n16165), .Q(n16171) );
  OR2X1 U19448 ( .IN2(n16170), .IN1(n16169), .Q(n16173) );
  OR2X1 U19449 ( .IN2(n16175), .IN1(n16174), .Q(n16179) );
  OR2X1 U19450 ( .IN2(n16177), .IN1(n16176), .Q(n16181) );
  OR2X1 U19451 ( .IN2(n16180), .IN1(n16178), .Q(n16191) );
  OR2X1 U19452 ( .IN2(n16183), .IN1(n16182), .Q(n16187) );
  OR2X1 U19453 ( .IN2(n16185), .IN1(n16184), .Q(n16189) );
  OR2X1 U19454 ( .IN2(n16188), .IN1(n16186), .Q(n16193) );
  OR2X1 U19455 ( .IN2(n16192), .IN1(n16190), .Q(n16205) );
  OR2X1 U19456 ( .IN2(n16195), .IN1(n16194), .Q(n16199) );
  OR2X1 U19457 ( .IN2(n16197), .IN1(n16196), .Q(n16201) );
  OR2X1 U19458 ( .IN2(n16200), .IN1(n16198), .Q(n16204) );
  OR2X1 U19459 ( .IN2(n16203), .IN1(n16202), .Q(n16206) );
  OR2X1 U19460 ( .IN2(n16208), .IN1(n16207), .Q(n16212) );
  OR2X1 U19461 ( .IN2(n16210), .IN1(n16209), .Q(n16214) );
  OR2X1 U19462 ( .IN2(n16213), .IN1(n16211), .Q(n16224) );
  OR2X1 U19463 ( .IN2(n16216), .IN1(n16215), .Q(n16220) );
  OR2X1 U19464 ( .IN2(n16218), .IN1(n16217), .Q(n16222) );
  OR2X1 U19465 ( .IN2(n16221), .IN1(n16219), .Q(n16226) );
  OR2X1 U19466 ( .IN2(n16225), .IN1(n16223), .Q(n16238) );
  OR2X1 U19281 ( .IN2(n15670), .IN1(n15668), .Q(n15681) );
  OR2X1 U19282 ( .IN2(n15673), .IN1(n15672), .Q(n15677) );
  OR2X1 U19283 ( .IN2(n15675), .IN1(n15674), .Q(n15679) );
  OR2X1 U19284 ( .IN2(n15678), .IN1(n15676), .Q(n15683) );
  OR2X1 U19285 ( .IN2(n15682), .IN1(n15680), .Q(n15698) );
  OR2X1 U19286 ( .IN2(n15685), .IN1(n15684), .Q(n15689) );
  OR2X1 U19287 ( .IN2(n15687), .IN1(n15686), .Q(n15691) );
  OR2X1 U19288 ( .IN2(n15690), .IN1(n15688), .Q(n15695) );
  OR2X1 U19289 ( .IN2(n15693), .IN1(n15692), .Q(n15697) );
  OR2X1 U19290 ( .IN2(n15696), .IN1(n15694), .Q(n15699) );
  OR2X1 U19291 ( .IN2(n15701), .IN1(n15700), .Q(n15705) );
  OR2X1 U19292 ( .IN2(n15703), .IN1(n15702), .Q(n15707) );
  OR2X1 U19293 ( .IN2(n15706), .IN1(n15704), .Q(n15717) );
  OR2X1 U19294 ( .IN2(n15709), .IN1(n15708), .Q(n15713) );
  OR2X1 U19295 ( .IN2(n15711), .IN1(n15710), .Q(n15715) );
  OR2X1 U19296 ( .IN2(n15714), .IN1(n15712), .Q(n15719) );
  OR2X1 U19297 ( .IN2(n15718), .IN1(n15716), .Q(n15734) );
  OR2X1 U19298 ( .IN2(n15721), .IN1(n15720), .Q(n15725) );
  OR2X1 U19299 ( .IN2(n15723), .IN1(n15722), .Q(n15727) );
  OR2X1 U19300 ( .IN2(n15726), .IN1(n15724), .Q(n15731) );
  OR2X1 U19301 ( .IN2(n15729), .IN1(n15728), .Q(n15733) );
  OR2X1 U19302 ( .IN2(n15732), .IN1(n15730), .Q(n15735) );
  OR2X1 U19303 ( .IN2(n15737), .IN1(n15736), .Q(n15741) );
  OR2X1 U19304 ( .IN2(n15739), .IN1(n15738), .Q(n15743) );
  OR2X1 U19305 ( .IN2(n15742), .IN1(n15740), .Q(n15753) );
  OR2X1 U19306 ( .IN2(n15745), .IN1(n15744), .Q(n15749) );
  OR2X1 U19307 ( .IN2(n15747), .IN1(n15746), .Q(n15751) );
  OR2X1 U19308 ( .IN2(n15750), .IN1(n15748), .Q(n15755) );
  OR2X1 U19309 ( .IN2(n15754), .IN1(n15752), .Q(n15770) );
  OR2X1 U19310 ( .IN2(n15757), .IN1(n15756), .Q(n15761) );
  OR2X1 U19311 ( .IN2(n15759), .IN1(n15758), .Q(n15763) );
  OR2X1 U19312 ( .IN2(n15762), .IN1(n15760), .Q(n15767) );
  OR2X1 U19313 ( .IN2(n15765), .IN1(n15764), .Q(n15769) );
  OR2X1 U19314 ( .IN2(n15768), .IN1(n15766), .Q(n15771) );
  OR2X1 U19315 ( .IN2(n15773), .IN1(n15772), .Q(n15777) );
  OR2X1 U19316 ( .IN2(n15775), .IN1(n15774), .Q(n15779) );
  OR2X1 U19317 ( .IN2(n15778), .IN1(n15776), .Q(n15789) );
  OR2X1 U19318 ( .IN2(n15781), .IN1(n15780), .Q(n15785) );
  OR2X1 U19319 ( .IN2(n15783), .IN1(n15782), .Q(n15787) );
  OR2X1 U19320 ( .IN2(n15786), .IN1(n15784), .Q(n15791) );
  OR2X1 U19321 ( .IN2(n15790), .IN1(n15788), .Q(n15806) );
  OR2X1 U19322 ( .IN2(n15793), .IN1(n15792), .Q(n15797) );
  OR2X1 U19323 ( .IN2(n15795), .IN1(n15794), .Q(n15799) );
  OR2X1 U19324 ( .IN2(n15798), .IN1(n15796), .Q(n15803) );
  OR2X1 U19325 ( .IN2(n15801), .IN1(n15800), .Q(n15805) );
  OR2X1 U19326 ( .IN2(n15804), .IN1(n15802), .Q(n15807) );
  OR2X1 U19327 ( .IN2(n15809), .IN1(n15808), .Q(n15813) );
  OR2X1 U19328 ( .IN2(n15811), .IN1(n15810), .Q(n15815) );
  OR2X1 U19329 ( .IN2(n15814), .IN1(n15812), .Q(n15825) );
  OR2X1 U19330 ( .IN2(n15817), .IN1(n15816), .Q(n15821) );
  OR2X1 U19331 ( .IN2(n15819), .IN1(n15818), .Q(n15823) );
  OR2X1 U19332 ( .IN2(n15822), .IN1(n15820), .Q(n15827) );
  OR2X1 U19333 ( .IN2(n15826), .IN1(n15824), .Q(n15842) );
  OR2X1 U19334 ( .IN2(n15829), .IN1(n15828), .Q(n15833) );
  OR2X1 U19335 ( .IN2(n15831), .IN1(n15830), .Q(n15835) );
  OR2X1 U19336 ( .IN2(n15834), .IN1(n15832), .Q(n15839) );
  OR2X1 U19337 ( .IN2(n15837), .IN1(n15836), .Q(n15841) );
  OR2X1 U19338 ( .IN2(n15840), .IN1(n15838), .Q(n15843) );
  OR2X1 U19339 ( .IN2(n15845), .IN1(n15844), .Q(n15849) );
  OR2X1 U19340 ( .IN2(n15847), .IN1(n15846), .Q(n15851) );
  OR2X1 U19341 ( .IN2(n15850), .IN1(n15848), .Q(n15861) );
  OR2X1 U19342 ( .IN2(n15853), .IN1(n15852), .Q(n15857) );
  OR2X1 U19343 ( .IN2(n15855), .IN1(n15854), .Q(n15859) );
  OR2X1 U19344 ( .IN2(n15858), .IN1(n15856), .Q(n15863) );
  OR2X1 U19345 ( .IN2(n15862), .IN1(n15860), .Q(n15875) );
  OR2X1 U19346 ( .IN2(n15865), .IN1(n15864), .Q(n15869) );
  OR2X1 U19347 ( .IN2(n15867), .IN1(n15866), .Q(n15871) );
  OR2X1 U19348 ( .IN2(n15870), .IN1(n15868), .Q(n15874) );
  OR2X1 U19349 ( .IN2(n15873), .IN1(n15872), .Q(n15876) );
  OR2X1 U19350 ( .IN2(n15878), .IN1(n15877), .Q(n15882) );
  OR2X1 U19351 ( .IN2(n15880), .IN1(n15879), .Q(n15884) );
  OR2X1 U19352 ( .IN2(n15883), .IN1(n15881), .Q(n15894) );
  OR2X1 U19353 ( .IN2(n15886), .IN1(n15885), .Q(n15890) );
  OR2X1 U19354 ( .IN2(n15888), .IN1(n15887), .Q(n15892) );
  OR2X1 U19355 ( .IN2(n15891), .IN1(n15889), .Q(n15896) );
  OR2X1 U19356 ( .IN2(n15895), .IN1(n15893), .Q(n15908) );
  OR2X1 U19357 ( .IN2(n15898), .IN1(n15897), .Q(n15902) );
  OR2X1 U19358 ( .IN2(n15900), .IN1(n15899), .Q(n15904) );
  OR2X1 U19359 ( .IN2(n15903), .IN1(n15901), .Q(n15907) );
  OR2X1 U19360 ( .IN2(n15906), .IN1(n15905), .Q(n15909) );
  OR2X1 U19361 ( .IN2(n15911), .IN1(n15910), .Q(n15915) );
  OR2X1 U19362 ( .IN2(n15913), .IN1(n15912), .Q(n15917) );
  OR2X1 U19363 ( .IN2(n15916), .IN1(n15914), .Q(n15927) );
  OR2X1 U19364 ( .IN2(n15919), .IN1(n15918), .Q(n15923) );
  OR2X1 U19365 ( .IN2(n15921), .IN1(n15920), .Q(n15925) );
  OR2X1 U19366 ( .IN2(n15924), .IN1(n15922), .Q(n15929) );
  OR2X1 U19367 ( .IN2(n15928), .IN1(n15926), .Q(n15941) );
  OR2X1 U19368 ( .IN2(n15931), .IN1(n15930), .Q(n15935) );
  OR2X1 U19369 ( .IN2(n15933), .IN1(n15932), .Q(n15937) );
  OR2X1 U19370 ( .IN2(n15936), .IN1(n15934), .Q(n15940) );
  OR2X1 U19371 ( .IN2(n15939), .IN1(n15938), .Q(n15942) );
  OR2X1 U19372 ( .IN2(n15944), .IN1(n15943), .Q(n15948) );
  OR2X1 U19373 ( .IN2(n15946), .IN1(n15945), .Q(n15950) );
  OR2X1 U19188 ( .IN2(n15390), .IN1(n15388), .Q(n15395) );
  OR2X1 U19189 ( .IN2(n15394), .IN1(n15392), .Q(n15410) );
  OR2X1 U19190 ( .IN2(n15397), .IN1(n15396), .Q(n15401) );
  OR2X1 U19191 ( .IN2(n15399), .IN1(n15398), .Q(n15403) );
  OR2X1 U19192 ( .IN2(n15402), .IN1(n15400), .Q(n15407) );
  OR2X1 U19193 ( .IN2(n15405), .IN1(n15404), .Q(n15409) );
  OR2X1 U19194 ( .IN2(n15408), .IN1(n15406), .Q(n15411) );
  OR2X1 U19195 ( .IN2(n15413), .IN1(n15412), .Q(n15417) );
  OR2X1 U19196 ( .IN2(n15415), .IN1(n15414), .Q(n15419) );
  OR2X1 U19197 ( .IN2(n15418), .IN1(n15416), .Q(n15429) );
  OR2X1 U19198 ( .IN2(n15421), .IN1(n15420), .Q(n15425) );
  OR2X1 U19199 ( .IN2(n15423), .IN1(n15422), .Q(n15427) );
  OR2X1 U19200 ( .IN2(n15426), .IN1(n15424), .Q(n15431) );
  OR2X1 U19201 ( .IN2(n15430), .IN1(n15428), .Q(n15446) );
  OR2X1 U19202 ( .IN2(n15433), .IN1(n15432), .Q(n15437) );
  OR2X1 U19203 ( .IN2(n15435), .IN1(n15434), .Q(n15439) );
  OR2X1 U19204 ( .IN2(n15438), .IN1(n15436), .Q(n15443) );
  OR2X1 U19205 ( .IN2(n15441), .IN1(n15440), .Q(n15445) );
  OR2X1 U19206 ( .IN2(n15444), .IN1(n15442), .Q(n15447) );
  OR2X1 U19207 ( .IN2(n15449), .IN1(n15448), .Q(n15453) );
  OR2X1 U19208 ( .IN2(n15451), .IN1(n15450), .Q(n15455) );
  OR2X1 U19209 ( .IN2(n15454), .IN1(n15452), .Q(n15465) );
  OR2X1 U19210 ( .IN2(n15457), .IN1(n15456), .Q(n15461) );
  OR2X1 U19211 ( .IN2(n15459), .IN1(n15458), .Q(n15463) );
  OR2X1 U19212 ( .IN2(n15462), .IN1(n15460), .Q(n15467) );
  OR2X1 U19213 ( .IN2(n15466), .IN1(n15464), .Q(n15482) );
  OR2X1 U19214 ( .IN2(n15469), .IN1(n15468), .Q(n15473) );
  OR2X1 U19215 ( .IN2(n15471), .IN1(n15470), .Q(n15475) );
  OR2X1 U19216 ( .IN2(n15474), .IN1(n15472), .Q(n15479) );
  OR2X1 U19217 ( .IN2(n15477), .IN1(n15476), .Q(n15481) );
  OR2X1 U19218 ( .IN2(n15480), .IN1(n15478), .Q(n15483) );
  OR2X1 U19219 ( .IN2(n15485), .IN1(n15484), .Q(n15489) );
  OR2X1 U19220 ( .IN2(n15487), .IN1(n15486), .Q(n15491) );
  OR2X1 U19221 ( .IN2(n15490), .IN1(n15488), .Q(n15501) );
  OR2X1 U19222 ( .IN2(n15493), .IN1(n15492), .Q(n15497) );
  OR2X1 U19223 ( .IN2(n15495), .IN1(n15494), .Q(n15499) );
  OR2X1 U19224 ( .IN2(n15498), .IN1(n15496), .Q(n15503) );
  OR2X1 U19225 ( .IN2(n15502), .IN1(n15500), .Q(n15518) );
  OR2X1 U19226 ( .IN2(n15505), .IN1(n15504), .Q(n15509) );
  OR2X1 U19227 ( .IN2(n15507), .IN1(n15506), .Q(n15511) );
  OR2X1 U19228 ( .IN2(n15510), .IN1(n15508), .Q(n15515) );
  OR2X1 U19229 ( .IN2(n15513), .IN1(n15512), .Q(n15517) );
  OR2X1 U19230 ( .IN2(n15516), .IN1(n15514), .Q(n15519) );
  OR2X1 U19231 ( .IN2(n15521), .IN1(n15520), .Q(n15525) );
  OR2X1 U19232 ( .IN2(n15523), .IN1(n15522), .Q(n15527) );
  OR2X1 U19233 ( .IN2(n15526), .IN1(n15524), .Q(n15537) );
  OR2X1 U19234 ( .IN2(n15529), .IN1(n15528), .Q(n15533) );
  OR2X1 U19235 ( .IN2(n15531), .IN1(n15530), .Q(n15535) );
  OR2X1 U19236 ( .IN2(n15534), .IN1(n15532), .Q(n15539) );
  OR2X1 U19237 ( .IN2(n15538), .IN1(n15536), .Q(n15554) );
  OR2X1 U19238 ( .IN2(n15541), .IN1(n15540), .Q(n15545) );
  OR2X1 U19239 ( .IN2(n15543), .IN1(n15542), .Q(n15547) );
  OR2X1 U19240 ( .IN2(n15546), .IN1(n15544), .Q(n15551) );
  OR2X1 U19241 ( .IN2(n15549), .IN1(n15548), .Q(n15553) );
  OR2X1 U19242 ( .IN2(n15552), .IN1(n15550), .Q(n15555) );
  OR2X1 U19243 ( .IN2(n15557), .IN1(n15556), .Q(n15561) );
  OR2X1 U19244 ( .IN2(n15559), .IN1(n15558), .Q(n15563) );
  OR2X1 U19245 ( .IN2(n15562), .IN1(n15560), .Q(n15573) );
  OR2X1 U19246 ( .IN2(n15565), .IN1(n15564), .Q(n15569) );
  OR2X1 U19247 ( .IN2(n15567), .IN1(n15566), .Q(n15571) );
  OR2X1 U19248 ( .IN2(n15570), .IN1(n15568), .Q(n15575) );
  OR2X1 U19249 ( .IN2(n15574), .IN1(n15572), .Q(n15590) );
  OR2X1 U19250 ( .IN2(n15577), .IN1(n15576), .Q(n15581) );
  OR2X1 U19251 ( .IN2(n15579), .IN1(n15578), .Q(n15583) );
  OR2X1 U19252 ( .IN2(n15582), .IN1(n15580), .Q(n15587) );
  OR2X1 U19253 ( .IN2(n15585), .IN1(n15584), .Q(n15589) );
  OR2X1 U19254 ( .IN2(n15588), .IN1(n15586), .Q(n15591) );
  OR2X1 U19255 ( .IN2(n15593), .IN1(n15592), .Q(n15597) );
  OR2X1 U19256 ( .IN2(n15595), .IN1(n15594), .Q(n15599) );
  OR2X1 U19257 ( .IN2(n15598), .IN1(n15596), .Q(n15609) );
  OR2X1 U19258 ( .IN2(n15601), .IN1(n15600), .Q(n15605) );
  OR2X1 U19259 ( .IN2(n15603), .IN1(n15602), .Q(n15607) );
  OR2X1 U19260 ( .IN2(n15606), .IN1(n15604), .Q(n15611) );
  OR2X1 U19261 ( .IN2(n15610), .IN1(n15608), .Q(n15626) );
  OR2X1 U19262 ( .IN2(n15613), .IN1(n15612), .Q(n15617) );
  OR2X1 U19263 ( .IN2(n15615), .IN1(n15614), .Q(n15619) );
  OR2X1 U19264 ( .IN2(n15618), .IN1(n15616), .Q(n15623) );
  OR2X1 U19265 ( .IN2(n15621), .IN1(n15620), .Q(n15625) );
  OR2X1 U19266 ( .IN2(n15624), .IN1(n15622), .Q(n15627) );
  OR2X1 U19267 ( .IN2(n15629), .IN1(n15628), .Q(n15633) );
  OR2X1 U19268 ( .IN2(n15631), .IN1(n15630), .Q(n15635) );
  OR2X1 U19269 ( .IN2(n15634), .IN1(n15632), .Q(n15645) );
  OR2X1 U19270 ( .IN2(n15637), .IN1(n15636), .Q(n15641) );
  OR2X1 U19271 ( .IN2(n15639), .IN1(n15638), .Q(n15643) );
  OR2X1 U19272 ( .IN2(n15642), .IN1(n15640), .Q(n15647) );
  OR2X1 U19273 ( .IN2(n15646), .IN1(n15644), .Q(n15662) );
  OR2X1 U19274 ( .IN2(n15649), .IN1(n15648), .Q(n15653) );
  OR2X1 U19275 ( .IN2(n15651), .IN1(n15650), .Q(n15655) );
  OR2X1 U19276 ( .IN2(n15654), .IN1(n15652), .Q(n15659) );
  OR2X1 U19277 ( .IN2(n15657), .IN1(n15656), .Q(n15661) );
  OR2X1 U19278 ( .IN2(n15660), .IN1(n15658), .Q(n15663) );
  OR2X1 U19279 ( .IN2(n15665), .IN1(n15664), .Q(n15669) );
  OR2X1 U19280 ( .IN2(n15667), .IN1(n15666), .Q(n15671) );
  OR2X1 U19095 ( .IN2(n15111), .IN1(n15110), .Q(n15115) );
  OR2X1 U19096 ( .IN2(n15114), .IN1(n15112), .Q(n15119) );
  OR2X1 U19097 ( .IN2(n15117), .IN1(n15116), .Q(n15121) );
  OR2X1 U19098 ( .IN2(n15120), .IN1(n15118), .Q(n15123) );
  OR2X1 U19099 ( .IN2(n15125), .IN1(n15124), .Q(n15129) );
  OR2X1 U19100 ( .IN2(n15127), .IN1(n15126), .Q(n15131) );
  OR2X1 U19101 ( .IN2(n15130), .IN1(n15128), .Q(n15141) );
  OR2X1 U19102 ( .IN2(n15133), .IN1(n15132), .Q(n15137) );
  OR2X1 U19103 ( .IN2(n15135), .IN1(n15134), .Q(n15139) );
  OR2X1 U19104 ( .IN2(n15138), .IN1(n15136), .Q(n15143) );
  OR2X1 U19105 ( .IN2(n15142), .IN1(n15140), .Q(n15158) );
  OR2X1 U19106 ( .IN2(n15145), .IN1(n15144), .Q(n15149) );
  OR2X1 U19107 ( .IN2(n15147), .IN1(n15146), .Q(n15151) );
  OR2X1 U19108 ( .IN2(n15150), .IN1(n15148), .Q(n15155) );
  OR2X1 U19109 ( .IN2(n15153), .IN1(n15152), .Q(n15157) );
  OR2X1 U19110 ( .IN2(n15156), .IN1(n15154), .Q(n15159) );
  OR2X1 U19111 ( .IN2(n15161), .IN1(n15160), .Q(n15165) );
  OR2X1 U19112 ( .IN2(n15163), .IN1(n15162), .Q(n15167) );
  OR2X1 U19113 ( .IN2(n15166), .IN1(n15164), .Q(n15177) );
  OR2X1 U19114 ( .IN2(n15169), .IN1(n15168), .Q(n15173) );
  OR2X1 U19115 ( .IN2(n15171), .IN1(n15170), .Q(n15175) );
  OR2X1 U19116 ( .IN2(n15174), .IN1(n15172), .Q(n15179) );
  OR2X1 U19117 ( .IN2(n15178), .IN1(n15176), .Q(n15194) );
  OR2X1 U19118 ( .IN2(n15181), .IN1(n15180), .Q(n15185) );
  OR2X1 U19119 ( .IN2(n15183), .IN1(n15182), .Q(n15187) );
  OR2X1 U19120 ( .IN2(n15186), .IN1(n15184), .Q(n15191) );
  OR2X1 U19121 ( .IN2(n15189), .IN1(n15188), .Q(n15193) );
  OR2X1 U19122 ( .IN2(n15192), .IN1(n15190), .Q(n15195) );
  OR2X1 U19123 ( .IN2(n15197), .IN1(n15196), .Q(n15201) );
  OR2X1 U19124 ( .IN2(n15199), .IN1(n15198), .Q(n15203) );
  OR2X1 U19125 ( .IN2(n15202), .IN1(n15200), .Q(n15213) );
  OR2X1 U19126 ( .IN2(n15205), .IN1(n15204), .Q(n15209) );
  OR2X1 U19127 ( .IN2(n15207), .IN1(n15206), .Q(n15211) );
  OR2X1 U19128 ( .IN2(n15210), .IN1(n15208), .Q(n15215) );
  OR2X1 U19129 ( .IN2(n15214), .IN1(n15212), .Q(n15230) );
  OR2X1 U19130 ( .IN2(n15217), .IN1(n15216), .Q(n15221) );
  OR2X1 U19131 ( .IN2(n15219), .IN1(n15218), .Q(n15223) );
  OR2X1 U19132 ( .IN2(n15222), .IN1(n15220), .Q(n15227) );
  OR2X1 U19133 ( .IN2(n15225), .IN1(n15224), .Q(n15229) );
  OR2X1 U19134 ( .IN2(n15228), .IN1(n15226), .Q(n15231) );
  OR2X1 U19135 ( .IN2(n15233), .IN1(n15232), .Q(n15237) );
  OR2X1 U19136 ( .IN2(n15235), .IN1(n15234), .Q(n15239) );
  OR2X1 U19137 ( .IN2(n15238), .IN1(n15236), .Q(n15249) );
  OR2X1 U19138 ( .IN2(n15241), .IN1(n15240), .Q(n15245) );
  OR2X1 U19139 ( .IN2(n15243), .IN1(n15242), .Q(n15247) );
  OR2X1 U19140 ( .IN2(n15246), .IN1(n15244), .Q(n15251) );
  OR2X1 U19141 ( .IN2(n15250), .IN1(n15248), .Q(n15266) );
  OR2X1 U19142 ( .IN2(n15253), .IN1(n15252), .Q(n15257) );
  OR2X1 U19143 ( .IN2(n15255), .IN1(n15254), .Q(n15259) );
  OR2X1 U19144 ( .IN2(n15258), .IN1(n15256), .Q(n15263) );
  OR2X1 U19145 ( .IN2(n15261), .IN1(n15260), .Q(n15265) );
  OR2X1 U19146 ( .IN2(n15264), .IN1(n15262), .Q(n15267) );
  OR2X1 U19147 ( .IN2(n15269), .IN1(n15268), .Q(n15273) );
  OR2X1 U19148 ( .IN2(n15271), .IN1(n15270), .Q(n15275) );
  OR2X1 U19149 ( .IN2(n15274), .IN1(n15272), .Q(n15285) );
  OR2X1 U19150 ( .IN2(n15277), .IN1(n15276), .Q(n15281) );
  OR2X1 U19151 ( .IN2(n15279), .IN1(n15278), .Q(n15283) );
  OR2X1 U19152 ( .IN2(n15282), .IN1(n15280), .Q(n15287) );
  OR2X1 U19153 ( .IN2(n15286), .IN1(n15284), .Q(n15302) );
  OR2X1 U19154 ( .IN2(n15289), .IN1(n15288), .Q(n15293) );
  OR2X1 U19155 ( .IN2(n15291), .IN1(n15290), .Q(n15295) );
  OR2X1 U19156 ( .IN2(n15294), .IN1(n15292), .Q(n15299) );
  OR2X1 U19157 ( .IN2(n15297), .IN1(n15296), .Q(n15301) );
  OR2X1 U19158 ( .IN2(n15300), .IN1(n15298), .Q(n15303) );
  OR2X1 U19159 ( .IN2(n15305), .IN1(n15304), .Q(n15309) );
  OR2X1 U19160 ( .IN2(n15307), .IN1(n15306), .Q(n15311) );
  OR2X1 U19161 ( .IN2(n15310), .IN1(n15308), .Q(n15321) );
  OR2X1 U19162 ( .IN2(n15313), .IN1(n15312), .Q(n15317) );
  OR2X1 U19163 ( .IN2(n15315), .IN1(n15314), .Q(n15319) );
  OR2X1 U19164 ( .IN2(n15318), .IN1(n15316), .Q(n15323) );
  OR2X1 U19165 ( .IN2(n15322), .IN1(n15320), .Q(n15338) );
  OR2X1 U19166 ( .IN2(n15325), .IN1(n15324), .Q(n15329) );
  OR2X1 U19167 ( .IN2(n15327), .IN1(n15326), .Q(n15331) );
  OR2X1 U19168 ( .IN2(n15330), .IN1(n15328), .Q(n15335) );
  OR2X1 U19169 ( .IN2(n15333), .IN1(n15332), .Q(n15337) );
  OR2X1 U19170 ( .IN2(n15336), .IN1(n15334), .Q(n15339) );
  OR2X1 U19171 ( .IN2(n15341), .IN1(n15340), .Q(n15345) );
  OR2X1 U19172 ( .IN2(n15343), .IN1(n15342), .Q(n15347) );
  OR2X1 U19173 ( .IN2(n15346), .IN1(n15344), .Q(n15357) );
  OR2X1 U19174 ( .IN2(n15349), .IN1(n15348), .Q(n15353) );
  OR2X1 U19175 ( .IN2(n15351), .IN1(n15350), .Q(n15355) );
  OR2X1 U19176 ( .IN2(n15354), .IN1(n15352), .Q(n15359) );
  OR2X1 U19177 ( .IN2(n15358), .IN1(n15356), .Q(n15374) );
  OR2X1 U19178 ( .IN2(n15361), .IN1(n15360), .Q(n15365) );
  OR2X1 U19179 ( .IN2(n15363), .IN1(n15362), .Q(n15367) );
  OR2X1 U19180 ( .IN2(n15366), .IN1(n15364), .Q(n15371) );
  OR2X1 U19181 ( .IN2(n15369), .IN1(n15368), .Q(n15373) );
  OR2X1 U19182 ( .IN2(n15372), .IN1(n15370), .Q(n15375) );
  OR2X1 U19183 ( .IN2(n15377), .IN1(n15376), .Q(n15381) );
  OR2X1 U19184 ( .IN2(n15379), .IN1(n15378), .Q(n15383) );
  OR2X1 U19185 ( .IN2(n15382), .IN1(n15380), .Q(n15393) );
  OR2X1 U19186 ( .IN2(n15385), .IN1(n15384), .Q(n15389) );
  OR2X1 U19187 ( .IN2(n15387), .IN1(n15386), .Q(n15391) );
  OR2X1 U19002 ( .IN2(n14832), .IN1(n14830), .Q(n14835) );
  OR2X1 U19003 ( .IN2(n14837), .IN1(n14836), .Q(n14841) );
  OR2X1 U19004 ( .IN2(n14839), .IN1(n14838), .Q(n14843) );
  OR2X1 U19005 ( .IN2(n14842), .IN1(n14840), .Q(n14853) );
  OR2X1 U19006 ( .IN2(n14845), .IN1(n14844), .Q(n14849) );
  OR2X1 U19007 ( .IN2(n14847), .IN1(n14846), .Q(n14851) );
  OR2X1 U19008 ( .IN2(n14850), .IN1(n14848), .Q(n14855) );
  OR2X1 U19009 ( .IN2(n14854), .IN1(n14852), .Q(n14870) );
  OR2X1 U19010 ( .IN2(n14857), .IN1(n14856), .Q(n14861) );
  OR2X1 U19011 ( .IN2(n14859), .IN1(n14858), .Q(n14863) );
  OR2X1 U19012 ( .IN2(n14862), .IN1(n14860), .Q(n14867) );
  OR2X1 U19013 ( .IN2(n14865), .IN1(n14864), .Q(n14869) );
  OR2X1 U19014 ( .IN2(n14868), .IN1(n14866), .Q(n14871) );
  OR2X1 U19015 ( .IN2(n14873), .IN1(n14872), .Q(n14877) );
  OR2X1 U19016 ( .IN2(n14875), .IN1(n14874), .Q(n14879) );
  OR2X1 U19017 ( .IN2(n14878), .IN1(n14876), .Q(n14889) );
  OR2X1 U19018 ( .IN2(n14881), .IN1(n14880), .Q(n14885) );
  OR2X1 U19019 ( .IN2(n14883), .IN1(n14882), .Q(n14887) );
  OR2X1 U19020 ( .IN2(n14886), .IN1(n14884), .Q(n14891) );
  OR2X1 U19021 ( .IN2(n14890), .IN1(n14888), .Q(n14906) );
  OR2X1 U19022 ( .IN2(n14893), .IN1(n14892), .Q(n14897) );
  OR2X1 U19023 ( .IN2(n14895), .IN1(n14894), .Q(n14899) );
  OR2X1 U19024 ( .IN2(n14898), .IN1(n14896), .Q(n14903) );
  OR2X1 U19025 ( .IN2(n14901), .IN1(n14900), .Q(n14905) );
  OR2X1 U19026 ( .IN2(n14904), .IN1(n14902), .Q(n14907) );
  OR2X1 U19027 ( .IN2(n14909), .IN1(n14908), .Q(n14913) );
  OR2X1 U19028 ( .IN2(n14911), .IN1(n14910), .Q(n14915) );
  OR2X1 U19029 ( .IN2(n14914), .IN1(n14912), .Q(n14925) );
  OR2X1 U19030 ( .IN2(n14917), .IN1(n14916), .Q(n14921) );
  OR2X1 U19031 ( .IN2(n14919), .IN1(n14918), .Q(n14923) );
  OR2X1 U19032 ( .IN2(n14922), .IN1(n14920), .Q(n14927) );
  OR2X1 U19033 ( .IN2(n14926), .IN1(n14924), .Q(n14942) );
  OR2X1 U19034 ( .IN2(n14929), .IN1(n14928), .Q(n14933) );
  OR2X1 U19035 ( .IN2(n14931), .IN1(n14930), .Q(n14935) );
  OR2X1 U19036 ( .IN2(n14934), .IN1(n14932), .Q(n14939) );
  OR2X1 U19037 ( .IN2(n14937), .IN1(n14936), .Q(n14941) );
  OR2X1 U19038 ( .IN2(n14940), .IN1(n14938), .Q(n14943) );
  OR2X1 U19039 ( .IN2(n14945), .IN1(n14944), .Q(n14949) );
  OR2X1 U19040 ( .IN2(n14947), .IN1(n14946), .Q(n14951) );
  OR2X1 U19041 ( .IN2(n14950), .IN1(n14948), .Q(n14961) );
  OR2X1 U19042 ( .IN2(n14953), .IN1(n14952), .Q(n14957) );
  OR2X1 U19043 ( .IN2(n14955), .IN1(n14954), .Q(n14959) );
  OR2X1 U19044 ( .IN2(n14958), .IN1(n14956), .Q(n14963) );
  OR2X1 U19045 ( .IN2(n14962), .IN1(n14960), .Q(n14978) );
  OR2X1 U19046 ( .IN2(n14965), .IN1(n14964), .Q(n14969) );
  OR2X1 U19047 ( .IN2(n14967), .IN1(n14966), .Q(n14971) );
  OR2X1 U19048 ( .IN2(n14970), .IN1(n14968), .Q(n14975) );
  OR2X1 U19049 ( .IN2(n14973), .IN1(n14972), .Q(n14977) );
  OR2X1 U19050 ( .IN2(n14976), .IN1(n14974), .Q(n14979) );
  OR2X1 U19051 ( .IN2(n14981), .IN1(n14980), .Q(n14985) );
  OR2X1 U19052 ( .IN2(n14983), .IN1(n14982), .Q(n14987) );
  OR2X1 U19053 ( .IN2(n14986), .IN1(n14984), .Q(n14997) );
  OR2X1 U19054 ( .IN2(n14989), .IN1(n14988), .Q(n14993) );
  OR2X1 U19055 ( .IN2(n14991), .IN1(n14990), .Q(n14995) );
  OR2X1 U19056 ( .IN2(n14994), .IN1(n14992), .Q(n14999) );
  OR2X1 U19057 ( .IN2(n14998), .IN1(n14996), .Q(n15014) );
  OR2X1 U19058 ( .IN2(n15001), .IN1(n15000), .Q(n15005) );
  OR2X1 U19059 ( .IN2(n15003), .IN1(n15002), .Q(n15007) );
  OR2X1 U19060 ( .IN2(n15006), .IN1(n15004), .Q(n15011) );
  OR2X1 U19061 ( .IN2(n15009), .IN1(n15008), .Q(n15013) );
  OR2X1 U19062 ( .IN2(n15012), .IN1(n15010), .Q(n15015) );
  OR2X1 U19063 ( .IN2(n15017), .IN1(n15016), .Q(n15021) );
  OR2X1 U19064 ( .IN2(n15019), .IN1(n15018), .Q(n15023) );
  OR2X1 U19065 ( .IN2(n15022), .IN1(n15020), .Q(n15033) );
  OR2X1 U19066 ( .IN2(n15025), .IN1(n15024), .Q(n15029) );
  OR2X1 U19067 ( .IN2(n15027), .IN1(n15026), .Q(n15031) );
  OR2X1 U19068 ( .IN2(n15030), .IN1(n15028), .Q(n15035) );
  OR2X1 U19069 ( .IN2(n15034), .IN1(n15032), .Q(n15050) );
  OR2X1 U19070 ( .IN2(n15037), .IN1(n15036), .Q(n15041) );
  OR2X1 U19071 ( .IN2(n15039), .IN1(n15038), .Q(n15043) );
  OR2X1 U19072 ( .IN2(n15042), .IN1(n15040), .Q(n15047) );
  OR2X1 U19073 ( .IN2(n15045), .IN1(n15044), .Q(n15049) );
  OR2X1 U19074 ( .IN2(n15048), .IN1(n15046), .Q(n15051) );
  OR2X1 U19075 ( .IN2(n15053), .IN1(n15052), .Q(n15057) );
  OR2X1 U19076 ( .IN2(n15055), .IN1(n15054), .Q(n15059) );
  OR2X1 U19077 ( .IN2(n15058), .IN1(n15056), .Q(n15069) );
  OR2X1 U19078 ( .IN2(n15061), .IN1(n15060), .Q(n15065) );
  OR2X1 U19079 ( .IN2(n15063), .IN1(n15062), .Q(n15067) );
  OR2X1 U19080 ( .IN2(n15066), .IN1(n15064), .Q(n15071) );
  OR2X1 U19081 ( .IN2(n15070), .IN1(n15068), .Q(n15086) );
  OR2X1 U19082 ( .IN2(n15073), .IN1(n15072), .Q(n15077) );
  OR2X1 U19083 ( .IN2(n15075), .IN1(n15074), .Q(n15079) );
  OR2X1 U19084 ( .IN2(n15078), .IN1(n15076), .Q(n15083) );
  OR2X1 U19085 ( .IN2(n15081), .IN1(n15080), .Q(n15085) );
  OR2X1 U19086 ( .IN2(n15084), .IN1(n15082), .Q(n15087) );
  OR2X1 U19087 ( .IN2(n15089), .IN1(n15088), .Q(n15093) );
  OR2X1 U19088 ( .IN2(n15091), .IN1(n15090), .Q(n15095) );
  OR2X1 U19089 ( .IN2(n15094), .IN1(n15092), .Q(n15105) );
  OR2X1 U19090 ( .IN2(n15097), .IN1(n15096), .Q(n15101) );
  OR2X1 U19091 ( .IN2(n15099), .IN1(n15098), .Q(n15103) );
  OR2X1 U19092 ( .IN2(n15102), .IN1(n15100), .Q(n15107) );
  OR2X1 U19093 ( .IN2(n15106), .IN1(n15104), .Q(n15122) );
  OR2X1 U19094 ( .IN2(n15109), .IN1(n15108), .Q(n15113) );
  AND2X1 U18909 ( .IN1(n17640), .IN2(n6804), .Q(n17639) );
  AND2X1 U18910 ( .IN1(n17642), .IN2(n6803), .Q(n17641) );
  AND2X1 U18911 ( .IN1(n17643), .IN2(n6974), .Q(n14752) );
  AND2X1 U18912 ( .IN1(n17644), .IN2(n6967), .Q(n14753) );
  AND2X1 U18913 ( .IN1(P2_N933), .IN2(n6808), .Q(n17645) );
  AND2X1 U18914 ( .IN1(P2_N933), .IN2(n6807), .Q(n17646) );
  AND2X1 U18915 ( .IN1(P2_N933), .IN2(n6808), .Q(n17647) );
  AND2X1 U18916 ( .IN1(P2_N933), .IN2(n6807), .Q(n17648) );
  AND2X1 U18917 ( .IN1(n17650), .IN2(n6804), .Q(n17649) );
  AND2X1 U18918 ( .IN1(n17652), .IN2(n6803), .Q(n17651) );
  AND2X1 U18919 ( .IN1(P2_N933), .IN2(n6848), .Q(n17653) );
  AND2X1 U18920 ( .IN1(P2_N933), .IN2(n6847), .Q(n17654) );
  AND2X1 U18921 ( .IN1(P2_N933), .IN2(n6808), .Q(n17655) );
  AND2X1 U18922 ( .IN1(P2_N933), .IN2(n6847), .Q(n17656) );
  AND2X1 U18923 ( .IN1(n17658), .IN2(n6804), .Q(n17657) );
  AND2X1 U18924 ( .IN1(n17660), .IN2(n6803), .Q(n17659) );
  AND2X1 U18925 ( .IN1(n17662), .IN2(n6932), .Q(n17661) );
  AND2X1 U18926 ( .IN1(n17664), .IN2(n6931), .Q(n17663) );
  AND2X1 U18927 ( .IN1(P2_N933), .IN2(n6848), .Q(n17665) );
  AND2X1 U18928 ( .IN1(P2_N933), .IN2(n6847), .Q(n17666) );
  AND2X1 U18929 ( .IN1(P2_N933), .IN2(n6848), .Q(n17667) );
  AND2X1 U18930 ( .IN1(P2_N933), .IN2(n6847), .Q(n17668) );
  AND2X1 U18931 ( .IN1(n17670), .IN2(n6804), .Q(n17669) );
  AND2X1 U18932 ( .IN1(n17672), .IN2(n6803), .Q(n17671) );
  AND2X1 U18933 ( .IN1(n17673), .IN2(n6974), .Q(n14754) );
  AND2X1 U18934 ( .IN1(n17674), .IN2(n6967), .Q(n14755) );
  AND2X1 U18935 ( .IN1(P2_N934), .IN2(n6808), .Q(n17675) );
  AND2X1 U18936 ( .IN1(P2_N934), .IN2(n6807), .Q(n17676) );
  AND2X1 U18937 ( .IN1(P2_N934), .IN2(n6808), .Q(n17677) );
  AND2X1 U18938 ( .IN1(P2_N934), .IN2(n6807), .Q(n17678) );
  AND2X1 U18939 ( .IN1(n17680), .IN2(n6804), .Q(n17679) );
  AND2X1 U18940 ( .IN1(n17682), .IN2(n6803), .Q(n17681) );
  AND2X1 U18941 ( .IN1(P2_N934), .IN2(n6848), .Q(n17683) );
  AND2X1 U18942 ( .IN1(P2_N934), .IN2(n6847), .Q(n17684) );
  AND2X1 U18943 ( .IN1(P2_N934), .IN2(n6808), .Q(n17685) );
  AND2X1 U18944 ( .IN1(P2_N934), .IN2(n6807), .Q(n17686) );
  AND2X1 U18945 ( .IN1(n17688), .IN2(n6780), .Q(n17687) );
  AND2X1 U18946 ( .IN1(n17690), .IN2(P2_N291), .Q(n17689) );
  AND2X1 U18947 ( .IN1(n17692), .IN2(n6932), .Q(n17691) );
  AND2X1 U18948 ( .IN1(n17694), .IN2(n6931), .Q(n17693) );
  AND2X1 U18949 ( .IN1(P2_N934), .IN2(n6848), .Q(n17695) );
  AND2X1 U18950 ( .IN1(P2_N934), .IN2(n6847), .Q(n17696) );
  AND2X1 U18951 ( .IN1(P2_N934), .IN2(n6848), .Q(n17697) );
  AND2X1 U18952 ( .IN1(P2_N934), .IN2(n6847), .Q(n17698) );
  AND2X1 U18953 ( .IN1(n17700), .IN2(n6780), .Q(n17699) );
  AND2X1 U18954 ( .IN1(n17702), .IN2(P2_N291), .Q(n17701) );
  AND2X1 U18955 ( .IN1(n17703), .IN2(n6970), .Q(n14756) );
  AND2X1 U18956 ( .IN1(n17704), .IN2(n6967), .Q(n14757) );
  AND2X1 U18957 ( .IN1(n7012), .IN2(n6838), .Q(n17705) );
  AND2X1 U18958 ( .IN1(n7012), .IN2(n6837), .Q(n17706) );
  AND2X1 U18959 ( .IN1(n7012), .IN2(n6838), .Q(n17707) );
  AND2X1 U18960 ( .IN1(n7012), .IN2(n6837), .Q(n17708) );
  AND2X1 U18961 ( .IN1(n17710), .IN2(n6784), .Q(n17709) );
  AND2X1 U18962 ( .IN1(n17712), .IN2(n6793), .Q(n17711) );
  AND2X1 U18963 ( .IN1(n7012), .IN2(n6838), .Q(n17713) );
  AND2X1 U18964 ( .IN1(n7012), .IN2(n6837), .Q(n17714) );
  AND2X1 U18965 ( .IN1(n7012), .IN2(n6838), .Q(n17715) );
  AND2X1 U18966 ( .IN1(n7012), .IN2(n6837), .Q(n17716) );
  AND2X1 U18967 ( .IN1(n17718), .IN2(n6784), .Q(n17717) );
  AND2X1 U18968 ( .IN1(n17720), .IN2(n6793), .Q(n17719) );
  AND2X1 U18969 ( .IN1(n17722), .IN2(n6940), .Q(n17721) );
  AND2X1 U18970 ( .IN1(n17724), .IN2(n6943), .Q(n17723) );
  AND2X1 U18971 ( .IN1(n17726), .IN2(n17727), .Q(n17725) );
  AND2X1 U18972 ( .IN1(n17729), .IN2(n17730), .Q(n17728) );
  AND2X1 U18973 ( .IN1(n17731), .IN2(n17732), .Q(n14759) );
  AND2X1 U18974 ( .IN1(n17733), .IN2(n6972), .Q(n14760) );
  AND2X1 U18975 ( .IN1(n14758), .IN2(n6969), .Q(n14761) );
  OR2X1 U18977 ( .IN2(n6838), .IN1(P2_N1413), .Q(n17019) );
  OR2X1 U18979 ( .IN2(n14764), .IN1(n14762), .Q(n14774) );
  OR2X1 U18980 ( .IN2(n14766), .IN1(n14765), .Q(n14770) );
  OR2X1 U18981 ( .IN2(n14768), .IN1(n14767), .Q(n14772) );
  OR2X1 U18982 ( .IN2(n14771), .IN1(n14769), .Q(n14776) );
  OR2X1 U18983 ( .IN2(n14775), .IN1(n14773), .Q(n14798) );
  OR2X1 U18984 ( .IN2(n14778), .IN1(n14777), .Q(n14782) );
  OR2X1 U18985 ( .IN2(n14780), .IN1(n14779), .Q(n14784) );
  OR2X1 U18986 ( .IN2(n14783), .IN1(n14781), .Q(n14794) );
  OR2X1 U18987 ( .IN2(n14786), .IN1(n14785), .Q(n14790) );
  OR2X1 U18988 ( .IN2(n14788), .IN1(n14787), .Q(n14792) );
  OR2X1 U18989 ( .IN2(n14791), .IN1(n14789), .Q(n14796) );
  OR2X1 U18990 ( .IN2(n14795), .IN1(n14793), .Q(n14799) );
  OR2X1 U18991 ( .IN2(n14801), .IN1(n14800), .Q(n14805) );
  OR2X1 U18992 ( .IN2(n14803), .IN1(n14802), .Q(n14807) );
  OR2X1 U18993 ( .IN2(n14806), .IN1(n14804), .Q(n14817) );
  OR2X1 U18994 ( .IN2(n14809), .IN1(n14808), .Q(n14813) );
  OR2X1 U18995 ( .IN2(n14811), .IN1(n14810), .Q(n14815) );
  OR2X1 U18996 ( .IN2(n14814), .IN1(n14812), .Q(n14819) );
  OR2X1 U18997 ( .IN2(n14818), .IN1(n14816), .Q(n14834) );
  OR2X1 U18998 ( .IN2(n14821), .IN1(n14820), .Q(n14825) );
  OR2X1 U18999 ( .IN2(n14823), .IN1(n14822), .Q(n14827) );
  OR2X1 U19000 ( .IN2(n14826), .IN1(n14824), .Q(n14831) );
  OR2X1 U19001 ( .IN2(n14829), .IN1(n14828), .Q(n14833) );
  AND2X1 U18816 ( .IN1(n17514), .IN2(n6931), .Q(n17513) );
  AND2X1 U18817 ( .IN1(P2_N928), .IN2(n6832), .Q(n17515) );
  AND2X1 U18818 ( .IN1(P2_N928), .IN2(n6831), .Q(n17516) );
  AND2X1 U18819 ( .IN1(P2_N928), .IN2(n6832), .Q(n17517) );
  AND2X1 U18820 ( .IN1(P2_N928), .IN2(n6831), .Q(n17518) );
  AND2X1 U18821 ( .IN1(n17520), .IN2(n6804), .Q(n17519) );
  AND2X1 U18822 ( .IN1(n17522), .IN2(n6803), .Q(n17521) );
  AND2X1 U18823 ( .IN1(n17523), .IN2(n6974), .Q(n14744) );
  AND2X1 U18824 ( .IN1(n17524), .IN2(n6967), .Q(n14745) );
  AND2X1 U18825 ( .IN1(P2_N929), .IN2(n6808), .Q(n17525) );
  AND2X1 U18826 ( .IN1(P2_N929), .IN2(n6807), .Q(n17526) );
  AND2X1 U18827 ( .IN1(P2_N929), .IN2(n6808), .Q(n17527) );
  AND2X1 U18828 ( .IN1(P2_N929), .IN2(n6807), .Q(n17528) );
  AND2X1 U18829 ( .IN1(n17530), .IN2(n6804), .Q(n17529) );
  AND2X1 U18830 ( .IN1(n17532), .IN2(n6803), .Q(n17531) );
  AND2X1 U18831 ( .IN1(P2_N929), .IN2(n6810), .Q(n17533) );
  AND2X1 U18832 ( .IN1(P2_N929), .IN2(n6807), .Q(n17534) );
  AND2X1 U18833 ( .IN1(P2_N929), .IN2(n6810), .Q(n17535) );
  AND2X1 U18834 ( .IN1(P2_N929), .IN2(n6807), .Q(n17536) );
  AND2X1 U18835 ( .IN1(n17538), .IN2(n6804), .Q(n17537) );
  AND2X1 U18836 ( .IN1(n17540), .IN2(n6803), .Q(n17539) );
  AND2X1 U18837 ( .IN1(n17542), .IN2(n6932), .Q(n17541) );
  AND2X1 U18838 ( .IN1(n17544), .IN2(n6931), .Q(n17543) );
  AND2X1 U18839 ( .IN1(P2_N929), .IN2(n6832), .Q(n17545) );
  AND2X1 U18840 ( .IN1(P2_N929), .IN2(n6807), .Q(n17546) );
  AND2X1 U18841 ( .IN1(P2_N929), .IN2(n6832), .Q(n17547) );
  AND2X1 U18842 ( .IN1(P2_N929), .IN2(n6807), .Q(n17548) );
  AND2X1 U18843 ( .IN1(n17550), .IN2(n6804), .Q(n17549) );
  AND2X1 U18844 ( .IN1(n17552), .IN2(n6803), .Q(n17551) );
  AND2X1 U18845 ( .IN1(n17553), .IN2(n6974), .Q(n14746) );
  AND2X1 U18846 ( .IN1(n17554), .IN2(n6967), .Q(n14747) );
  AND2X1 U18847 ( .IN1(P2_N930), .IN2(n6808), .Q(n17555) );
  AND2X1 U18848 ( .IN1(P2_N930), .IN2(n6807), .Q(n17556) );
  AND2X1 U18849 ( .IN1(P2_N930), .IN2(n6808), .Q(n17557) );
  AND2X1 U18850 ( .IN1(P2_N930), .IN2(n6807), .Q(n17558) );
  AND2X1 U18851 ( .IN1(n17560), .IN2(n6804), .Q(n17559) );
  AND2X1 U18852 ( .IN1(n17562), .IN2(n6803), .Q(n17561) );
  AND2X1 U18853 ( .IN1(P2_N930), .IN2(n6810), .Q(n17563) );
  AND2X1 U18854 ( .IN1(P2_N930), .IN2(n6807), .Q(n17564) );
  AND2X1 U18855 ( .IN1(P2_N930), .IN2(n6808), .Q(n17565) );
  AND2X1 U18856 ( .IN1(P2_N930), .IN2(n6807), .Q(n17566) );
  AND2X1 U18857 ( .IN1(n17568), .IN2(n6804), .Q(n17567) );
  AND2X1 U18858 ( .IN1(n17570), .IN2(n6803), .Q(n17569) );
  AND2X1 U18859 ( .IN1(n17572), .IN2(n6932), .Q(n17571) );
  AND2X1 U18860 ( .IN1(n17574), .IN2(n6931), .Q(n17573) );
  AND2X1 U18861 ( .IN1(P2_N930), .IN2(n6832), .Q(n17575) );
  AND2X1 U18862 ( .IN1(P2_N930), .IN2(n6807), .Q(n17576) );
  AND2X1 U18863 ( .IN1(P2_N930), .IN2(n6832), .Q(n17577) );
  AND2X1 U18864 ( .IN1(P2_N930), .IN2(n6807), .Q(n17578) );
  AND2X1 U18865 ( .IN1(n17580), .IN2(n6804), .Q(n17579) );
  AND2X1 U18866 ( .IN1(n17582), .IN2(n6803), .Q(n17581) );
  AND2X1 U18867 ( .IN1(n17583), .IN2(n6974), .Q(n14748) );
  AND2X1 U18868 ( .IN1(n17584), .IN2(n6967), .Q(n14749) );
  AND2X1 U18869 ( .IN1(P2_N931), .IN2(n6808), .Q(n17585) );
  AND2X1 U18870 ( .IN1(P2_N931), .IN2(n6807), .Q(n17586) );
  AND2X1 U18871 ( .IN1(P2_N931), .IN2(n6808), .Q(n17587) );
  AND2X1 U18872 ( .IN1(P2_N931), .IN2(n6807), .Q(n17588) );
  AND2X1 U18873 ( .IN1(n17590), .IN2(n6804), .Q(n17589) );
  AND2X1 U18874 ( .IN1(n17592), .IN2(n6803), .Q(n17591) );
  AND2X1 U18875 ( .IN1(P2_N931), .IN2(n6808), .Q(n17593) );
  AND2X1 U18876 ( .IN1(P2_N931), .IN2(n6807), .Q(n17594) );
  AND2X1 U18877 ( .IN1(P2_N931), .IN2(n6808), .Q(n17595) );
  AND2X1 U18878 ( .IN1(P2_N931), .IN2(n6807), .Q(n17596) );
  AND2X1 U18879 ( .IN1(n17598), .IN2(n6804), .Q(n17597) );
  AND2X1 U18880 ( .IN1(n17600), .IN2(n6803), .Q(n17599) );
  AND2X1 U18881 ( .IN1(n17602), .IN2(n6932), .Q(n17601) );
  AND2X1 U18882 ( .IN1(n17604), .IN2(n6931), .Q(n17603) );
  AND2X1 U18883 ( .IN1(P2_N931), .IN2(n6808), .Q(n17605) );
  AND2X1 U18884 ( .IN1(P2_N931), .IN2(n6807), .Q(n17606) );
  AND2X1 U18885 ( .IN1(P2_N931), .IN2(n6808), .Q(n17607) );
  AND2X1 U18886 ( .IN1(P2_N931), .IN2(n6807), .Q(n17608) );
  AND2X1 U18887 ( .IN1(n17610), .IN2(n6804), .Q(n17609) );
  AND2X1 U18888 ( .IN1(n17612), .IN2(n6803), .Q(n17611) );
  AND2X1 U18889 ( .IN1(n17613), .IN2(n6974), .Q(n14750) );
  AND2X1 U18890 ( .IN1(n17614), .IN2(n6967), .Q(n14751) );
  AND2X1 U18891 ( .IN1(P2_N932), .IN2(n6808), .Q(n17615) );
  AND2X1 U18892 ( .IN1(P2_N932), .IN2(n6807), .Q(n17616) );
  AND2X1 U18893 ( .IN1(P2_N932), .IN2(n6808), .Q(n17617) );
  AND2X1 U18894 ( .IN1(P2_N932), .IN2(n6807), .Q(n17618) );
  AND2X1 U18895 ( .IN1(n17620), .IN2(n6804), .Q(n17619) );
  AND2X1 U18896 ( .IN1(n17622), .IN2(n6803), .Q(n17621) );
  AND2X1 U18897 ( .IN1(P2_N932), .IN2(n6808), .Q(n17623) );
  AND2X1 U18898 ( .IN1(P2_N932), .IN2(n6807), .Q(n17624) );
  AND2X1 U18899 ( .IN1(P2_N932), .IN2(n6808), .Q(n17625) );
  AND2X1 U18900 ( .IN1(P2_N932), .IN2(n6807), .Q(n17626) );
  AND2X1 U18901 ( .IN1(n17628), .IN2(n6804), .Q(n17627) );
  AND2X1 U18902 ( .IN1(n17630), .IN2(n6803), .Q(n17629) );
  AND2X1 U18903 ( .IN1(n17632), .IN2(n6932), .Q(n17631) );
  AND2X1 U18904 ( .IN1(n17634), .IN2(n6931), .Q(n17633) );
  AND2X1 U18905 ( .IN1(P2_N932), .IN2(n6808), .Q(n17635) );
  AND2X1 U18906 ( .IN1(P2_N932), .IN2(n6807), .Q(n17636) );
  AND2X1 U18907 ( .IN1(P2_N932), .IN2(n6808), .Q(n17637) );
  AND2X1 U18908 ( .IN1(P2_N932), .IN2(n6807), .Q(n17638) );
  AND2X1 U18723 ( .IN1(P2_N924), .IN2(n6832), .Q(n17385) );
  AND2X1 U18724 ( .IN1(P2_N924), .IN2(n6837), .Q(n17386) );
  AND2X1 U18725 ( .IN1(n17388), .IN2(n6780), .Q(n17387) );
  AND2X1 U18726 ( .IN1(n17390), .IN2(n6779), .Q(n17389) );
  AND2X1 U18727 ( .IN1(n17392), .IN2(n6932), .Q(n17391) );
  AND2X1 U18728 ( .IN1(n17394), .IN2(n6931), .Q(n17393) );
  AND2X1 U18729 ( .IN1(P2_N924), .IN2(n6832), .Q(n17395) );
  AND2X1 U18730 ( .IN1(P2_N924), .IN2(n6831), .Q(n17396) );
  AND2X1 U18731 ( .IN1(P2_N924), .IN2(n6832), .Q(n17397) );
  AND2X1 U18732 ( .IN1(P2_N924), .IN2(n6831), .Q(n17398) );
  AND2X1 U18733 ( .IN1(n17400), .IN2(n6780), .Q(n17399) );
  AND2X1 U18734 ( .IN1(n17402), .IN2(n6779), .Q(n17401) );
  AND2X1 U18735 ( .IN1(n17403), .IN2(n6972), .Q(n14736) );
  AND2X1 U18736 ( .IN1(n17404), .IN2(n6963), .Q(n14737) );
  AND2X1 U18737 ( .IN1(P2_N925), .IN2(n6848), .Q(n17405) );
  AND2X1 U18738 ( .IN1(P2_N925), .IN2(n6847), .Q(n17406) );
  AND2X1 U18739 ( .IN1(P2_N925), .IN2(n6848), .Q(n17407) );
  AND2X1 U18740 ( .IN1(P2_N925), .IN2(n6847), .Q(n17408) );
  AND2X1 U18741 ( .IN1(n17410), .IN2(n6780), .Q(n17409) );
  AND2X1 U18742 ( .IN1(n17412), .IN2(n6803), .Q(n17411) );
  AND2X1 U18743 ( .IN1(P2_N925), .IN2(n6810), .Q(n17413) );
  AND2X1 U18744 ( .IN1(P2_N925), .IN2(n6809), .Q(n17414) );
  AND2X1 U18745 ( .IN1(P2_N925), .IN2(n6810), .Q(n17415) );
  AND2X1 U18746 ( .IN1(P2_N925), .IN2(n6809), .Q(n17416) );
  AND2X1 U18747 ( .IN1(n17418), .IN2(n6780), .Q(n17417) );
  AND2X1 U18748 ( .IN1(n17420), .IN2(n6779), .Q(n17419) );
  AND2X1 U18749 ( .IN1(n17422), .IN2(n6932), .Q(n17421) );
  AND2X1 U18750 ( .IN1(n17424), .IN2(n6931), .Q(n17423) );
  AND2X1 U18751 ( .IN1(P2_N925), .IN2(n6832), .Q(n17425) );
  AND2X1 U18752 ( .IN1(P2_N925), .IN2(n6831), .Q(n17426) );
  AND2X1 U18753 ( .IN1(P2_N925), .IN2(n6832), .Q(n17427) );
  AND2X1 U18754 ( .IN1(P2_N925), .IN2(n6831), .Q(n17428) );
  AND2X1 U18755 ( .IN1(n17430), .IN2(n6804), .Q(n17429) );
  AND2X1 U18756 ( .IN1(n17432), .IN2(n6803), .Q(n17431) );
  AND2X1 U18757 ( .IN1(n17433), .IN2(n6974), .Q(n14738) );
  AND2X1 U18758 ( .IN1(n17434), .IN2(n6967), .Q(n14739) );
  AND2X1 U18759 ( .IN1(P2_N926), .IN2(n6810), .Q(n17435) );
  AND2X1 U18760 ( .IN1(P2_N926), .IN2(n6809), .Q(n17436) );
  AND2X1 U18761 ( .IN1(P2_N926), .IN2(n6810), .Q(n17437) );
  AND2X1 U18762 ( .IN1(P2_N926), .IN2(n6809), .Q(n17438) );
  AND2X1 U18763 ( .IN1(n17440), .IN2(n6780), .Q(n17439) );
  AND2X1 U18764 ( .IN1(n17442), .IN2(n6779), .Q(n17441) );
  AND2X1 U18765 ( .IN1(P2_N926), .IN2(n6810), .Q(n17443) );
  AND2X1 U18766 ( .IN1(P2_N926), .IN2(n6809), .Q(n17444) );
  AND2X1 U18767 ( .IN1(P2_N926), .IN2(n6810), .Q(n17445) );
  AND2X1 U18768 ( .IN1(P2_N926), .IN2(n6809), .Q(n17446) );
  AND2X1 U18769 ( .IN1(n17448), .IN2(n6780), .Q(n17447) );
  AND2X1 U18770 ( .IN1(n17450), .IN2(n6779), .Q(n17449) );
  AND2X1 U18771 ( .IN1(n17452), .IN2(n6932), .Q(n17451) );
  AND2X1 U18772 ( .IN1(n17454), .IN2(n6931), .Q(n17453) );
  AND2X1 U18773 ( .IN1(P2_N926), .IN2(n6810), .Q(n17455) );
  AND2X1 U18774 ( .IN1(P2_N926), .IN2(n6809), .Q(n17456) );
  AND2X1 U18775 ( .IN1(P2_N926), .IN2(n6810), .Q(n17457) );
  AND2X1 U18776 ( .IN1(P2_N926), .IN2(n6809), .Q(n17458) );
  AND2X1 U18777 ( .IN1(n17460), .IN2(n6780), .Q(n17459) );
  AND2X1 U18778 ( .IN1(n17462), .IN2(n6779), .Q(n17461) );
  AND2X1 U18779 ( .IN1(n17463), .IN2(n6974), .Q(n14740) );
  AND2X1 U18780 ( .IN1(n17464), .IN2(n6967), .Q(n14741) );
  AND2X1 U18781 ( .IN1(P2_N927), .IN2(n6848), .Q(n17465) );
  AND2X1 U18782 ( .IN1(P2_N927), .IN2(n6807), .Q(n17466) );
  AND2X1 U18783 ( .IN1(P2_N927), .IN2(n6848), .Q(n17467) );
  AND2X1 U18784 ( .IN1(P2_N927), .IN2(n6847), .Q(n17468) );
  AND2X1 U18785 ( .IN1(n17470), .IN2(n6804), .Q(n17469) );
  AND2X1 U18786 ( .IN1(n17472), .IN2(n6803), .Q(n17471) );
  AND2X1 U18787 ( .IN1(P2_N927), .IN2(n6808), .Q(n17473) );
  AND2X1 U18788 ( .IN1(P2_N927), .IN2(n6807), .Q(n17474) );
  AND2X1 U18789 ( .IN1(P2_N927), .IN2(n6848), .Q(n17475) );
  AND2X1 U18790 ( .IN1(P2_N927), .IN2(n6807), .Q(n17476) );
  AND2X1 U18791 ( .IN1(n17478), .IN2(n6804), .Q(n17477) );
  AND2X1 U18792 ( .IN1(n17480), .IN2(n6803), .Q(n17479) );
  AND2X1 U18793 ( .IN1(n17482), .IN2(n6932), .Q(n17481) );
  AND2X1 U18794 ( .IN1(n17484), .IN2(n6931), .Q(n17483) );
  AND2X1 U18795 ( .IN1(P2_N927), .IN2(n6832), .Q(n17485) );
  AND2X1 U18796 ( .IN1(P2_N927), .IN2(n6807), .Q(n17486) );
  AND2X1 U18797 ( .IN1(P2_N927), .IN2(n6832), .Q(n17487) );
  AND2X1 U18798 ( .IN1(P2_N927), .IN2(n6807), .Q(n17488) );
  AND2X1 U18799 ( .IN1(n17490), .IN2(n6804), .Q(n17489) );
  AND2X1 U18800 ( .IN1(n17492), .IN2(n6803), .Q(n17491) );
  AND2X1 U18801 ( .IN1(n17493), .IN2(n6970), .Q(n14742) );
  AND2X1 U18802 ( .IN1(n17494), .IN2(n6967), .Q(n14743) );
  AND2X1 U18803 ( .IN1(P2_N928), .IN2(n6810), .Q(n17495) );
  AND2X1 U18804 ( .IN1(P2_N928), .IN2(n6807), .Q(n17496) );
  AND2X1 U18805 ( .IN1(P2_N928), .IN2(n6808), .Q(n17497) );
  AND2X1 U18806 ( .IN1(P2_N928), .IN2(n6807), .Q(n17498) );
  AND2X1 U18807 ( .IN1(n17500), .IN2(n6804), .Q(n17499) );
  AND2X1 U18808 ( .IN1(n17502), .IN2(n6803), .Q(n17501) );
  AND2X1 U18809 ( .IN1(P2_N928), .IN2(n6810), .Q(n17503) );
  AND2X1 U18810 ( .IN1(P2_N928), .IN2(n6807), .Q(n17504) );
  AND2X1 U18811 ( .IN1(P2_N928), .IN2(n6810), .Q(n17505) );
  AND2X1 U18812 ( .IN1(P2_N928), .IN2(n6807), .Q(n17506) );
  AND2X1 U18813 ( .IN1(n17508), .IN2(n6804), .Q(n17507) );
  AND2X1 U18814 ( .IN1(n17510), .IN2(n6803), .Q(n17509) );
  AND2X1 U18815 ( .IN1(n17512), .IN2(n6932), .Q(n17511) );
  AND2X1 U18630 ( .IN1(P2_N920), .IN2(n6831), .Q(n17258) );
  AND2X1 U18631 ( .IN1(n17260), .IN2(n6780), .Q(n17259) );
  AND2X1 U18632 ( .IN1(n17262), .IN2(n6779), .Q(n17261) );
  AND2X1 U18633 ( .IN1(P2_N920), .IN2(n6832), .Q(n17263) );
  AND2X1 U18634 ( .IN1(P2_N920), .IN2(n6831), .Q(n17264) );
  AND2X1 U18635 ( .IN1(P2_N920), .IN2(n6832), .Q(n17265) );
  AND2X1 U18636 ( .IN1(P2_N920), .IN2(n6831), .Q(n17266) );
  AND2X1 U18637 ( .IN1(n17268), .IN2(n6780), .Q(n17267) );
  AND2X1 U18638 ( .IN1(n17270), .IN2(n6779), .Q(n17269) );
  AND2X1 U18639 ( .IN1(n17272), .IN2(n6940), .Q(n17271) );
  AND2X1 U18640 ( .IN1(n17274), .IN2(n6931), .Q(n17273) );
  AND2X1 U18641 ( .IN1(P2_N920), .IN2(n6832), .Q(n17275) );
  AND2X1 U18642 ( .IN1(P2_N920), .IN2(n6831), .Q(n17276) );
  AND2X1 U18643 ( .IN1(P2_N920), .IN2(n6832), .Q(n17277) );
  AND2X1 U18644 ( .IN1(P2_N920), .IN2(n6831), .Q(n17278) );
  AND2X1 U18645 ( .IN1(n17280), .IN2(n6780), .Q(n17279) );
  AND2X1 U18646 ( .IN1(n17282), .IN2(n6779), .Q(n17281) );
  AND2X1 U18647 ( .IN1(n17283), .IN2(n6972), .Q(n14728) );
  AND2X1 U18648 ( .IN1(n17284), .IN2(n6963), .Q(n14729) );
  AND2X1 U18649 ( .IN1(P2_N921), .IN2(n6832), .Q(n17285) );
  AND2X1 U18650 ( .IN1(P2_N921), .IN2(n6831), .Q(n17286) );
  AND2X1 U18651 ( .IN1(P2_N921), .IN2(n6832), .Q(n17287) );
  AND2X1 U18652 ( .IN1(P2_N921), .IN2(n6831), .Q(n17288) );
  AND2X1 U18653 ( .IN1(n17290), .IN2(n6780), .Q(n17289) );
  AND2X1 U18654 ( .IN1(n17292), .IN2(n6779), .Q(n17291) );
  AND2X1 U18655 ( .IN1(P2_N921), .IN2(n6832), .Q(n17293) );
  AND2X1 U18656 ( .IN1(P2_N921), .IN2(n6831), .Q(n17294) );
  AND2X1 U18657 ( .IN1(P2_N921), .IN2(n6832), .Q(n17295) );
  AND2X1 U18658 ( .IN1(P2_N921), .IN2(n6831), .Q(n17296) );
  AND2X1 U18659 ( .IN1(n17298), .IN2(n6780), .Q(n17297) );
  AND2X1 U18660 ( .IN1(n17300), .IN2(n6779), .Q(n17299) );
  AND2X1 U18661 ( .IN1(n17302), .IN2(n6940), .Q(n17301) );
  AND2X1 U18662 ( .IN1(n17304), .IN2(n6931), .Q(n17303) );
  AND2X1 U18663 ( .IN1(P2_N921), .IN2(n6832), .Q(n17305) );
  AND2X1 U18664 ( .IN1(P2_N921), .IN2(n6831), .Q(n17306) );
  AND2X1 U18665 ( .IN1(P2_N921), .IN2(n6832), .Q(n17307) );
  AND2X1 U18666 ( .IN1(P2_N921), .IN2(n6831), .Q(n17308) );
  AND2X1 U18667 ( .IN1(n17310), .IN2(n6780), .Q(n17309) );
  AND2X1 U18668 ( .IN1(n17312), .IN2(n6779), .Q(n17311) );
  AND2X1 U18669 ( .IN1(n17313), .IN2(n6972), .Q(n14730) );
  AND2X1 U18670 ( .IN1(n17314), .IN2(n6963), .Q(n14731) );
  AND2X1 U18671 ( .IN1(P2_N922), .IN2(n6832), .Q(n17315) );
  AND2X1 U18672 ( .IN1(P2_N922), .IN2(n6831), .Q(n17316) );
  AND2X1 U18673 ( .IN1(P2_N922), .IN2(n6832), .Q(n17317) );
  AND2X1 U18674 ( .IN1(P2_N922), .IN2(n6831), .Q(n17318) );
  AND2X1 U18675 ( .IN1(n17320), .IN2(n6780), .Q(n17319) );
  AND2X1 U18676 ( .IN1(n17322), .IN2(n6779), .Q(n17321) );
  AND2X1 U18677 ( .IN1(P2_N922), .IN2(n6832), .Q(n17323) );
  AND2X1 U18678 ( .IN1(P2_N922), .IN2(n6831), .Q(n17324) );
  AND2X1 U18679 ( .IN1(P2_N922), .IN2(n6832), .Q(n17325) );
  AND2X1 U18680 ( .IN1(P2_N922), .IN2(n6831), .Q(n17326) );
  AND2X1 U18681 ( .IN1(n17328), .IN2(n6780), .Q(n17327) );
  AND2X1 U18682 ( .IN1(n17330), .IN2(n6779), .Q(n17329) );
  AND2X1 U18683 ( .IN1(n17332), .IN2(n6932), .Q(n17331) );
  AND2X1 U18684 ( .IN1(n17334), .IN2(n6931), .Q(n17333) );
  AND2X1 U18685 ( .IN1(P2_N922), .IN2(n6832), .Q(n17335) );
  AND2X1 U18686 ( .IN1(P2_N922), .IN2(n6831), .Q(n17336) );
  AND2X1 U18687 ( .IN1(P2_N922), .IN2(n6832), .Q(n17337) );
  AND2X1 U18688 ( .IN1(P2_N922), .IN2(n6831), .Q(n17338) );
  AND2X1 U18689 ( .IN1(n17340), .IN2(n6780), .Q(n17339) );
  AND2X1 U18690 ( .IN1(n17342), .IN2(n6779), .Q(n17341) );
  AND2X1 U18691 ( .IN1(n17343), .IN2(n6972), .Q(n14732) );
  AND2X1 U18692 ( .IN1(n17344), .IN2(n6963), .Q(n14733) );
  AND2X1 U18693 ( .IN1(P2_N923), .IN2(n6832), .Q(n17345) );
  AND2X1 U18694 ( .IN1(P2_N923), .IN2(n6831), .Q(n17346) );
  AND2X1 U18695 ( .IN1(P2_N923), .IN2(n6832), .Q(n17347) );
  AND2X1 U18696 ( .IN1(P2_N923), .IN2(n6831), .Q(n17348) );
  AND2X1 U18697 ( .IN1(n17350), .IN2(n6780), .Q(n17349) );
  AND2X1 U18698 ( .IN1(n17352), .IN2(n6779), .Q(n17351) );
  AND2X1 U18699 ( .IN1(P2_N923), .IN2(n6832), .Q(n17353) );
  AND2X1 U18700 ( .IN1(P2_N923), .IN2(n6831), .Q(n17354) );
  AND2X1 U18701 ( .IN1(P2_N923), .IN2(n6832), .Q(n17355) );
  AND2X1 U18702 ( .IN1(P2_N923), .IN2(n6831), .Q(n17356) );
  AND2X1 U18703 ( .IN1(n17358), .IN2(n6780), .Q(n17357) );
  AND2X1 U18704 ( .IN1(n17360), .IN2(n6779), .Q(n17359) );
  AND2X1 U18705 ( .IN1(n17362), .IN2(n6940), .Q(n17361) );
  AND2X1 U18706 ( .IN1(n17364), .IN2(n6931), .Q(n17363) );
  AND2X1 U18707 ( .IN1(P2_N923), .IN2(n6832), .Q(n17365) );
  AND2X1 U18708 ( .IN1(P2_N923), .IN2(n6831), .Q(n17366) );
  AND2X1 U18709 ( .IN1(P2_N923), .IN2(n6832), .Q(n17367) );
  AND2X1 U18710 ( .IN1(P2_N923), .IN2(n6831), .Q(n17368) );
  AND2X1 U18711 ( .IN1(n17370), .IN2(n6780), .Q(n17369) );
  AND2X1 U18712 ( .IN1(n17372), .IN2(n6779), .Q(n17371) );
  AND2X1 U18713 ( .IN1(n17373), .IN2(n6972), .Q(n14734) );
  AND2X1 U18714 ( .IN1(n17374), .IN2(n6963), .Q(n14735) );
  AND2X1 U18715 ( .IN1(P2_N924), .IN2(n6832), .Q(n17375) );
  AND2X1 U18716 ( .IN1(P2_N924), .IN2(n6831), .Q(n17376) );
  AND2X1 U18717 ( .IN1(P2_N924), .IN2(n6832), .Q(n17377) );
  AND2X1 U18718 ( .IN1(P2_N924), .IN2(n6831), .Q(n17378) );
  AND2X1 U18719 ( .IN1(n17380), .IN2(n6780), .Q(n17379) );
  AND2X1 U18720 ( .IN1(n17382), .IN2(n6779), .Q(n17381) );
  AND2X1 U18721 ( .IN1(P2_N924), .IN2(n6832), .Q(n17383) );
  AND2X1 U18722 ( .IN1(P2_N924), .IN2(n6831), .Q(n17384) );
  AND2X1 U18537 ( .IN1(n17133), .IN2(n6974), .Q(n14718) );
  AND2X1 U18538 ( .IN1(n17134), .IN2(n6967), .Q(n14719) );
  AND2X1 U18539 ( .IN1(P2_N916), .IN2(n6848), .Q(n17135) );
  AND2X1 U18540 ( .IN1(P2_N916), .IN2(n6847), .Q(n17136) );
  AND2X1 U18541 ( .IN1(P2_N916), .IN2(n6848), .Q(n17137) );
  AND2X1 U18542 ( .IN1(P2_N916), .IN2(n6847), .Q(n17138) );
  AND2X1 U18543 ( .IN1(n17140), .IN2(n6780), .Q(n17139) );
  AND2X1 U18544 ( .IN1(n17142), .IN2(P2_N291), .Q(n17141) );
  AND2X1 U18545 ( .IN1(P2_N916), .IN2(n6848), .Q(n17143) );
  AND2X1 U18546 ( .IN1(P2_N916), .IN2(n6847), .Q(n17144) );
  AND2X1 U18547 ( .IN1(P2_N916), .IN2(n6848), .Q(n17145) );
  AND2X1 U18548 ( .IN1(P2_N916), .IN2(n6847), .Q(n17146) );
  AND2X1 U18549 ( .IN1(n17148), .IN2(n6780), .Q(n17147) );
  AND2X1 U18550 ( .IN1(n17150), .IN2(P2_N291), .Q(n17149) );
  AND2X1 U18551 ( .IN1(n17152), .IN2(n6932), .Q(n17151) );
  AND2X1 U18552 ( .IN1(n17154), .IN2(n6931), .Q(n17153) );
  AND2X1 U18553 ( .IN1(P2_N916), .IN2(n6848), .Q(n17155) );
  AND2X1 U18554 ( .IN1(P2_N916), .IN2(n6847), .Q(n17156) );
  AND2X1 U18555 ( .IN1(P2_N916), .IN2(n6848), .Q(n17157) );
  AND2X1 U18556 ( .IN1(P2_N916), .IN2(n6847), .Q(n17158) );
  AND2X1 U18557 ( .IN1(n17160), .IN2(n6780), .Q(n17159) );
  AND2X1 U18558 ( .IN1(n17162), .IN2(P2_N291), .Q(n17161) );
  AND2X1 U18559 ( .IN1(n17163), .IN2(n6974), .Q(n14720) );
  AND2X1 U18560 ( .IN1(n17164), .IN2(n6967), .Q(n14721) );
  AND2X1 U18561 ( .IN1(P2_N917), .IN2(n6810), .Q(n17165) );
  AND2X1 U18562 ( .IN1(P2_N917), .IN2(n6809), .Q(n17166) );
  AND2X1 U18563 ( .IN1(P2_N917), .IN2(n6810), .Q(n17167) );
  AND2X1 U18564 ( .IN1(P2_N917), .IN2(n6809), .Q(n17168) );
  AND2X1 U18565 ( .IN1(n17170), .IN2(n6780), .Q(n17169) );
  AND2X1 U18566 ( .IN1(n17172), .IN2(P2_N291), .Q(n17171) );
  AND2X1 U18567 ( .IN1(P2_N917), .IN2(n6810), .Q(n17173) );
  AND2X1 U18568 ( .IN1(P2_N917), .IN2(n6809), .Q(n17174) );
  AND2X1 U18569 ( .IN1(P2_N917), .IN2(n6810), .Q(n17175) );
  AND2X1 U18570 ( .IN1(P2_N917), .IN2(n6809), .Q(n17176) );
  AND2X1 U18571 ( .IN1(n17178), .IN2(n6780), .Q(n17177) );
  AND2X1 U18572 ( .IN1(n17180), .IN2(P2_N291), .Q(n17179) );
  AND2X1 U18573 ( .IN1(n17182), .IN2(n6932), .Q(n17181) );
  AND2X1 U18574 ( .IN1(n17184), .IN2(n6931), .Q(n17183) );
  AND2X1 U18575 ( .IN1(P2_N917), .IN2(n6810), .Q(n17185) );
  AND2X1 U18576 ( .IN1(P2_N917), .IN2(n6809), .Q(n17186) );
  AND2X1 U18577 ( .IN1(P2_N917), .IN2(n6810), .Q(n17187) );
  AND2X1 U18578 ( .IN1(P2_N917), .IN2(n6809), .Q(n17188) );
  AND2X1 U18579 ( .IN1(n17190), .IN2(n6780), .Q(n17189) );
  AND2X1 U18580 ( .IN1(n17192), .IN2(P2_N291), .Q(n17191) );
  AND2X1 U18581 ( .IN1(n17193), .IN2(n6970), .Q(n14722) );
  AND2X1 U18582 ( .IN1(n17194), .IN2(n6967), .Q(n14723) );
  AND2X1 U18583 ( .IN1(P2_N918), .IN2(n6810), .Q(n17195) );
  AND2X1 U18584 ( .IN1(P2_N918), .IN2(n6809), .Q(n17196) );
  AND2X1 U18585 ( .IN1(P2_N918), .IN2(n6810), .Q(n17197) );
  AND2X1 U18586 ( .IN1(P2_N918), .IN2(n6809), .Q(n17198) );
  AND2X1 U18587 ( .IN1(n17200), .IN2(n6780), .Q(n17199) );
  AND2X1 U18588 ( .IN1(n17202), .IN2(P2_N291), .Q(n17201) );
  AND2X1 U18589 ( .IN1(P2_N918), .IN2(n6810), .Q(n17203) );
  AND2X1 U18590 ( .IN1(P2_N918), .IN2(n6809), .Q(n17204) );
  AND2X1 U18591 ( .IN1(P2_N918), .IN2(n6810), .Q(n17205) );
  AND2X1 U18592 ( .IN1(P2_N918), .IN2(n6809), .Q(n17206) );
  AND2X1 U18593 ( .IN1(n17208), .IN2(n6780), .Q(n17207) );
  AND2X1 U18594 ( .IN1(n17210), .IN2(P2_N291), .Q(n17209) );
  AND2X1 U18595 ( .IN1(n17212), .IN2(n6932), .Q(n17211) );
  AND2X1 U18596 ( .IN1(n17214), .IN2(n6931), .Q(n17213) );
  AND2X1 U18597 ( .IN1(P2_N918), .IN2(n6810), .Q(n17215) );
  AND2X1 U18598 ( .IN1(P2_N918), .IN2(n6809), .Q(n17216) );
  AND2X1 U18599 ( .IN1(P2_N918), .IN2(n6810), .Q(n17217) );
  AND2X1 U18600 ( .IN1(P2_N918), .IN2(n6809), .Q(n17218) );
  AND2X1 U18601 ( .IN1(n17220), .IN2(n6780), .Q(n17219) );
  AND2X1 U18602 ( .IN1(n17222), .IN2(P2_N291), .Q(n17221) );
  AND2X1 U18603 ( .IN1(n17223), .IN2(n6970), .Q(n14724) );
  AND2X1 U18604 ( .IN1(n17224), .IN2(n6967), .Q(n14725) );
  AND2X1 U18605 ( .IN1(P2_N919), .IN2(n6810), .Q(n17225) );
  AND2X1 U18606 ( .IN1(P2_N919), .IN2(n6809), .Q(n17226) );
  AND2X1 U18607 ( .IN1(P2_N919), .IN2(n6810), .Q(n17227) );
  AND2X1 U18608 ( .IN1(P2_N919), .IN2(n6809), .Q(n17228) );
  AND2X1 U18609 ( .IN1(n17230), .IN2(n6780), .Q(n17229) );
  AND2X1 U18610 ( .IN1(n17232), .IN2(P2_N291), .Q(n17231) );
  AND2X1 U18611 ( .IN1(P2_N919), .IN2(n6810), .Q(n17233) );
  AND2X1 U18612 ( .IN1(P2_N919), .IN2(n6809), .Q(n17234) );
  AND2X1 U18613 ( .IN1(P2_N919), .IN2(n6810), .Q(n17235) );
  AND2X1 U18614 ( .IN1(P2_N919), .IN2(n6809), .Q(n17236) );
  AND2X1 U18615 ( .IN1(n17238), .IN2(n6780), .Q(n17237) );
  AND2X1 U18616 ( .IN1(n17240), .IN2(P2_N291), .Q(n17239) );
  AND2X1 U18617 ( .IN1(n17242), .IN2(n6932), .Q(n17241) );
  AND2X1 U18618 ( .IN1(n17244), .IN2(n6931), .Q(n17243) );
  AND2X1 U18619 ( .IN1(P2_N919), .IN2(n6810), .Q(n17245) );
  AND2X1 U18620 ( .IN1(P2_N919), .IN2(n6809), .Q(n17246) );
  AND2X1 U18621 ( .IN1(P2_N919), .IN2(n6810), .Q(n17247) );
  AND2X1 U18622 ( .IN1(P2_N919), .IN2(n6809), .Q(n17248) );
  AND2X1 U18623 ( .IN1(n17250), .IN2(n6780), .Q(n17249) );
  AND2X1 U18624 ( .IN1(n17252), .IN2(n6779), .Q(n17251) );
  AND2X1 U18625 ( .IN1(n17253), .IN2(n6974), .Q(n14726) );
  AND2X1 U18626 ( .IN1(n17254), .IN2(n6967), .Q(n14727) );
  AND2X1 U18627 ( .IN1(P2_N920), .IN2(n6832), .Q(n17255) );
  AND2X1 U18628 ( .IN1(P2_N920), .IN2(n6831), .Q(n17256) );
  AND2X1 U18629 ( .IN1(P2_N920), .IN2(n6832), .Q(n17257) );
  AND2X1 U18444 ( .IN1(n17007), .IN2(n6974), .Q(n14703) );
  AND2X1 U18445 ( .IN1(P2_N1260), .IN2(n6803), .Q(n17008) );
  AND2X1 U18446 ( .IN1(n16806), .IN2(n6804), .Q(n17009) );
  AND2X1 U18447 ( .IN1(n16820), .IN2(n6931), .Q(n17010) );
  AND2X1 U18448 ( .IN1(n17012), .IN2(n6932), .Q(n17011) );
  AND2X1 U18449 ( .IN1(n16833), .IN2(n6967), .Q(n14704) );
  AND2X1 U18450 ( .IN1(n17013), .IN2(n6970), .Q(n14705) );
  AND2X1 U18451 ( .IN1(P2_N812), .IN2(n6838), .Q(n17014) );
  AND2X1 U18452 ( .IN1(P2_N1158), .IN2(n6837), .Q(n17015) );
  AND2X1 U18453 ( .IN1(n17017), .IN2(n6794), .Q(n17016) );
  AND2X1 U18454 ( .IN1(n6793), .IN2(n17019), .Q(n17018) );
  AND2X1 U18455 ( .IN1(P2_N1786), .IN2(n6834), .Q(n17020) );
  AND2X1 U18456 ( .IN1(P2_N2532), .IN2(n7484), .Q(n17021) );
  AND2X1 U18457 ( .IN1(P2_N2159), .IN2(n6834), .Q(n17022) );
  AND2X1 U18458 ( .IN1(P2_N2905), .IN2(n7484), .Q(n17023) );
  AND2X1 U18459 ( .IN1(n17025), .IN2(n6802), .Q(n17024) );
  AND2X1 U18460 ( .IN1(n17027), .IN2(n6779), .Q(n17026) );
  AND2X1 U18461 ( .IN1(n17029), .IN2(n6934), .Q(n17028) );
  AND2X1 U18462 ( .IN1(n17031), .IN2(n6943), .Q(n17030) );
  AND2X1 U18463 ( .IN1(P2_N3278), .IN2(n6838), .Q(n17032) );
  AND2X1 U18464 ( .IN1(P2_N4055), .IN2(n7485), .Q(n17033) );
  AND2X1 U18465 ( .IN1(P2_N3651), .IN2(n6838), .Q(n17034) );
  AND2X1 U18466 ( .IN1(n7397), .IN2(n7485), .Q(n17035) );
  AND2X1 U18467 ( .IN1(n17037), .IN2(n6802), .Q(n17036) );
  AND2X1 U18468 ( .IN1(n17039), .IN2(P2_N291), .Q(n17038) );
  AND2X1 U18469 ( .IN1(n17041), .IN2(n6934), .Q(n17040) );
  AND2X1 U18470 ( .IN1(n14706), .IN2(n6943), .Q(n17042) );
  AND2X1 U18471 ( .IN1(n17043), .IN2(n6966), .Q(n14708) );
  AND2X1 U18472 ( .IN1(n17044), .IN2(P2_N294), .Q(n14709) );
  AND2X1 U18473 ( .IN1(P2_N843), .IN2(n6838), .Q(n17045) );
  AND2X1 U18474 ( .IN1(P2_N1189), .IN2(n6837), .Q(n17046) );
  AND2X1 U18475 ( .IN1(n17048), .IN2(n6784), .Q(n17047) );
  AND2X1 U18476 ( .IN1(n14711), .IN2(n6793), .Q(n17049) );
  AND2X1 U18477 ( .IN1(P2_N1817), .IN2(n6834), .Q(n17050) );
  AND2X1 U18478 ( .IN1(P2_N2563), .IN2(n7484), .Q(n17051) );
  AND2X1 U18479 ( .IN1(P2_N2190), .IN2(n6834), .Q(n17052) );
  AND2X1 U18480 ( .IN1(P2_N2936), .IN2(n7484), .Q(n17053) );
  AND2X1 U18481 ( .IN1(n17055), .IN2(n6802), .Q(n17054) );
  AND2X1 U18482 ( .IN1(n17057), .IN2(n6803), .Q(n17056) );
  AND2X1 U18483 ( .IN1(n17059), .IN2(n6934), .Q(n17058) );
  AND2X1 U18484 ( .IN1(n17061), .IN2(n6943), .Q(n17060) );
  AND2X1 U18485 ( .IN1(P2_N3309), .IN2(n6820), .Q(n17062) );
  AND2X1 U18486 ( .IN1(P2_N4024), .IN2(n7485), .Q(n17063) );
  AND2X1 U18487 ( .IN1(P2_N3682), .IN2(n6828), .Q(n17064) );
  AND2X1 U18488 ( .IN1(P2_N4428), .IN2(n7485), .Q(n17065) );
  AND2X1 U18489 ( .IN1(n17067), .IN2(n6802), .Q(n17066) );
  AND2X1 U18490 ( .IN1(n17069), .IN2(n6803), .Q(n17068) );
  AND2X1 U18491 ( .IN1(n17071), .IN2(n6934), .Q(n17070) );
  AND2X1 U18492 ( .IN1(n14710), .IN2(n6943), .Q(n17072) );
  AND2X1 U18493 ( .IN1(n17073), .IN2(n6966), .Q(n14712) );
  AND2X1 U18494 ( .IN1(n17074), .IN2(P2_N294), .Q(n14713) );
  AND2X1 U18495 ( .IN1(P2_N842), .IN2(n6838), .Q(n17075) );
  AND2X1 U18496 ( .IN1(P2_N1188), .IN2(n6837), .Q(n17076) );
  AND2X1 U18497 ( .IN1(n17078), .IN2(n6784), .Q(n17077) );
  AND2X1 U18498 ( .IN1(n14715), .IN2(n6793), .Q(n17079) );
  AND2X1 U18499 ( .IN1(P2_N1816), .IN2(n6834), .Q(n17080) );
  AND2X1 U18500 ( .IN1(P2_N2562), .IN2(n7484), .Q(n17081) );
  AND2X1 U18501 ( .IN1(P2_N2189), .IN2(n6848), .Q(n17082) );
  AND2X1 U18502 ( .IN1(P2_N2935), .IN2(n6847), .Q(n17083) );
  AND2X1 U18503 ( .IN1(n17085), .IN2(n6782), .Q(n17084) );
  AND2X1 U18504 ( .IN1(n17087), .IN2(P2_N291), .Q(n17086) );
  AND2X1 U18505 ( .IN1(n17089), .IN2(n6934), .Q(n17088) );
  AND2X1 U18506 ( .IN1(n17091), .IN2(n6943), .Q(n17090) );
  AND2X1 U18507 ( .IN1(P2_N3308), .IN2(n6842), .Q(n17092) );
  AND2X1 U18508 ( .IN1(P2_N4054), .IN2(n7485), .Q(n17093) );
  AND2X1 U18509 ( .IN1(P2_N3681), .IN2(n6842), .Q(n17094) );
  AND2X1 U18510 ( .IN1(P2_N4398), .IN2(n7485), .Q(n17095) );
  AND2X1 U18511 ( .IN1(n17097), .IN2(n6782), .Q(n17096) );
  AND2X1 U18512 ( .IN1(n17099), .IN2(P2_N291), .Q(n17098) );
  AND2X1 U18513 ( .IN1(n17101), .IN2(n6934), .Q(n17100) );
  AND2X1 U18514 ( .IN1(n14714), .IN2(n6943), .Q(n17102) );
  AND2X1 U18515 ( .IN1(n17103), .IN2(n6966), .Q(n14716) );
  AND2X1 U18516 ( .IN1(n17104), .IN2(P2_N294), .Q(n14717) );
  AND2X1 U18517 ( .IN1(P2_N915), .IN2(n6848), .Q(n17105) );
  AND2X1 U18518 ( .IN1(P2_N915), .IN2(n6847), .Q(n17106) );
  AND2X1 U18519 ( .IN1(P2_N915), .IN2(n6848), .Q(n17107) );
  AND2X1 U18520 ( .IN1(P2_N915), .IN2(n6847), .Q(n17108) );
  AND2X1 U18521 ( .IN1(n17110), .IN2(n6780), .Q(n17109) );
  AND2X1 U18522 ( .IN1(n17112), .IN2(P2_N291), .Q(n17111) );
  AND2X1 U18523 ( .IN1(P2_N915), .IN2(n6848), .Q(n17113) );
  AND2X1 U18524 ( .IN1(P2_N915), .IN2(n6847), .Q(n17114) );
  AND2X1 U18525 ( .IN1(P2_N915), .IN2(n6848), .Q(n17115) );
  AND2X1 U18526 ( .IN1(P2_N915), .IN2(n6847), .Q(n17116) );
  AND2X1 U18527 ( .IN1(n17118), .IN2(n6780), .Q(n17117) );
  AND2X1 U18528 ( .IN1(n17120), .IN2(P2_N291), .Q(n17119) );
  AND2X1 U18529 ( .IN1(n17122), .IN2(n6932), .Q(n17121) );
  AND2X1 U18530 ( .IN1(n17124), .IN2(n6931), .Q(n17123) );
  AND2X1 U18531 ( .IN1(P2_N915), .IN2(n6848), .Q(n17125) );
  AND2X1 U18532 ( .IN1(P2_N915), .IN2(n6847), .Q(n17126) );
  AND2X1 U18533 ( .IN1(P2_N915), .IN2(n6848), .Q(n17127) );
  AND2X1 U18534 ( .IN1(P2_N915), .IN2(n6847), .Q(n17128) );
  AND2X1 U18535 ( .IN1(n17130), .IN2(n6780), .Q(n17129) );
  AND2X1 U18536 ( .IN1(n17132), .IN2(P2_N291), .Q(n17131) );
  AND2X1 U18351 ( .IN1(n16292), .IN2(n6937), .Q(n16914) );
  AND2X1 U18352 ( .IN1(n16916), .IN2(n6946), .Q(n16915) );
  AND2X1 U18353 ( .IN1(n16305), .IN2(n6967), .Q(n14672) );
  AND2X1 U18354 ( .IN1(n16917), .IN2(n6974), .Q(n14673) );
  AND2X1 U18355 ( .IN1(P2_N1245), .IN2(n6789), .Q(n16918) );
  AND2X1 U18356 ( .IN1(n16311), .IN2(n6790), .Q(n16919) );
  AND2X1 U18357 ( .IN1(n16325), .IN2(n6937), .Q(n16920) );
  AND2X1 U18358 ( .IN1(n16922), .IN2(n6948), .Q(n16921) );
  AND2X1 U18359 ( .IN1(n16338), .IN2(n6969), .Q(n14674) );
  AND2X1 U18360 ( .IN1(n16923), .IN2(n6970), .Q(n14675) );
  AND2X1 U18361 ( .IN1(P2_N1246), .IN2(n6789), .Q(n16924) );
  AND2X1 U18362 ( .IN1(n16344), .IN2(n6790), .Q(n16925) );
  AND2X1 U18363 ( .IN1(n16358), .IN2(n6937), .Q(n16926) );
  AND2X1 U18364 ( .IN1(n16928), .IN2(n6946), .Q(n16927) );
  AND2X1 U18365 ( .IN1(n16371), .IN2(n6969), .Q(n14676) );
  AND2X1 U18366 ( .IN1(n16929), .IN2(n6970), .Q(n14677) );
  AND2X1 U18367 ( .IN1(P2_N1247), .IN2(n6789), .Q(n16930) );
  AND2X1 U18368 ( .IN1(n16377), .IN2(n6790), .Q(n16931) );
  AND2X1 U18369 ( .IN1(n16391), .IN2(n6937), .Q(n16932) );
  AND2X1 U18370 ( .IN1(n16934), .IN2(n6948), .Q(n16933) );
  AND2X1 U18371 ( .IN1(n16404), .IN2(n6969), .Q(n14678) );
  AND2X1 U18372 ( .IN1(n16935), .IN2(n6970), .Q(n14679) );
  AND2X1 U18373 ( .IN1(P2_N1248), .IN2(n6789), .Q(n16936) );
  AND2X1 U18374 ( .IN1(n16410), .IN2(n6790), .Q(n16937) );
  AND2X1 U18375 ( .IN1(n16424), .IN2(n6937), .Q(n16938) );
  AND2X1 U18376 ( .IN1(n16940), .IN2(n6948), .Q(n16939) );
  AND2X1 U18377 ( .IN1(n16437), .IN2(n6969), .Q(n14680) );
  AND2X1 U18378 ( .IN1(n16941), .IN2(n6970), .Q(n14681) );
  AND2X1 U18379 ( .IN1(P2_N1249), .IN2(n6793), .Q(n16942) );
  AND2X1 U18380 ( .IN1(n16443), .IN2(n6784), .Q(n16943) );
  AND2X1 U18381 ( .IN1(n16457), .IN2(n6931), .Q(n16944) );
  AND2X1 U18382 ( .IN1(n16946), .IN2(n6940), .Q(n16945) );
  AND2X1 U18383 ( .IN1(n16470), .IN2(n6969), .Q(n14682) );
  AND2X1 U18384 ( .IN1(n16947), .IN2(n6970), .Q(n14683) );
  AND2X1 U18385 ( .IN1(P2_N1250), .IN2(n7488), .Q(n16948) );
  AND2X1 U18386 ( .IN1(n16476), .IN2(n6784), .Q(n16949) );
  AND2X1 U18387 ( .IN1(n16490), .IN2(n6943), .Q(n16950) );
  AND2X1 U18388 ( .IN1(n16952), .IN2(n6940), .Q(n16951) );
  AND2X1 U18389 ( .IN1(n16503), .IN2(n6963), .Q(n14684) );
  AND2X1 U18390 ( .IN1(n16953), .IN2(n6972), .Q(n14685) );
  AND2X1 U18391 ( .IN1(P2_N1251), .IN2(n7488), .Q(n16954) );
  AND2X1 U18392 ( .IN1(n16509), .IN2(n6784), .Q(n16955) );
  AND2X1 U18393 ( .IN1(n16523), .IN2(n6943), .Q(n16956) );
  AND2X1 U18394 ( .IN1(n16958), .IN2(n6940), .Q(n16957) );
  AND2X1 U18395 ( .IN1(n16536), .IN2(n6963), .Q(n14686) );
  AND2X1 U18396 ( .IN1(n16959), .IN2(n6972), .Q(n14687) );
  AND2X1 U18397 ( .IN1(P2_N1252), .IN2(n6793), .Q(n16960) );
  AND2X1 U18398 ( .IN1(n16542), .IN2(n6784), .Q(n16961) );
  AND2X1 U18399 ( .IN1(n16556), .IN2(n7460), .Q(n16962) );
  AND2X1 U18400 ( .IN1(n16964), .IN2(n6934), .Q(n16963) );
  AND2X1 U18401 ( .IN1(n16569), .IN2(P2_N294), .Q(n14688) );
  AND2X1 U18402 ( .IN1(n16965), .IN2(n6966), .Q(n14689) );
  AND2X1 U18403 ( .IN1(P2_N1253), .IN2(P2_N291), .Q(n16966) );
  AND2X1 U18404 ( .IN1(n16575), .IN2(n6802), .Q(n16967) );
  AND2X1 U18405 ( .IN1(n16589), .IN2(n7460), .Q(n16968) );
  AND2X1 U18406 ( .IN1(n16970), .IN2(n6934), .Q(n16969) );
  AND2X1 U18407 ( .IN1(n16602), .IN2(P2_N294), .Q(n14690) );
  AND2X1 U18408 ( .IN1(n16971), .IN2(n6966), .Q(n14691) );
  AND2X1 U18409 ( .IN1(P2_N1254), .IN2(P2_N291), .Q(n16972) );
  AND2X1 U18410 ( .IN1(n16608), .IN2(n6802), .Q(n16973) );
  AND2X1 U18411 ( .IN1(n16622), .IN2(n7460), .Q(n16974) );
  AND2X1 U18412 ( .IN1(n16976), .IN2(n6934), .Q(n16975) );
  AND2X1 U18413 ( .IN1(n16635), .IN2(P2_N294), .Q(n14692) );
  AND2X1 U18414 ( .IN1(n16977), .IN2(n6966), .Q(n14693) );
  AND2X1 U18415 ( .IN1(P2_N1255), .IN2(P2_N291), .Q(n16978) );
  AND2X1 U18416 ( .IN1(n16641), .IN2(n6802), .Q(n16979) );
  AND2X1 U18417 ( .IN1(n16655), .IN2(n7460), .Q(n16980) );
  AND2X1 U18418 ( .IN1(n16982), .IN2(n6934), .Q(n16981) );
  AND2X1 U18419 ( .IN1(n16668), .IN2(P2_N294), .Q(n14694) );
  AND2X1 U18420 ( .IN1(n16983), .IN2(n6966), .Q(n14695) );
  AND2X1 U18421 ( .IN1(P2_N1256), .IN2(n6781), .Q(n16984) );
  AND2X1 U18422 ( .IN1(n16674), .IN2(n6782), .Q(n16985) );
  AND2X1 U18423 ( .IN1(n16688), .IN2(n7460), .Q(n16986) );
  AND2X1 U18424 ( .IN1(n16988), .IN2(n6934), .Q(n16987) );
  AND2X1 U18425 ( .IN1(n16701), .IN2(P2_N294), .Q(n14696) );
  AND2X1 U18426 ( .IN1(n16989), .IN2(n6966), .Q(n14697) );
  AND2X1 U18427 ( .IN1(P2_N1257), .IN2(n6781), .Q(n16990) );
  AND2X1 U18428 ( .IN1(n16707), .IN2(n6782), .Q(n16991) );
  AND2X1 U18429 ( .IN1(n16721), .IN2(n7460), .Q(n16992) );
  AND2X1 U18430 ( .IN1(n16994), .IN2(n6934), .Q(n16993) );
  AND2X1 U18431 ( .IN1(n16734), .IN2(P2_N294), .Q(n14698) );
  AND2X1 U18432 ( .IN1(n16995), .IN2(n6966), .Q(n14699) );
  AND2X1 U18433 ( .IN1(P2_N1258), .IN2(n6781), .Q(n16996) );
  AND2X1 U18434 ( .IN1(n16740), .IN2(n6782), .Q(n16997) );
  AND2X1 U18435 ( .IN1(n16754), .IN2(n6943), .Q(n16998) );
  AND2X1 U18436 ( .IN1(n17000), .IN2(n6932), .Q(n16999) );
  AND2X1 U18437 ( .IN1(n16767), .IN2(P2_N294), .Q(n14700) );
  AND2X1 U18438 ( .IN1(n17001), .IN2(n6966), .Q(n14701) );
  AND2X1 U18439 ( .IN1(P2_N1259), .IN2(n6803), .Q(n17002) );
  AND2X1 U18440 ( .IN1(n16773), .IN2(n6804), .Q(n17003) );
  AND2X1 U18441 ( .IN1(n16787), .IN2(n6943), .Q(n17004) );
  AND2X1 U18442 ( .IN1(n17006), .IN2(n6932), .Q(n17005) );
  AND2X1 U18443 ( .IN1(n16800), .IN2(n6967), .Q(n14702) );
  AND2X1 U18258 ( .IN1(n16816), .IN2(n6803), .Q(n16815) );
  AND2X1 U18259 ( .IN1(n16818), .IN2(n6932), .Q(n16817) );
  AND2X1 U18260 ( .IN1(n16820), .IN2(n6931), .Q(n16819) );
  AND2X1 U18261 ( .IN1(P2_N3159), .IN2(n6834), .Q(n16821) );
  AND2X1 U18262 ( .IN1(P2_N3905), .IN2(n7484), .Q(n16822) );
  AND2X1 U18263 ( .IN1(P2_N3532), .IN2(n6834), .Q(n16823) );
  AND2X1 U18264 ( .IN1(P2_N4307), .IN2(n7484), .Q(n16824) );
  AND2X1 U18265 ( .IN1(n16826), .IN2(n6804), .Q(n16825) );
  AND2X1 U18266 ( .IN1(n16828), .IN2(n6803), .Q(n16827) );
  AND2X1 U18267 ( .IN1(P2_N4528), .IN2(n6943), .Q(n16829) );
  AND2X1 U18268 ( .IN1(n16831), .IN2(n6932), .Q(n16830) );
  AND2X1 U18269 ( .IN1(n16832), .IN2(n6974), .Q(n14644) );
  AND2X1 U18270 ( .IN1(n16833), .IN2(n6967), .Q(n14645) );
  AND2X1 U18271 ( .IN1(P2_N1231), .IN2(n6775), .Q(n16834) );
  AND2X1 U18272 ( .IN1(n15849), .IN2(n6776), .Q(n16835) );
  AND2X1 U18273 ( .IN1(n15863), .IN2(n6937), .Q(n16836) );
  AND2X1 U18274 ( .IN1(n16838), .IN2(n6946), .Q(n16837) );
  AND2X1 U18275 ( .IN1(n15876), .IN2(n6967), .Q(n14646) );
  AND2X1 U18276 ( .IN1(n16839), .IN2(n6974), .Q(n14647) );
  AND2X1 U18277 ( .IN1(P2_N1232), .IN2(n6775), .Q(n16840) );
  AND2X1 U18278 ( .IN1(n15882), .IN2(n6776), .Q(n16841) );
  AND2X1 U18279 ( .IN1(n15896), .IN2(n6941), .Q(n16842) );
  AND2X1 U18280 ( .IN1(n16844), .IN2(n6942), .Q(n16843) );
  AND2X1 U18281 ( .IN1(n15909), .IN2(n6967), .Q(n14648) );
  AND2X1 U18282 ( .IN1(n16845), .IN2(n6974), .Q(n14649) );
  AND2X1 U18283 ( .IN1(P2_N1233), .IN2(n6775), .Q(n16846) );
  AND2X1 U18284 ( .IN1(n15915), .IN2(n6776), .Q(n16847) );
  AND2X1 U18285 ( .IN1(n15929), .IN2(n6941), .Q(n16848) );
  AND2X1 U18286 ( .IN1(n16850), .IN2(n6942), .Q(n16849) );
  AND2X1 U18287 ( .IN1(n15942), .IN2(n6967), .Q(n14650) );
  AND2X1 U18288 ( .IN1(n16851), .IN2(n6974), .Q(n14651) );
  AND2X1 U18289 ( .IN1(P2_N1234), .IN2(n6775), .Q(n16852) );
  AND2X1 U18290 ( .IN1(n15948), .IN2(n6776), .Q(n16853) );
  AND2X1 U18291 ( .IN1(n15962), .IN2(n6941), .Q(n16854) );
  AND2X1 U18292 ( .IN1(n16856), .IN2(n6942), .Q(n16855) );
  AND2X1 U18293 ( .IN1(n15975), .IN2(n6963), .Q(n14652) );
  AND2X1 U18294 ( .IN1(n16857), .IN2(n6970), .Q(n14653) );
  AND2X1 U18295 ( .IN1(P2_N1235), .IN2(n7487), .Q(n16858) );
  AND2X1 U18296 ( .IN1(n15981), .IN2(n6790), .Q(n16859) );
  AND2X1 U18297 ( .IN1(n15995), .IN2(P2_N293), .Q(n16860) );
  AND2X1 U18298 ( .IN1(n16862), .IN2(n6948), .Q(n16861) );
  AND2X1 U18299 ( .IN1(n16008), .IN2(n6963), .Q(n14654) );
  AND2X1 U18300 ( .IN1(n16863), .IN2(n6970), .Q(n14655) );
  AND2X1 U18301 ( .IN1(P2_N1236), .IN2(n7487), .Q(n16864) );
  AND2X1 U18302 ( .IN1(n16014), .IN2(n6786), .Q(n16865) );
  AND2X1 U18303 ( .IN1(n16028), .IN2(P2_N293), .Q(n16866) );
  AND2X1 U18304 ( .IN1(n16868), .IN2(n6946), .Q(n16867) );
  AND2X1 U18305 ( .IN1(n16041), .IN2(n6963), .Q(n14656) );
  AND2X1 U18306 ( .IN1(n16869), .IN2(n6970), .Q(n14657) );
  AND2X1 U18307 ( .IN1(P2_N1237), .IN2(n7487), .Q(n16870) );
  AND2X1 U18308 ( .IN1(n16047), .IN2(n6790), .Q(n16871) );
  AND2X1 U18309 ( .IN1(n16061), .IN2(P2_N293), .Q(n16872) );
  AND2X1 U18310 ( .IN1(n16874), .IN2(n6946), .Q(n16873) );
  AND2X1 U18311 ( .IN1(n16074), .IN2(n6963), .Q(n14658) );
  AND2X1 U18312 ( .IN1(n16875), .IN2(n6970), .Q(n14659) );
  AND2X1 U18313 ( .IN1(P2_N1238), .IN2(n6787), .Q(n16876) );
  AND2X1 U18314 ( .IN1(n16080), .IN2(n6786), .Q(n16877) );
  AND2X1 U18315 ( .IN1(n16094), .IN2(P2_N293), .Q(n16878) );
  AND2X1 U18316 ( .IN1(n16880), .IN2(n6942), .Q(n16879) );
  AND2X1 U18317 ( .IN1(n16107), .IN2(n6963), .Q(n14660) );
  AND2X1 U18318 ( .IN1(n16881), .IN2(n6970), .Q(n14661) );
  AND2X1 U18319 ( .IN1(P2_N1239), .IN2(n6787), .Q(n16882) );
  AND2X1 U18320 ( .IN1(n16113), .IN2(n6786), .Q(n16883) );
  AND2X1 U18321 ( .IN1(n16127), .IN2(P2_N293), .Q(n16884) );
  AND2X1 U18322 ( .IN1(n16886), .IN2(n6946), .Q(n16885) );
  AND2X1 U18323 ( .IN1(n16140), .IN2(n6963), .Q(n14662) );
  AND2X1 U18324 ( .IN1(n16887), .IN2(n6970), .Q(n14663) );
  AND2X1 U18325 ( .IN1(P2_N1240), .IN2(n6787), .Q(n16888) );
  AND2X1 U18326 ( .IN1(n16146), .IN2(n6790), .Q(n16889) );
  AND2X1 U18327 ( .IN1(n16160), .IN2(P2_N293), .Q(n16890) );
  AND2X1 U18328 ( .IN1(n16892), .IN2(n6948), .Q(n16891) );
  AND2X1 U18329 ( .IN1(n16173), .IN2(n6963), .Q(n14664) );
  AND2X1 U18330 ( .IN1(n16893), .IN2(n6970), .Q(n14665) );
  AND2X1 U18331 ( .IN1(P2_N1241), .IN2(n6787), .Q(n16894) );
  AND2X1 U18332 ( .IN1(n16179), .IN2(n6790), .Q(n16895) );
  AND2X1 U18333 ( .IN1(n16193), .IN2(P2_N293), .Q(n16896) );
  AND2X1 U18334 ( .IN1(n16898), .IN2(n6948), .Q(n16897) );
  AND2X1 U18335 ( .IN1(n16206), .IN2(n6963), .Q(n14666) );
  AND2X1 U18336 ( .IN1(n16899), .IN2(n6974), .Q(n14667) );
  AND2X1 U18337 ( .IN1(P2_N1242), .IN2(n6789), .Q(n16900) );
  AND2X1 U18338 ( .IN1(n16212), .IN2(n6786), .Q(n16901) );
  AND2X1 U18339 ( .IN1(n16226), .IN2(n6937), .Q(n16902) );
  AND2X1 U18340 ( .IN1(n16904), .IN2(n6946), .Q(n16903) );
  AND2X1 U18341 ( .IN1(n16239), .IN2(n6967), .Q(n14668) );
  AND2X1 U18342 ( .IN1(n16905), .IN2(n6974), .Q(n14669) );
  AND2X1 U18343 ( .IN1(P2_N1243), .IN2(n6789), .Q(n16906) );
  AND2X1 U18344 ( .IN1(n16245), .IN2(n6786), .Q(n16907) );
  AND2X1 U18345 ( .IN1(n16259), .IN2(n6941), .Q(n16908) );
  AND2X1 U18346 ( .IN1(n16910), .IN2(n6946), .Q(n16909) );
  AND2X1 U18347 ( .IN1(n16272), .IN2(n6967), .Q(n14670) );
  AND2X1 U18348 ( .IN1(n16911), .IN2(n6974), .Q(n14671) );
  AND2X1 U18349 ( .IN1(P2_N1244), .IN2(n6789), .Q(n16912) );
  AND2X1 U18350 ( .IN1(n16278), .IN2(n6786), .Q(n16913) );
  AND2X1 U18165 ( .IN1(P2_N3155), .IN2(n6830), .Q(n16689) );
  AND2X1 U18166 ( .IN1(P2_N3901), .IN2(n6829), .Q(n16690) );
  AND2X1 U18167 ( .IN1(P2_N3528), .IN2(n6830), .Q(n16691) );
  AND2X1 U18168 ( .IN1(P2_N4303), .IN2(n6829), .Q(n16692) );
  AND2X1 U18169 ( .IN1(n16694), .IN2(n6794), .Q(n16693) );
  AND2X1 U18170 ( .IN1(n16696), .IN2(n6793), .Q(n16695) );
  AND2X1 U18171 ( .IN1(P2_N4524), .IN2(n6943), .Q(n16697) );
  AND2X1 U18172 ( .IN1(n16699), .IN2(n6934), .Q(n16698) );
  AND2X1 U18173 ( .IN1(n16700), .IN2(n6966), .Q(n14636) );
  AND2X1 U18174 ( .IN1(n16701), .IN2(P2_N294), .Q(n14637) );
  AND2X1 U18175 ( .IN1(P2_N656), .IN2(n6828), .Q(n16702) );
  AND2X1 U18176 ( .IN1(P2_N1002), .IN2(n7485), .Q(n16703) );
  AND2X1 U18177 ( .IN1(P2_N390), .IN2(n6828), .Q(n16704) );
  AND2X1 U18178 ( .IN1(P2_N1257), .IN2(n7485), .Q(n16705) );
  AND2X1 U18179 ( .IN1(n16707), .IN2(n6782), .Q(n16706) );
  AND2X1 U18180 ( .IN1(n16709), .IN2(n6781), .Q(n16708) );
  AND2X1 U18181 ( .IN1(P2_N1664), .IN2(n6830), .Q(n16710) );
  AND2X1 U18182 ( .IN1(P2_N2410), .IN2(n6829), .Q(n16711) );
  AND2X1 U18183 ( .IN1(P2_N2037), .IN2(n6830), .Q(n16712) );
  AND2X1 U18184 ( .IN1(P2_N2783), .IN2(n6829), .Q(n16713) );
  AND2X1 U18185 ( .IN1(n16715), .IN2(n6794), .Q(n16714) );
  AND2X1 U18186 ( .IN1(n16717), .IN2(n6793), .Q(n16716) );
  AND2X1 U18187 ( .IN1(n16719), .IN2(n6934), .Q(n16718) );
  AND2X1 U18188 ( .IN1(n16721), .IN2(n7460), .Q(n16720) );
  AND2X1 U18189 ( .IN1(P2_N3156), .IN2(n6830), .Q(n16722) );
  AND2X1 U18190 ( .IN1(P2_N3902), .IN2(n6829), .Q(n16723) );
  AND2X1 U18191 ( .IN1(P2_N3529), .IN2(n6830), .Q(n16724) );
  AND2X1 U18192 ( .IN1(P2_N4304), .IN2(n6829), .Q(n16725) );
  AND2X1 U18193 ( .IN1(n16727), .IN2(n6804), .Q(n16726) );
  AND2X1 U18194 ( .IN1(n16729), .IN2(n6803), .Q(n16728) );
  AND2X1 U18195 ( .IN1(P2_N4525), .IN2(n6943), .Q(n16730) );
  AND2X1 U18196 ( .IN1(n16732), .IN2(n6932), .Q(n16731) );
  AND2X1 U18197 ( .IN1(n16733), .IN2(n6966), .Q(n14638) );
  AND2X1 U18198 ( .IN1(n16734), .IN2(P2_N294), .Q(n14639) );
  AND2X1 U18199 ( .IN1(P2_N657), .IN2(n6820), .Q(n16735) );
  AND2X1 U18200 ( .IN1(P2_N1003), .IN2(n7485), .Q(n16736) );
  AND2X1 U18201 ( .IN1(P2_N391), .IN2(n6828), .Q(n16737) );
  AND2X1 U18202 ( .IN1(P2_N1258), .IN2(n7485), .Q(n16738) );
  AND2X1 U18203 ( .IN1(n16740), .IN2(n6782), .Q(n16739) );
  AND2X1 U18204 ( .IN1(n16742), .IN2(n6781), .Q(n16741) );
  AND2X1 U18205 ( .IN1(P2_N1665), .IN2(n6834), .Q(n16743) );
  AND2X1 U18206 ( .IN1(P2_N2411), .IN2(n7484), .Q(n16744) );
  AND2X1 U18207 ( .IN1(P2_N2038), .IN2(n6834), .Q(n16745) );
  AND2X1 U18208 ( .IN1(P2_N2784), .IN2(n7484), .Q(n16746) );
  AND2X1 U18209 ( .IN1(n16748), .IN2(n6804), .Q(n16747) );
  AND2X1 U18210 ( .IN1(n16750), .IN2(n6803), .Q(n16749) );
  AND2X1 U18211 ( .IN1(n16752), .IN2(n6932), .Q(n16751) );
  AND2X1 U18212 ( .IN1(n16754), .IN2(n6943), .Q(n16753) );
  AND2X1 U18213 ( .IN1(P2_N3157), .IN2(n6834), .Q(n16755) );
  AND2X1 U18214 ( .IN1(P2_N3903), .IN2(n7484), .Q(n16756) );
  AND2X1 U18215 ( .IN1(P2_N3530), .IN2(n6834), .Q(n16757) );
  AND2X1 U18216 ( .IN1(P2_N4305), .IN2(n7484), .Q(n16758) );
  AND2X1 U18217 ( .IN1(n16760), .IN2(n6804), .Q(n16759) );
  AND2X1 U18218 ( .IN1(n16762), .IN2(n6803), .Q(n16761) );
  AND2X1 U18219 ( .IN1(P2_N4526), .IN2(n6943), .Q(n16763) );
  AND2X1 U18220 ( .IN1(n16765), .IN2(n6932), .Q(n16764) );
  AND2X1 U18221 ( .IN1(n16766), .IN2(n6966), .Q(n14640) );
  AND2X1 U18222 ( .IN1(n16767), .IN2(P2_N294), .Q(n14641) );
  AND2X1 U18223 ( .IN1(P2_N658), .IN2(n6828), .Q(n16768) );
  AND2X1 U18224 ( .IN1(P2_N1004), .IN2(n7485), .Q(n16769) );
  AND2X1 U18225 ( .IN1(P2_N392), .IN2(n6820), .Q(n16770) );
  AND2X1 U18226 ( .IN1(P2_N1259), .IN2(n7485), .Q(n16771) );
  AND2X1 U18227 ( .IN1(n16773), .IN2(n6804), .Q(n16772) );
  AND2X1 U18228 ( .IN1(n16775), .IN2(n6803), .Q(n16774) );
  AND2X1 U18229 ( .IN1(P2_N1666), .IN2(n6834), .Q(n16776) );
  AND2X1 U18230 ( .IN1(P2_N2412), .IN2(n7484), .Q(n16777) );
  AND2X1 U18231 ( .IN1(P2_N2039), .IN2(n6834), .Q(n16778) );
  AND2X1 U18232 ( .IN1(P2_N2785), .IN2(n7484), .Q(n16779) );
  AND2X1 U18233 ( .IN1(n16781), .IN2(n6804), .Q(n16780) );
  AND2X1 U18234 ( .IN1(n16783), .IN2(n6803), .Q(n16782) );
  AND2X1 U18235 ( .IN1(n16785), .IN2(n6932), .Q(n16784) );
  AND2X1 U18236 ( .IN1(n16787), .IN2(n6943), .Q(n16786) );
  AND2X1 U18237 ( .IN1(P2_N3158), .IN2(n6834), .Q(n16788) );
  AND2X1 U18238 ( .IN1(P2_N3904), .IN2(n7484), .Q(n16789) );
  AND2X1 U18239 ( .IN1(P2_N3531), .IN2(n6834), .Q(n16790) );
  AND2X1 U18240 ( .IN1(P2_N4306), .IN2(n7484), .Q(n16791) );
  AND2X1 U18241 ( .IN1(n16793), .IN2(n6804), .Q(n16792) );
  AND2X1 U18242 ( .IN1(n16795), .IN2(n6803), .Q(n16794) );
  AND2X1 U18243 ( .IN1(P2_N4527), .IN2(n6943), .Q(n16796) );
  AND2X1 U18244 ( .IN1(n16798), .IN2(n6932), .Q(n16797) );
  AND2X1 U18245 ( .IN1(n16799), .IN2(n6970), .Q(n14642) );
  AND2X1 U18246 ( .IN1(n16800), .IN2(n6967), .Q(n14643) );
  AND2X1 U18247 ( .IN1(P2_N659), .IN2(n6834), .Q(n16801) );
  AND2X1 U18248 ( .IN1(P2_N1005), .IN2(n7484), .Q(n16802) );
  AND2X1 U18249 ( .IN1(P2_N393), .IN2(n6820), .Q(n16803) );
  AND2X1 U18250 ( .IN1(P2_N1260), .IN2(n7484), .Q(n16804) );
  AND2X1 U18251 ( .IN1(n16806), .IN2(n6804), .Q(n16805) );
  AND2X1 U18252 ( .IN1(n16808), .IN2(n6803), .Q(n16807) );
  AND2X1 U18253 ( .IN1(P2_N1667), .IN2(n6834), .Q(n16809) );
  AND2X1 U18254 ( .IN1(P2_N2413), .IN2(n7484), .Q(n16810) );
  AND2X1 U18255 ( .IN1(P2_N2040), .IN2(n6808), .Q(n16811) );
  AND2X1 U18256 ( .IN1(P2_N2786), .IN2(n7484), .Q(n16812) );
  AND2X1 U18257 ( .IN1(n16814), .IN2(n6804), .Q(n16813) );
  AND2X1 U18072 ( .IN1(P2_N4299), .IN2(n6825), .Q(n16560) );
  AND2X1 U18073 ( .IN1(n16562), .IN2(n6802), .Q(n16561) );
  AND2X1 U18074 ( .IN1(n16564), .IN2(P2_N291), .Q(n16563) );
  AND2X1 U18075 ( .IN1(P2_N4520), .IN2(n7460), .Q(n16565) );
  AND2X1 U18076 ( .IN1(n16567), .IN2(n6934), .Q(n16566) );
  AND2X1 U18077 ( .IN1(n16568), .IN2(n6966), .Q(n14628) );
  AND2X1 U18078 ( .IN1(n16569), .IN2(P2_N294), .Q(n14629) );
  AND2X1 U18079 ( .IN1(P2_N652), .IN2(n6828), .Q(n16570) );
  AND2X1 U18080 ( .IN1(P2_N998), .IN2(n6827), .Q(n16571) );
  AND2X1 U18081 ( .IN1(P2_N386), .IN2(n6828), .Q(n16572) );
  AND2X1 U18082 ( .IN1(P2_N1253), .IN2(n6827), .Q(n16573) );
  AND2X1 U18083 ( .IN1(n16575), .IN2(n6802), .Q(n16574) );
  AND2X1 U18084 ( .IN1(n16577), .IN2(P2_N291), .Q(n16576) );
  AND2X1 U18085 ( .IN1(P2_N1660), .IN2(n6822), .Q(n16578) );
  AND2X1 U18086 ( .IN1(P2_N2406), .IN2(n7486), .Q(n16579) );
  AND2X1 U18087 ( .IN1(P2_N2033), .IN2(n6822), .Q(n16580) );
  AND2X1 U18088 ( .IN1(P2_N2779), .IN2(n6825), .Q(n16581) );
  AND2X1 U18089 ( .IN1(n16583), .IN2(n6802), .Q(n16582) );
  AND2X1 U18090 ( .IN1(n16585), .IN2(P2_N291), .Q(n16584) );
  AND2X1 U18091 ( .IN1(n16587), .IN2(n6934), .Q(n16586) );
  AND2X1 U18092 ( .IN1(n16589), .IN2(n7460), .Q(n16588) );
  AND2X1 U18093 ( .IN1(P2_N3152), .IN2(n6822), .Q(n16590) );
  AND2X1 U18094 ( .IN1(P2_N3898), .IN2(n7486), .Q(n16591) );
  AND2X1 U18095 ( .IN1(P2_N3525), .IN2(n6816), .Q(n16592) );
  AND2X1 U18096 ( .IN1(P2_N4300), .IN2(n7486), .Q(n16593) );
  AND2X1 U18097 ( .IN1(n16595), .IN2(n6794), .Q(n16594) );
  AND2X1 U18098 ( .IN1(n16597), .IN2(n6793), .Q(n16596) );
  AND2X1 U18099 ( .IN1(P2_N4521), .IN2(n7460), .Q(n16598) );
  AND2X1 U18100 ( .IN1(n16600), .IN2(n6934), .Q(n16599) );
  AND2X1 U18101 ( .IN1(n16601), .IN2(n6966), .Q(n14630) );
  AND2X1 U18102 ( .IN1(n16602), .IN2(P2_N294), .Q(n14631) );
  AND2X1 U18103 ( .IN1(P2_N653), .IN2(n6828), .Q(n16603) );
  AND2X1 U18104 ( .IN1(P2_N999), .IN2(n6827), .Q(n16604) );
  AND2X1 U18105 ( .IN1(P2_N387), .IN2(n6828), .Q(n16605) );
  AND2X1 U18106 ( .IN1(P2_N1254), .IN2(n6827), .Q(n16606) );
  AND2X1 U18107 ( .IN1(n16608), .IN2(n6802), .Q(n16607) );
  AND2X1 U18108 ( .IN1(n16610), .IN2(P2_N291), .Q(n16609) );
  AND2X1 U18109 ( .IN1(P2_N1661), .IN2(n6816), .Q(n16611) );
  AND2X1 U18110 ( .IN1(P2_N2407), .IN2(n6825), .Q(n16612) );
  AND2X1 U18111 ( .IN1(P2_N2034), .IN2(n6816), .Q(n16613) );
  AND2X1 U18112 ( .IN1(P2_N2780), .IN2(n6825), .Q(n16614) );
  AND2X1 U18113 ( .IN1(n16616), .IN2(n6794), .Q(n16615) );
  AND2X1 U18114 ( .IN1(n16618), .IN2(n6793), .Q(n16617) );
  AND2X1 U18115 ( .IN1(n16620), .IN2(n6934), .Q(n16619) );
  AND2X1 U18116 ( .IN1(n16622), .IN2(n7460), .Q(n16621) );
  AND2X1 U18117 ( .IN1(P2_N3153), .IN2(n6822), .Q(n16623) );
  AND2X1 U18118 ( .IN1(P2_N3899), .IN2(n7486), .Q(n16624) );
  AND2X1 U18119 ( .IN1(P2_N3526), .IN2(n6830), .Q(n16625) );
  AND2X1 U18120 ( .IN1(P2_N4301), .IN2(n6829), .Q(n16626) );
  AND2X1 U18121 ( .IN1(n16628), .IN2(n6794), .Q(n16627) );
  AND2X1 U18122 ( .IN1(n16630), .IN2(n6793), .Q(n16629) );
  AND2X1 U18123 ( .IN1(P2_N4522), .IN2(n7460), .Q(n16631) );
  AND2X1 U18124 ( .IN1(n16633), .IN2(n6934), .Q(n16632) );
  AND2X1 U18125 ( .IN1(n16634), .IN2(n6966), .Q(n14632) );
  AND2X1 U18126 ( .IN1(n16635), .IN2(P2_N294), .Q(n14633) );
  AND2X1 U18127 ( .IN1(P2_N654), .IN2(n6828), .Q(n16636) );
  AND2X1 U18128 ( .IN1(P2_N1000), .IN2(n6827), .Q(n16637) );
  AND2X1 U18129 ( .IN1(P2_N388), .IN2(n6812), .Q(n16638) );
  AND2X1 U18130 ( .IN1(P2_N1255), .IN2(n7486), .Q(n16639) );
  AND2X1 U18131 ( .IN1(n16641), .IN2(n6802), .Q(n16640) );
  AND2X1 U18132 ( .IN1(n16643), .IN2(n6781), .Q(n16642) );
  AND2X1 U18133 ( .IN1(P2_N1662), .IN2(n6830), .Q(n16644) );
  AND2X1 U18134 ( .IN1(P2_N2408), .IN2(n6829), .Q(n16645) );
  AND2X1 U18135 ( .IN1(P2_N2035), .IN2(n6830), .Q(n16646) );
  AND2X1 U18136 ( .IN1(P2_N2781), .IN2(n6829), .Q(n16647) );
  AND2X1 U18137 ( .IN1(n16649), .IN2(n6794), .Q(n16648) );
  AND2X1 U18138 ( .IN1(n16651), .IN2(n6793), .Q(n16650) );
  AND2X1 U18139 ( .IN1(n16653), .IN2(n6934), .Q(n16652) );
  AND2X1 U18140 ( .IN1(n16655), .IN2(n7460), .Q(n16654) );
  AND2X1 U18141 ( .IN1(P2_N3154), .IN2(n6830), .Q(n16656) );
  AND2X1 U18142 ( .IN1(P2_N3900), .IN2(n6829), .Q(n16657) );
  AND2X1 U18143 ( .IN1(P2_N3527), .IN2(n6830), .Q(n16658) );
  AND2X1 U18144 ( .IN1(P2_N4302), .IN2(n6829), .Q(n16659) );
  AND2X1 U18145 ( .IN1(n16661), .IN2(n6794), .Q(n16660) );
  AND2X1 U18146 ( .IN1(n16663), .IN2(n6793), .Q(n16662) );
  AND2X1 U18147 ( .IN1(P2_N4523), .IN2(n6943), .Q(n16664) );
  AND2X1 U18148 ( .IN1(n16666), .IN2(n6934), .Q(n16665) );
  AND2X1 U18149 ( .IN1(n16667), .IN2(n6966), .Q(n14634) );
  AND2X1 U18150 ( .IN1(n16668), .IN2(P2_N294), .Q(n14635) );
  AND2X1 U18151 ( .IN1(P2_N655), .IN2(n6812), .Q(n16669) );
  AND2X1 U18152 ( .IN1(P2_N1001), .IN2(n7486), .Q(n16670) );
  AND2X1 U18153 ( .IN1(P2_N389), .IN2(n6812), .Q(n16671) );
  AND2X1 U18154 ( .IN1(P2_N1256), .IN2(n7486), .Q(n16672) );
  AND2X1 U18155 ( .IN1(n16674), .IN2(n6782), .Q(n16673) );
  AND2X1 U18156 ( .IN1(n16676), .IN2(n6781), .Q(n16675) );
  AND2X1 U18157 ( .IN1(P2_N1663), .IN2(n6830), .Q(n16677) );
  AND2X1 U18158 ( .IN1(P2_N2409), .IN2(n6829), .Q(n16678) );
  AND2X1 U18159 ( .IN1(P2_N2036), .IN2(n6830), .Q(n16679) );
  AND2X1 U18160 ( .IN1(P2_N2782), .IN2(n6829), .Q(n16680) );
  AND2X1 U18161 ( .IN1(n16682), .IN2(n6794), .Q(n16681) );
  AND2X1 U18162 ( .IN1(n16684), .IN2(n6793), .Q(n16683) );
  AND2X1 U18163 ( .IN1(n16686), .IN2(n6934), .Q(n16685) );
  AND2X1 U18164 ( .IN1(n16688), .IN2(n7460), .Q(n16687) );
  AND2X1 U17979 ( .IN1(P2_N4516), .IN2(n6937), .Q(n16433) );
  AND2X1 U17980 ( .IN1(n16435), .IN2(n6946), .Q(n16434) );
  AND2X1 U17981 ( .IN1(n16436), .IN2(n6970), .Q(n14620) );
  AND2X1 U17982 ( .IN1(n16437), .IN2(n6969), .Q(n14621) );
  AND2X1 U17983 ( .IN1(P2_N648), .IN2(n6820), .Q(n16438) );
  AND2X1 U17984 ( .IN1(P2_N994), .IN2(n6819), .Q(n16439) );
  AND2X1 U17985 ( .IN1(P2_N382), .IN2(n6820), .Q(n16440) );
  AND2X1 U17986 ( .IN1(P2_N1249), .IN2(n6813), .Q(n16441) );
  AND2X1 U17987 ( .IN1(n16443), .IN2(n6784), .Q(n16442) );
  AND2X1 U17988 ( .IN1(n16445), .IN2(n7488), .Q(n16444) );
  AND2X1 U17989 ( .IN1(P2_N1656), .IN2(n6842), .Q(n16446) );
  AND2X1 U17990 ( .IN1(P2_N2402), .IN2(n6827), .Q(n16447) );
  AND2X1 U17991 ( .IN1(P2_N2029), .IN2(n6842), .Q(n16448) );
  AND2X1 U17992 ( .IN1(P2_N2775), .IN2(n6827), .Q(n16449) );
  AND2X1 U17993 ( .IN1(n16451), .IN2(n6784), .Q(n16450) );
  AND2X1 U17994 ( .IN1(n16453), .IN2(n7488), .Q(n16452) );
  AND2X1 U17995 ( .IN1(n16455), .IN2(n6940), .Q(n16454) );
  AND2X1 U17996 ( .IN1(n16457), .IN2(n6931), .Q(n16456) );
  AND2X1 U17997 ( .IN1(P2_N3148), .IN2(n6842), .Q(n16458) );
  AND2X1 U17998 ( .IN1(P2_N3894), .IN2(n6827), .Q(n16459) );
  AND2X1 U17999 ( .IN1(P2_N3521), .IN2(n6842), .Q(n16460) );
  AND2X1 U18000 ( .IN1(P2_N4296), .IN2(n6819), .Q(n16461) );
  AND2X1 U18001 ( .IN1(n16463), .IN2(n6784), .Q(n16462) );
  AND2X1 U18002 ( .IN1(n16465), .IN2(n7488), .Q(n16464) );
  AND2X1 U18003 ( .IN1(P2_N4517), .IN2(n6931), .Q(n16466) );
  AND2X1 U18004 ( .IN1(n16468), .IN2(n6940), .Q(n16467) );
  AND2X1 U18005 ( .IN1(n16469), .IN2(n6970), .Q(n14622) );
  AND2X1 U18006 ( .IN1(n16470), .IN2(n6969), .Q(n14623) );
  AND2X1 U18007 ( .IN1(P2_N649), .IN2(n6820), .Q(n16471) );
  AND2X1 U18008 ( .IN1(P2_N995), .IN2(n6813), .Q(n16472) );
  AND2X1 U18009 ( .IN1(P2_N383), .IN2(n6828), .Q(n16473) );
  AND2X1 U18010 ( .IN1(P2_N1250), .IN2(n6813), .Q(n16474) );
  AND2X1 U18011 ( .IN1(n16476), .IN2(n6784), .Q(n16475) );
  AND2X1 U18012 ( .IN1(n16478), .IN2(n7488), .Q(n16477) );
  AND2X1 U18013 ( .IN1(P2_N1657), .IN2(n6842), .Q(n16479) );
  AND2X1 U18014 ( .IN1(P2_N2403), .IN2(n6819), .Q(n16480) );
  AND2X1 U18015 ( .IN1(P2_N2030), .IN2(n6842), .Q(n16481) );
  AND2X1 U18016 ( .IN1(P2_N2776), .IN2(n6827), .Q(n16482) );
  AND2X1 U18017 ( .IN1(n16484), .IN2(n6784), .Q(n16483) );
  AND2X1 U18018 ( .IN1(n16486), .IN2(n7488), .Q(n16485) );
  AND2X1 U18019 ( .IN1(n16488), .IN2(n6940), .Q(n16487) );
  AND2X1 U18020 ( .IN1(n16490), .IN2(n6943), .Q(n16489) );
  AND2X1 U18021 ( .IN1(P2_N3149), .IN2(n6842), .Q(n16491) );
  AND2X1 U18022 ( .IN1(P2_N3895), .IN2(n6819), .Q(n16492) );
  AND2X1 U18023 ( .IN1(P2_N3522), .IN2(n6842), .Q(n16493) );
  AND2X1 U18024 ( .IN1(P2_N4297), .IN2(n6819), .Q(n16494) );
  AND2X1 U18025 ( .IN1(n16496), .IN2(n6784), .Q(n16495) );
  AND2X1 U18026 ( .IN1(n16498), .IN2(n7488), .Q(n16497) );
  AND2X1 U18027 ( .IN1(P2_N4518), .IN2(n6931), .Q(n16499) );
  AND2X1 U18028 ( .IN1(n16501), .IN2(n6940), .Q(n16500) );
  AND2X1 U18029 ( .IN1(n16502), .IN2(n6970), .Q(n14624) );
  AND2X1 U18030 ( .IN1(n16503), .IN2(n6969), .Q(n14625) );
  AND2X1 U18031 ( .IN1(P2_N650), .IN2(n6828), .Q(n16504) );
  AND2X1 U18032 ( .IN1(P2_N996), .IN2(n6813), .Q(n16505) );
  AND2X1 U18033 ( .IN1(P2_N384), .IN2(n6828), .Q(n16506) );
  AND2X1 U18034 ( .IN1(P2_N1251), .IN2(n6813), .Q(n16507) );
  AND2X1 U18035 ( .IN1(n16509), .IN2(n6784), .Q(n16508) );
  AND2X1 U18036 ( .IN1(n16511), .IN2(n6793), .Q(n16510) );
  AND2X1 U18037 ( .IN1(P2_N1658), .IN2(n6842), .Q(n16512) );
  AND2X1 U18038 ( .IN1(P2_N2404), .IN2(n6827), .Q(n16513) );
  AND2X1 U18039 ( .IN1(P2_N2031), .IN2(n6842), .Q(n16514) );
  AND2X1 U18040 ( .IN1(P2_N2777), .IN2(n6827), .Q(n16515) );
  AND2X1 U18041 ( .IN1(n16517), .IN2(n6784), .Q(n16516) );
  AND2X1 U18042 ( .IN1(n16519), .IN2(n6793), .Q(n16518) );
  AND2X1 U18043 ( .IN1(n16521), .IN2(n6940), .Q(n16520) );
  AND2X1 U18044 ( .IN1(n16523), .IN2(n6931), .Q(n16522) );
  AND2X1 U18045 ( .IN1(P2_N3150), .IN2(n6842), .Q(n16524) );
  AND2X1 U18046 ( .IN1(P2_N3896), .IN2(n6827), .Q(n16525) );
  AND2X1 U18047 ( .IN1(P2_N3523), .IN2(n6842), .Q(n16526) );
  AND2X1 U18048 ( .IN1(P2_N4298), .IN2(n6827), .Q(n16527) );
  AND2X1 U18049 ( .IN1(n16529), .IN2(n6784), .Q(n16528) );
  AND2X1 U18050 ( .IN1(n16531), .IN2(n7488), .Q(n16530) );
  AND2X1 U18051 ( .IN1(P2_N4519), .IN2(n6931), .Q(n16532) );
  AND2X1 U18052 ( .IN1(n16534), .IN2(n6940), .Q(n16533) );
  AND2X1 U18053 ( .IN1(n16535), .IN2(n6972), .Q(n14626) );
  AND2X1 U18054 ( .IN1(n16536), .IN2(n6963), .Q(n14627) );
  AND2X1 U18055 ( .IN1(P2_N651), .IN2(n6828), .Q(n16537) );
  AND2X1 U18056 ( .IN1(P2_N997), .IN2(n6813), .Q(n16538) );
  AND2X1 U18057 ( .IN1(P2_N385), .IN2(n6828), .Q(n16539) );
  AND2X1 U18058 ( .IN1(P2_N1252), .IN2(n6813), .Q(n16540) );
  AND2X1 U18059 ( .IN1(n16542), .IN2(n6784), .Q(n16541) );
  AND2X1 U18060 ( .IN1(n16544), .IN2(n7488), .Q(n16543) );
  AND2X1 U18061 ( .IN1(P2_N1659), .IN2(n6828), .Q(n16545) );
  AND2X1 U18062 ( .IN1(P2_N2405), .IN2(n6827), .Q(n16546) );
  AND2X1 U18063 ( .IN1(P2_N2032), .IN2(n6830), .Q(n16547) );
  AND2X1 U18064 ( .IN1(P2_N2778), .IN2(n6825), .Q(n16548) );
  AND2X1 U18065 ( .IN1(n16550), .IN2(n6802), .Q(n16549) );
  AND2X1 U18066 ( .IN1(n16552), .IN2(P2_N291), .Q(n16551) );
  AND2X1 U18067 ( .IN1(n16554), .IN2(n6934), .Q(n16553) );
  AND2X1 U18068 ( .IN1(n16556), .IN2(n7460), .Q(n16555) );
  AND2X1 U18069 ( .IN1(P2_N3151), .IN2(n6816), .Q(n16557) );
  AND2X1 U18070 ( .IN1(P2_N3897), .IN2(n7486), .Q(n16558) );
  AND2X1 U18071 ( .IN1(P2_N3524), .IN2(n6822), .Q(n16559) );
  AND2X1 U17886 ( .IN1(n16305), .IN2(n6967), .Q(n14613) );
  AND2X1 U17887 ( .IN1(P2_N644), .IN2(n6822), .Q(n16306) );
  AND2X1 U17888 ( .IN1(P2_N990), .IN2(n6825), .Q(n16307) );
  AND2X1 U17889 ( .IN1(P2_N378), .IN2(n6822), .Q(n16308) );
  AND2X1 U17890 ( .IN1(P2_N1245), .IN2(n6825), .Q(n16309) );
  AND2X1 U17891 ( .IN1(n16311), .IN2(n6790), .Q(n16310) );
  AND2X1 U17892 ( .IN1(n16313), .IN2(n6789), .Q(n16312) );
  AND2X1 U17893 ( .IN1(P2_N1652), .IN2(n6816), .Q(n16314) );
  AND2X1 U17894 ( .IN1(P2_N2398), .IN2(n6825), .Q(n16315) );
  AND2X1 U17895 ( .IN1(P2_N2025), .IN2(n6812), .Q(n16316) );
  AND2X1 U17896 ( .IN1(P2_N2771), .IN2(n6825), .Q(n16317) );
  AND2X1 U17897 ( .IN1(n16319), .IN2(n6786), .Q(n16318) );
  AND2X1 U17898 ( .IN1(n16321), .IN2(n6789), .Q(n16320) );
  AND2X1 U17899 ( .IN1(n16323), .IN2(n6942), .Q(n16322) );
  AND2X1 U17900 ( .IN1(n16325), .IN2(n6937), .Q(n16324) );
  AND2X1 U17901 ( .IN1(P2_N3144), .IN2(n6816), .Q(n16326) );
  AND2X1 U17902 ( .IN1(P2_N3890), .IN2(n6825), .Q(n16327) );
  AND2X1 U17903 ( .IN1(P2_N3517), .IN2(n6816), .Q(n16328) );
  AND2X1 U17904 ( .IN1(P2_N4292), .IN2(n6825), .Q(n16329) );
  AND2X1 U17905 ( .IN1(n16331), .IN2(n6786), .Q(n16330) );
  AND2X1 U17906 ( .IN1(n16333), .IN2(n6789), .Q(n16332) );
  AND2X1 U17907 ( .IN1(P2_N4513), .IN2(n6937), .Q(n16334) );
  AND2X1 U17908 ( .IN1(n16336), .IN2(n6946), .Q(n16335) );
  AND2X1 U17909 ( .IN1(n16337), .IN2(n6970), .Q(n14614) );
  AND2X1 U17910 ( .IN1(n16338), .IN2(n6969), .Q(n14615) );
  AND2X1 U17911 ( .IN1(P2_N645), .IN2(n6822), .Q(n16339) );
  AND2X1 U17912 ( .IN1(P2_N991), .IN2(n7486), .Q(n16340) );
  AND2X1 U17913 ( .IN1(P2_N379), .IN2(n6822), .Q(n16341) );
  AND2X1 U17914 ( .IN1(P2_N1246), .IN2(n7486), .Q(n16342) );
  AND2X1 U17915 ( .IN1(n16344), .IN2(n6790), .Q(n16343) );
  AND2X1 U17916 ( .IN1(n16346), .IN2(n6789), .Q(n16345) );
  AND2X1 U17917 ( .IN1(P2_N1653), .IN2(n6822), .Q(n16347) );
  AND2X1 U17918 ( .IN1(P2_N2399), .IN2(n6825), .Q(n16348) );
  AND2X1 U17919 ( .IN1(P2_N2026), .IN2(n6822), .Q(n16349) );
  AND2X1 U17920 ( .IN1(P2_N2772), .IN2(n6825), .Q(n16350) );
  AND2X1 U17921 ( .IN1(n16352), .IN2(n6790), .Q(n16351) );
  AND2X1 U17922 ( .IN1(n16354), .IN2(n6789), .Q(n16353) );
  AND2X1 U17923 ( .IN1(n16356), .IN2(n6942), .Q(n16355) );
  AND2X1 U17924 ( .IN1(n16358), .IN2(n6937), .Q(n16357) );
  AND2X1 U17925 ( .IN1(P2_N3145), .IN2(n6822), .Q(n16359) );
  AND2X1 U17926 ( .IN1(P2_N3891), .IN2(n6825), .Q(n16360) );
  AND2X1 U17927 ( .IN1(P2_N3518), .IN2(n6822), .Q(n16361) );
  AND2X1 U17928 ( .IN1(P2_N4293), .IN2(n7486), .Q(n16362) );
  AND2X1 U17929 ( .IN1(n16364), .IN2(n6790), .Q(n16363) );
  AND2X1 U17930 ( .IN1(n16366), .IN2(n6789), .Q(n16365) );
  AND2X1 U17931 ( .IN1(P2_N4514), .IN2(n6937), .Q(n16367) );
  AND2X1 U17932 ( .IN1(n16369), .IN2(n6946), .Q(n16368) );
  AND2X1 U17933 ( .IN1(n16370), .IN2(n6970), .Q(n14616) );
  AND2X1 U17934 ( .IN1(n16371), .IN2(n6969), .Q(n14617) );
  AND2X1 U17935 ( .IN1(P2_N646), .IN2(n6820), .Q(n16372) );
  AND2X1 U17936 ( .IN1(P2_N992), .IN2(n6819), .Q(n16373) );
  AND2X1 U17937 ( .IN1(P2_N380), .IN2(n6820), .Q(n16374) );
  AND2X1 U17938 ( .IN1(P2_N1247), .IN2(n6819), .Q(n16375) );
  AND2X1 U17939 ( .IN1(n16377), .IN2(n6790), .Q(n16376) );
  AND2X1 U17940 ( .IN1(n16379), .IN2(n6789), .Q(n16378) );
  AND2X1 U17941 ( .IN1(P2_N1654), .IN2(n6822), .Q(n16380) );
  AND2X1 U17942 ( .IN1(P2_N2400), .IN2(n6825), .Q(n16381) );
  AND2X1 U17943 ( .IN1(P2_N2027), .IN2(n6822), .Q(n16382) );
  AND2X1 U17944 ( .IN1(P2_N2773), .IN2(n7486), .Q(n16383) );
  AND2X1 U17945 ( .IN1(n16385), .IN2(n6790), .Q(n16384) );
  AND2X1 U17946 ( .IN1(n16387), .IN2(n6789), .Q(n16386) );
  AND2X1 U17947 ( .IN1(n16389), .IN2(n6946), .Q(n16388) );
  AND2X1 U17948 ( .IN1(n16391), .IN2(n6937), .Q(n16390) );
  AND2X1 U17949 ( .IN1(P2_N3146), .IN2(n6820), .Q(n16392) );
  AND2X1 U17950 ( .IN1(P2_N3892), .IN2(n6819), .Q(n16393) );
  AND2X1 U17951 ( .IN1(P2_N3519), .IN2(n6820), .Q(n16394) );
  AND2X1 U17952 ( .IN1(P2_N4294), .IN2(n6819), .Q(n16395) );
  AND2X1 U17953 ( .IN1(n16397), .IN2(n6790), .Q(n16396) );
  AND2X1 U17954 ( .IN1(n16399), .IN2(n6789), .Q(n16398) );
  AND2X1 U17955 ( .IN1(P2_N4515), .IN2(n6937), .Q(n16400) );
  AND2X1 U17956 ( .IN1(n16402), .IN2(n6942), .Q(n16401) );
  AND2X1 U17957 ( .IN1(n16403), .IN2(n6970), .Q(n14618) );
  AND2X1 U17958 ( .IN1(n16404), .IN2(n6969), .Q(n14619) );
  AND2X1 U17959 ( .IN1(P2_N647), .IN2(n6820), .Q(n16405) );
  AND2X1 U17960 ( .IN1(P2_N993), .IN2(n6819), .Q(n16406) );
  AND2X1 U17961 ( .IN1(P2_N381), .IN2(n6820), .Q(n16407) );
  AND2X1 U17962 ( .IN1(P2_N1248), .IN2(n6819), .Q(n16408) );
  AND2X1 U17963 ( .IN1(n16410), .IN2(n6790), .Q(n16409) );
  AND2X1 U17964 ( .IN1(n16412), .IN2(n6789), .Q(n16411) );
  AND2X1 U17965 ( .IN1(P2_N1655), .IN2(n6820), .Q(n16413) );
  AND2X1 U17966 ( .IN1(P2_N2401), .IN2(n6819), .Q(n16414) );
  AND2X1 U17967 ( .IN1(P2_N2028), .IN2(n6820), .Q(n16415) );
  AND2X1 U17968 ( .IN1(P2_N2774), .IN2(n6819), .Q(n16416) );
  AND2X1 U17969 ( .IN1(n16418), .IN2(n6790), .Q(n16417) );
  AND2X1 U17970 ( .IN1(n16420), .IN2(n6789), .Q(n16419) );
  AND2X1 U17971 ( .IN1(n16422), .IN2(n6948), .Q(n16421) );
  AND2X1 U17972 ( .IN1(n16424), .IN2(n6937), .Q(n16423) );
  AND2X1 U17973 ( .IN1(P2_N3147), .IN2(n6820), .Q(n16425) );
  AND2X1 U17974 ( .IN1(P2_N3893), .IN2(n6819), .Q(n16426) );
  AND2X1 U17975 ( .IN1(P2_N3520), .IN2(n6820), .Q(n16427) );
  AND2X1 U17976 ( .IN1(P2_N4295), .IN2(n6819), .Q(n16428) );
  AND2X1 U17977 ( .IN1(n16430), .IN2(n6790), .Q(n16429) );
  AND2X1 U17978 ( .IN1(n16432), .IN2(n6789), .Q(n16431) );
  AND2X1 U17793 ( .IN1(P2_N374), .IN2(n6816), .Q(n16176) );
  AND2X1 U17794 ( .IN1(P2_N1241), .IN2(n6815), .Q(n16177) );
  AND2X1 U17795 ( .IN1(n16179), .IN2(n6786), .Q(n16178) );
  AND2X1 U17796 ( .IN1(n16181), .IN2(n6787), .Q(n16180) );
  AND2X1 U17797 ( .IN1(P2_N1648), .IN2(n6818), .Q(n16182) );
  AND2X1 U17798 ( .IN1(P2_N2394), .IN2(n6823), .Q(n16183) );
  AND2X1 U17799 ( .IN1(P2_N2021), .IN2(n6818), .Q(n16184) );
  AND2X1 U17800 ( .IN1(P2_N2767), .IN2(n6823), .Q(n16185) );
  AND2X1 U17801 ( .IN1(n16187), .IN2(n6776), .Q(n16186) );
  AND2X1 U17802 ( .IN1(n16189), .IN2(n6787), .Q(n16188) );
  AND2X1 U17803 ( .IN1(n16191), .IN2(n6948), .Q(n16190) );
  AND2X1 U17804 ( .IN1(n16193), .IN2(P2_N293), .Q(n16192) );
  AND2X1 U17805 ( .IN1(P2_N3140), .IN2(n6818), .Q(n16194) );
  AND2X1 U17806 ( .IN1(P2_N3886), .IN2(n6823), .Q(n16195) );
  AND2X1 U17807 ( .IN1(P2_N3513), .IN2(n6818), .Q(n16196) );
  AND2X1 U17808 ( .IN1(P2_N4288), .IN2(n6823), .Q(n16197) );
  AND2X1 U17809 ( .IN1(n16199), .IN2(n6786), .Q(n16198) );
  AND2X1 U17810 ( .IN1(n16201), .IN2(n6787), .Q(n16200) );
  AND2X1 U17811 ( .IN1(P2_N4509), .IN2(n6941), .Q(n16202) );
  AND2X1 U17812 ( .IN1(n16204), .IN2(n6948), .Q(n16203) );
  AND2X1 U17813 ( .IN1(n16205), .IN2(n6970), .Q(n14606) );
  AND2X1 U17814 ( .IN1(n16206), .IN2(n6963), .Q(n14607) );
  AND2X1 U17815 ( .IN1(P2_N641), .IN2(n6816), .Q(n16207) );
  AND2X1 U17816 ( .IN1(P2_N987), .IN2(n6815), .Q(n16208) );
  AND2X1 U17817 ( .IN1(P2_N375), .IN2(n6816), .Q(n16209) );
  AND2X1 U17818 ( .IN1(P2_N1242), .IN2(n6815), .Q(n16210) );
  AND2X1 U17819 ( .IN1(n16212), .IN2(n6786), .Q(n16211) );
  AND2X1 U17820 ( .IN1(n16214), .IN2(n6789), .Q(n16213) );
  AND2X1 U17821 ( .IN1(P2_N1649), .IN2(n6816), .Q(n16215) );
  AND2X1 U17822 ( .IN1(P2_N2395), .IN2(n6815), .Q(n16216) );
  AND2X1 U17823 ( .IN1(P2_N2022), .IN2(n6816), .Q(n16217) );
  AND2X1 U17824 ( .IN1(P2_N2768), .IN2(n6815), .Q(n16218) );
  AND2X1 U17825 ( .IN1(n16220), .IN2(n6786), .Q(n16219) );
  AND2X1 U17826 ( .IN1(n16222), .IN2(n6789), .Q(n16221) );
  AND2X1 U17827 ( .IN1(n16224), .IN2(n6946), .Q(n16223) );
  AND2X1 U17828 ( .IN1(n16226), .IN2(n6937), .Q(n16225) );
  AND2X1 U17829 ( .IN1(P2_N3141), .IN2(n6816), .Q(n16227) );
  AND2X1 U17830 ( .IN1(P2_N3887), .IN2(n6815), .Q(n16228) );
  AND2X1 U17831 ( .IN1(P2_N3514), .IN2(n6816), .Q(n16229) );
  AND2X1 U17832 ( .IN1(P2_N4289), .IN2(n6815), .Q(n16230) );
  AND2X1 U17833 ( .IN1(n16232), .IN2(n6786), .Q(n16231) );
  AND2X1 U17834 ( .IN1(n16234), .IN2(n6789), .Q(n16233) );
  AND2X1 U17835 ( .IN1(P2_N4510), .IN2(n6937), .Q(n16235) );
  AND2X1 U17836 ( .IN1(n16237), .IN2(n6946), .Q(n16236) );
  AND2X1 U17837 ( .IN1(n16238), .IN2(n6974), .Q(n14608) );
  AND2X1 U17838 ( .IN1(n16239), .IN2(n6967), .Q(n14609) );
  AND2X1 U17839 ( .IN1(P2_N642), .IN2(n6816), .Q(n16240) );
  AND2X1 U17840 ( .IN1(P2_N988), .IN2(n6815), .Q(n16241) );
  AND2X1 U17841 ( .IN1(P2_N376), .IN2(n6816), .Q(n16242) );
  AND2X1 U17842 ( .IN1(P2_N1243), .IN2(n6815), .Q(n16243) );
  AND2X1 U17843 ( .IN1(n16245), .IN2(n6786), .Q(n16244) );
  AND2X1 U17844 ( .IN1(n16247), .IN2(n6775), .Q(n16246) );
  AND2X1 U17845 ( .IN1(P2_N1650), .IN2(n6816), .Q(n16248) );
  AND2X1 U17846 ( .IN1(P2_N2396), .IN2(n6825), .Q(n16249) );
  AND2X1 U17847 ( .IN1(P2_N2023), .IN2(n6812), .Q(n16250) );
  AND2X1 U17848 ( .IN1(P2_N2769), .IN2(n6825), .Q(n16251) );
  AND2X1 U17849 ( .IN1(n16253), .IN2(n6786), .Q(n16252) );
  AND2X1 U17850 ( .IN1(n16255), .IN2(n6775), .Q(n16254) );
  AND2X1 U17851 ( .IN1(n16257), .IN2(n6946), .Q(n16256) );
  AND2X1 U17852 ( .IN1(n16259), .IN2(n6941), .Q(n16258) );
  AND2X1 U17853 ( .IN1(P2_N3142), .IN2(n6816), .Q(n16260) );
  AND2X1 U17854 ( .IN1(P2_N3888), .IN2(n6825), .Q(n16261) );
  AND2X1 U17855 ( .IN1(P2_N3515), .IN2(n6812), .Q(n16262) );
  AND2X1 U17856 ( .IN1(P2_N4290), .IN2(n6825), .Q(n16263) );
  AND2X1 U17857 ( .IN1(n16265), .IN2(n6786), .Q(n16264) );
  AND2X1 U17858 ( .IN1(n16267), .IN2(n6787), .Q(n16266) );
  AND2X1 U17859 ( .IN1(P2_N4511), .IN2(n6941), .Q(n16268) );
  AND2X1 U17860 ( .IN1(n16270), .IN2(n6946), .Q(n16269) );
  AND2X1 U17861 ( .IN1(n16271), .IN2(n6974), .Q(n14610) );
  AND2X1 U17862 ( .IN1(n16272), .IN2(n6967), .Q(n14611) );
  AND2X1 U17863 ( .IN1(P2_N643), .IN2(n6816), .Q(n16273) );
  AND2X1 U17864 ( .IN1(P2_N989), .IN2(n6815), .Q(n16274) );
  AND2X1 U17865 ( .IN1(P2_N377), .IN2(n6812), .Q(n16275) );
  AND2X1 U17866 ( .IN1(P2_N1244), .IN2(n6825), .Q(n16276) );
  AND2X1 U17867 ( .IN1(n16278), .IN2(n6786), .Q(n16277) );
  AND2X1 U17868 ( .IN1(n16280), .IN2(n6789), .Q(n16279) );
  AND2X1 U17869 ( .IN1(P2_N1651), .IN2(n6812), .Q(n16281) );
  AND2X1 U17870 ( .IN1(P2_N2397), .IN2(n6825), .Q(n16282) );
  AND2X1 U17871 ( .IN1(P2_N2024), .IN2(n6812), .Q(n16283) );
  AND2X1 U17872 ( .IN1(P2_N2770), .IN2(n6825), .Q(n16284) );
  AND2X1 U17873 ( .IN1(n16286), .IN2(n6786), .Q(n16285) );
  AND2X1 U17874 ( .IN1(n16288), .IN2(n6775), .Q(n16287) );
  AND2X1 U17875 ( .IN1(n16290), .IN2(n6946), .Q(n16289) );
  AND2X1 U17876 ( .IN1(n16292), .IN2(n6937), .Q(n16291) );
  AND2X1 U17877 ( .IN1(P2_N3143), .IN2(n6816), .Q(n16293) );
  AND2X1 U17878 ( .IN1(P2_N3889), .IN2(n6825), .Q(n16294) );
  AND2X1 U17879 ( .IN1(P2_N3516), .IN2(n6816), .Q(n16295) );
  AND2X1 U17880 ( .IN1(P2_N4291), .IN2(n6825), .Q(n16296) );
  AND2X1 U17881 ( .IN1(n16298), .IN2(n6786), .Q(n16297) );
  AND2X1 U17882 ( .IN1(n16300), .IN2(n6787), .Q(n16299) );
  AND2X1 U17883 ( .IN1(P2_N4512), .IN2(n6941), .Q(n16301) );
  AND2X1 U17884 ( .IN1(n16303), .IN2(n6946), .Q(n16302) );
  AND2X1 U17885 ( .IN1(n16304), .IN2(n6974), .Q(n14612) );
  AND2X1 U17700 ( .IN1(n16049), .IN2(n7487), .Q(n16048) );
  AND2X1 U17701 ( .IN1(P2_N1644), .IN2(n6824), .Q(n16050) );
  AND2X1 U17702 ( .IN1(P2_N2390), .IN2(n6823), .Q(n16051) );
  AND2X1 U17703 ( .IN1(P2_N2017), .IN2(n6824), .Q(n16052) );
  AND2X1 U17704 ( .IN1(P2_N2763), .IN2(n6823), .Q(n16053) );
  AND2X1 U17705 ( .IN1(n16055), .IN2(n6776), .Q(n16054) );
  AND2X1 U17706 ( .IN1(n16057), .IN2(n6787), .Q(n16056) );
  AND2X1 U17707 ( .IN1(n16059), .IN2(n6946), .Q(n16058) );
  AND2X1 U17708 ( .IN1(n16061), .IN2(P2_N293), .Q(n16060) );
  AND2X1 U17709 ( .IN1(P2_N3136), .IN2(n6852), .Q(n16062) );
  AND2X1 U17710 ( .IN1(P2_N3882), .IN2(n6851), .Q(n16063) );
  AND2X1 U17711 ( .IN1(P2_N3509), .IN2(n6824), .Q(n16064) );
  AND2X1 U17712 ( .IN1(P2_N4284), .IN2(n6823), .Q(n16065) );
  AND2X1 U17713 ( .IN1(n16067), .IN2(n6776), .Q(n16066) );
  AND2X1 U17714 ( .IN1(n16069), .IN2(n6775), .Q(n16068) );
  AND2X1 U17715 ( .IN1(P2_N4505), .IN2(P2_N293), .Q(n16070) );
  AND2X1 U17716 ( .IN1(n16072), .IN2(n6946), .Q(n16071) );
  AND2X1 U17717 ( .IN1(n16073), .IN2(n6970), .Q(n14598) );
  AND2X1 U17718 ( .IN1(n16074), .IN2(n6963), .Q(n14599) );
  AND2X1 U17719 ( .IN1(P2_N637), .IN2(n6852), .Q(n16075) );
  AND2X1 U17720 ( .IN1(P2_N983), .IN2(n6843), .Q(n16076) );
  AND2X1 U17721 ( .IN1(P2_N371), .IN2(n6824), .Q(n16077) );
  AND2X1 U17722 ( .IN1(P2_N1238), .IN2(n6843), .Q(n16078) );
  AND2X1 U17723 ( .IN1(n16080), .IN2(n6790), .Q(n16079) );
  AND2X1 U17724 ( .IN1(n16082), .IN2(n6787), .Q(n16081) );
  AND2X1 U17725 ( .IN1(P2_N1645), .IN2(n6824), .Q(n16083) );
  AND2X1 U17726 ( .IN1(P2_N2391), .IN2(n6823), .Q(n16084) );
  AND2X1 U17727 ( .IN1(P2_N2018), .IN2(n6824), .Q(n16085) );
  AND2X1 U17728 ( .IN1(P2_N2764), .IN2(n6823), .Q(n16086) );
  AND2X1 U17729 ( .IN1(n16088), .IN2(n6792), .Q(n16087) );
  AND2X1 U17730 ( .IN1(n16090), .IN2(n6787), .Q(n16089) );
  AND2X1 U17731 ( .IN1(n16092), .IN2(n6946), .Q(n16091) );
  AND2X1 U17732 ( .IN1(n16094), .IN2(P2_N293), .Q(n16093) );
  AND2X1 U17733 ( .IN1(P2_N3137), .IN2(n6824), .Q(n16095) );
  AND2X1 U17734 ( .IN1(P2_N3883), .IN2(n6823), .Q(n16096) );
  AND2X1 U17735 ( .IN1(P2_N3510), .IN2(n6824), .Q(n16097) );
  AND2X1 U17736 ( .IN1(P2_N4285), .IN2(n6823), .Q(n16098) );
  AND2X1 U17737 ( .IN1(n16100), .IN2(n6792), .Q(n16099) );
  AND2X1 U17738 ( .IN1(n16102), .IN2(n6787), .Q(n16101) );
  AND2X1 U17739 ( .IN1(P2_N4506), .IN2(P2_N293), .Q(n16103) );
  AND2X1 U17740 ( .IN1(n16105), .IN2(n6948), .Q(n16104) );
  AND2X1 U17741 ( .IN1(n16106), .IN2(n6970), .Q(n14600) );
  AND2X1 U17742 ( .IN1(n16107), .IN2(n6963), .Q(n14601) );
  AND2X1 U17743 ( .IN1(P2_N638), .IN2(n6852), .Q(n16108) );
  AND2X1 U17744 ( .IN1(P2_N984), .IN2(n6843), .Q(n16109) );
  AND2X1 U17745 ( .IN1(P2_N372), .IN2(n6836), .Q(n16110) );
  AND2X1 U17746 ( .IN1(P2_N1239), .IN2(n6843), .Q(n16111) );
  AND2X1 U17747 ( .IN1(n16113), .IN2(n6776), .Q(n16112) );
  AND2X1 U17748 ( .IN1(n16115), .IN2(n6787), .Q(n16114) );
  AND2X1 U17749 ( .IN1(P2_N1646), .IN2(n6824), .Q(n16116) );
  AND2X1 U17750 ( .IN1(P2_N2392), .IN2(n6823), .Q(n16117) );
  AND2X1 U17751 ( .IN1(P2_N2019), .IN2(n6824), .Q(n16118) );
  AND2X1 U17752 ( .IN1(P2_N2765), .IN2(n6823), .Q(n16119) );
  AND2X1 U17753 ( .IN1(n16121), .IN2(n6792), .Q(n16120) );
  AND2X1 U17754 ( .IN1(n16123), .IN2(n6775), .Q(n16122) );
  AND2X1 U17755 ( .IN1(n16125), .IN2(n6942), .Q(n16124) );
  AND2X1 U17756 ( .IN1(n16127), .IN2(P2_N293), .Q(n16126) );
  AND2X1 U17757 ( .IN1(P2_N3138), .IN2(n6824), .Q(n16128) );
  AND2X1 U17758 ( .IN1(P2_N3884), .IN2(n6823), .Q(n16129) );
  AND2X1 U17759 ( .IN1(P2_N3511), .IN2(n6824), .Q(n16130) );
  AND2X1 U17760 ( .IN1(P2_N4286), .IN2(n6823), .Q(n16131) );
  AND2X1 U17761 ( .IN1(n16133), .IN2(n6792), .Q(n16132) );
  AND2X1 U17762 ( .IN1(n16135), .IN2(n6775), .Q(n16134) );
  AND2X1 U17763 ( .IN1(P2_N4507), .IN2(P2_N293), .Q(n16136) );
  AND2X1 U17764 ( .IN1(n16138), .IN2(n6942), .Q(n16137) );
  AND2X1 U17765 ( .IN1(n16139), .IN2(n6974), .Q(n14602) );
  AND2X1 U17766 ( .IN1(n16140), .IN2(n6963), .Q(n14603) );
  AND2X1 U17767 ( .IN1(P2_N639), .IN2(n6836), .Q(n16141) );
  AND2X1 U17768 ( .IN1(P2_N985), .IN2(n6843), .Q(n16142) );
  AND2X1 U17769 ( .IN1(P2_N373), .IN2(n6836), .Q(n16143) );
  AND2X1 U17770 ( .IN1(P2_N1240), .IN2(n6843), .Q(n16144) );
  AND2X1 U17771 ( .IN1(n16146), .IN2(n6790), .Q(n16145) );
  AND2X1 U17772 ( .IN1(n16148), .IN2(n6787), .Q(n16147) );
  AND2X1 U17773 ( .IN1(P2_N1647), .IN2(n6824), .Q(n16149) );
  AND2X1 U17774 ( .IN1(P2_N2393), .IN2(n6823), .Q(n16150) );
  AND2X1 U17775 ( .IN1(P2_N2020), .IN2(n6824), .Q(n16151) );
  AND2X1 U17776 ( .IN1(P2_N2766), .IN2(n6823), .Q(n16152) );
  AND2X1 U17777 ( .IN1(n16154), .IN2(n6792), .Q(n16153) );
  AND2X1 U17778 ( .IN1(n16156), .IN2(n6787), .Q(n16155) );
  AND2X1 U17779 ( .IN1(n16158), .IN2(n6948), .Q(n16157) );
  AND2X1 U17780 ( .IN1(n16160), .IN2(P2_N293), .Q(n16159) );
  AND2X1 U17781 ( .IN1(P2_N3139), .IN2(n6824), .Q(n16161) );
  AND2X1 U17782 ( .IN1(P2_N3885), .IN2(n6823), .Q(n16162) );
  AND2X1 U17783 ( .IN1(P2_N3512), .IN2(n6824), .Q(n16163) );
  AND2X1 U17784 ( .IN1(P2_N4287), .IN2(n6823), .Q(n16164) );
  AND2X1 U17785 ( .IN1(n16166), .IN2(n6792), .Q(n16165) );
  AND2X1 U17786 ( .IN1(n16168), .IN2(n6775), .Q(n16167) );
  AND2X1 U17787 ( .IN1(P2_N4508), .IN2(P2_N293), .Q(n16169) );
  AND2X1 U17788 ( .IN1(n16171), .IN2(n6948), .Q(n16170) );
  AND2X1 U17789 ( .IN1(n16172), .IN2(n6974), .Q(n14604) );
  AND2X1 U17790 ( .IN1(n16173), .IN2(n6963), .Q(n14605) );
  AND2X1 U17791 ( .IN1(P2_N640), .IN2(n6818), .Q(n16174) );
  AND2X1 U17792 ( .IN1(P2_N986), .IN2(n6843), .Q(n16175) );
  AND2X1 U17607 ( .IN1(P2_N2013), .IN2(n6818), .Q(n15920) );
  AND2X1 U17608 ( .IN1(P2_N2759), .IN2(P2_N292), .Q(n15921) );
  AND2X1 U17609 ( .IN1(n15923), .IN2(n6790), .Q(n15922) );
  AND2X1 U17610 ( .IN1(n15925), .IN2(n6775), .Q(n15924) );
  AND2X1 U17611 ( .IN1(n15927), .IN2(n6942), .Q(n15926) );
  AND2X1 U17612 ( .IN1(n15929), .IN2(n6941), .Q(n15928) );
  AND2X1 U17613 ( .IN1(P2_N3132), .IN2(n6852), .Q(n15930) );
  AND2X1 U17614 ( .IN1(P2_N3878), .IN2(n6851), .Q(n15931) );
  AND2X1 U17615 ( .IN1(P2_N3505), .IN2(n6852), .Q(n15932) );
  AND2X1 U17616 ( .IN1(P2_N4280), .IN2(P2_N292), .Q(n15933) );
  AND2X1 U17617 ( .IN1(n15935), .IN2(n6786), .Q(n15934) );
  AND2X1 U17618 ( .IN1(n15937), .IN2(n7487), .Q(n15936) );
  AND2X1 U17619 ( .IN1(P2_N4501), .IN2(n6941), .Q(n15938) );
  AND2X1 U17620 ( .IN1(n15940), .IN2(n6942), .Q(n15939) );
  AND2X1 U17621 ( .IN1(n15941), .IN2(n6974), .Q(n14590) );
  AND2X1 U17622 ( .IN1(n15942), .IN2(n6967), .Q(n14591) );
  AND2X1 U17623 ( .IN1(P2_N633), .IN2(n6818), .Q(n15943) );
  AND2X1 U17624 ( .IN1(P2_N979), .IN2(P2_N292), .Q(n15944) );
  AND2X1 U17625 ( .IN1(n18813), .IN2(n6818), .Q(n15945) );
  AND2X1 U17626 ( .IN1(P2_N1234), .IN2(P2_N292), .Q(n15946) );
  AND2X1 U17627 ( .IN1(n15948), .IN2(n6776), .Q(n15947) );
  AND2X1 U17628 ( .IN1(n15950), .IN2(n6775), .Q(n15949) );
  AND2X1 U17629 ( .IN1(P2_N1641), .IN2(n6852), .Q(n15951) );
  AND2X1 U17630 ( .IN1(P2_N2387), .IN2(n6851), .Q(n15952) );
  AND2X1 U17631 ( .IN1(P2_N2014), .IN2(n6818), .Q(n15953) );
  AND2X1 U17632 ( .IN1(P2_N2760), .IN2(P2_N292), .Q(n15954) );
  AND2X1 U17633 ( .IN1(n15956), .IN2(n6776), .Q(n15955) );
  AND2X1 U17634 ( .IN1(n15958), .IN2(n7487), .Q(n15957) );
  AND2X1 U17635 ( .IN1(n15960), .IN2(n6942), .Q(n15959) );
  AND2X1 U17636 ( .IN1(n15962), .IN2(n6941), .Q(n15961) );
  AND2X1 U17637 ( .IN1(P2_N3133), .IN2(n6852), .Q(n15963) );
  AND2X1 U17638 ( .IN1(P2_N3879), .IN2(n6851), .Q(n15964) );
  AND2X1 U17639 ( .IN1(P2_N3506), .IN2(n6852), .Q(n15965) );
  AND2X1 U17640 ( .IN1(P2_N4281), .IN2(n6851), .Q(n15966) );
  AND2X1 U17641 ( .IN1(n15968), .IN2(n6792), .Q(n15967) );
  AND2X1 U17642 ( .IN1(n15970), .IN2(n7487), .Q(n15969) );
  AND2X1 U17643 ( .IN1(P2_N4502), .IN2(n6941), .Q(n15971) );
  AND2X1 U17644 ( .IN1(n15973), .IN2(n6942), .Q(n15972) );
  AND2X1 U17645 ( .IN1(n15974), .IN2(n6970), .Q(n14592) );
  AND2X1 U17646 ( .IN1(n15975), .IN2(n6963), .Q(n14593) );
  AND2X1 U17647 ( .IN1(P2_N634), .IN2(n6818), .Q(n15976) );
  AND2X1 U17648 ( .IN1(P2_N980), .IN2(P2_N292), .Q(n15977) );
  AND2X1 U17649 ( .IN1(P2_N368), .IN2(n6818), .Q(n15978) );
  AND2X1 U17650 ( .IN1(P2_N1235), .IN2(n6843), .Q(n15979) );
  AND2X1 U17651 ( .IN1(n15981), .IN2(n6790), .Q(n15980) );
  AND2X1 U17652 ( .IN1(n15983), .IN2(n7487), .Q(n15982) );
  AND2X1 U17653 ( .IN1(P2_N1642), .IN2(n6852), .Q(n15984) );
  AND2X1 U17654 ( .IN1(P2_N2388), .IN2(n6851), .Q(n15985) );
  AND2X1 U17655 ( .IN1(P2_N2015), .IN2(n6852), .Q(n15986) );
  AND2X1 U17656 ( .IN1(P2_N2761), .IN2(n6851), .Q(n15987) );
  AND2X1 U17657 ( .IN1(n15989), .IN2(n6792), .Q(n15988) );
  AND2X1 U17658 ( .IN1(n15991), .IN2(n7487), .Q(n15990) );
  AND2X1 U17659 ( .IN1(n15993), .IN2(n6942), .Q(n15992) );
  AND2X1 U17660 ( .IN1(n15995), .IN2(P2_N293), .Q(n15994) );
  AND2X1 U17661 ( .IN1(P2_N3134), .IN2(n6852), .Q(n15996) );
  AND2X1 U17662 ( .IN1(P2_N3880), .IN2(n6851), .Q(n15997) );
  AND2X1 U17663 ( .IN1(P2_N3507), .IN2(n6852), .Q(n15998) );
  AND2X1 U17664 ( .IN1(P2_N4282), .IN2(n6851), .Q(n15999) );
  AND2X1 U17665 ( .IN1(n16001), .IN2(n6792), .Q(n16000) );
  AND2X1 U17666 ( .IN1(n16003), .IN2(n7487), .Q(n16002) );
  AND2X1 U17667 ( .IN1(P2_N4503), .IN2(P2_N293), .Q(n16004) );
  AND2X1 U17668 ( .IN1(n16006), .IN2(n6946), .Q(n16005) );
  AND2X1 U17669 ( .IN1(n16007), .IN2(n6970), .Q(n14594) );
  AND2X1 U17670 ( .IN1(n16008), .IN2(n6963), .Q(n14595) );
  AND2X1 U17671 ( .IN1(P2_N635), .IN2(n6836), .Q(n16009) );
  AND2X1 U17672 ( .IN1(P2_N981), .IN2(n6843), .Q(n16010) );
  AND2X1 U17673 ( .IN1(P2_N369), .IN2(n6836), .Q(n16011) );
  AND2X1 U17674 ( .IN1(P2_N1236), .IN2(n6843), .Q(n16012) );
  AND2X1 U17675 ( .IN1(n16014), .IN2(n6786), .Q(n16013) );
  AND2X1 U17676 ( .IN1(n16016), .IN2(n7487), .Q(n16015) );
  AND2X1 U17677 ( .IN1(P2_N1643), .IN2(n6852), .Q(n16017) );
  AND2X1 U17678 ( .IN1(P2_N2389), .IN2(n6851), .Q(n16018) );
  AND2X1 U17679 ( .IN1(P2_N2016), .IN2(n6852), .Q(n16019) );
  AND2X1 U17680 ( .IN1(P2_N2762), .IN2(n6851), .Q(n16020) );
  AND2X1 U17681 ( .IN1(n16022), .IN2(n6792), .Q(n16021) );
  AND2X1 U17682 ( .IN1(n16024), .IN2(n7487), .Q(n16023) );
  AND2X1 U17683 ( .IN1(n16026), .IN2(n6942), .Q(n16025) );
  AND2X1 U17684 ( .IN1(n16028), .IN2(P2_N293), .Q(n16027) );
  AND2X1 U17685 ( .IN1(P2_N3135), .IN2(n6852), .Q(n16029) );
  AND2X1 U17686 ( .IN1(P2_N3881), .IN2(n6851), .Q(n16030) );
  AND2X1 U17687 ( .IN1(P2_N3508), .IN2(n6852), .Q(n16031) );
  AND2X1 U17688 ( .IN1(P2_N4283), .IN2(n6851), .Q(n16032) );
  AND2X1 U17689 ( .IN1(n16034), .IN2(n6792), .Q(n16033) );
  AND2X1 U17690 ( .IN1(n16036), .IN2(n7487), .Q(n16035) );
  AND2X1 U17691 ( .IN1(P2_N4504), .IN2(P2_N293), .Q(n16037) );
  AND2X1 U17692 ( .IN1(n16039), .IN2(n6946), .Q(n16038) );
  AND2X1 U17693 ( .IN1(n16040), .IN2(n6974), .Q(n14596) );
  AND2X1 U17694 ( .IN1(n16041), .IN2(n6963), .Q(n14597) );
  AND2X1 U17695 ( .IN1(P2_N636), .IN2(n6852), .Q(n16042) );
  AND2X1 U17696 ( .IN1(P2_N982), .IN2(n6843), .Q(n16043) );
  AND2X1 U17697 ( .IN1(P2_N370), .IN2(n6852), .Q(n16044) );
  AND2X1 U17698 ( .IN1(P2_N1237), .IN2(n6843), .Q(n16045) );
  AND2X1 U17699 ( .IN1(n16047), .IN2(n6792), .Q(n16046) );
  AND2X1 U17514 ( .IN1(P2_N4052), .IN2(n7485), .Q(n15793) );
  AND2X1 U17515 ( .IN1(P2_N3679), .IN2(n6820), .Q(n15794) );
  AND2X1 U17516 ( .IN1(P2_N4426), .IN2(n7485), .Q(n15795) );
  AND2X1 U17517 ( .IN1(n15797), .IN2(n6782), .Q(n15796) );
  AND2X1 U17518 ( .IN1(n15799), .IN2(n6781), .Q(n15798) );
  AND2X1 U17519 ( .IN1(P2_N391), .IN2(n14522), .Q(n15800) );
  AND2X1 U17520 ( .IN1(P2_N4689), .IN2(n6986), .Q(n15801) );
  AND2X1 U17521 ( .IN1(n15803), .IN2(n6932), .Q(n15802) );
  AND2X1 U17522 ( .IN1(n15805), .IN2(n6943), .Q(n15804) );
  AND2X1 U17523 ( .IN1(n15806), .IN2(n6966), .Q(n14582) );
  AND2X1 U17524 ( .IN1(n15807), .IN2(P2_N294), .Q(n14583) );
  AND2X1 U17525 ( .IN1(P2_N841), .IN2(n6820), .Q(n15808) );
  AND2X1 U17526 ( .IN1(P2_N1187), .IN2(n7485), .Q(n15809) );
  AND2X1 U17527 ( .IN1(P2_N913), .IN2(n6820), .Q(n15810) );
  AND2X1 U17528 ( .IN1(P2_N1442), .IN2(n7485), .Q(n15811) );
  AND2X1 U17529 ( .IN1(n15813), .IN2(n6782), .Q(n15812) );
  AND2X1 U17530 ( .IN1(n15815), .IN2(n6781), .Q(n15814) );
  AND2X1 U17531 ( .IN1(P2_N1815), .IN2(n6828), .Q(n15816) );
  AND2X1 U17532 ( .IN1(P2_N2561), .IN2(n7485), .Q(n15817) );
  AND2X1 U17533 ( .IN1(P2_N2188), .IN2(n6820), .Q(n15818) );
  AND2X1 U17534 ( .IN1(P2_N2934), .IN2(n7485), .Q(n15819) );
  AND2X1 U17535 ( .IN1(n15821), .IN2(n6782), .Q(n15820) );
  AND2X1 U17536 ( .IN1(n15823), .IN2(n6781), .Q(n15822) );
  AND2X1 U17537 ( .IN1(n15825), .IN2(n6932), .Q(n15824) );
  AND2X1 U17538 ( .IN1(n15827), .IN2(n6943), .Q(n15826) );
  AND2X1 U17539 ( .IN1(P2_N3307), .IN2(n6828), .Q(n15828) );
  AND2X1 U17540 ( .IN1(P2_N4053), .IN2(n7485), .Q(n15829) );
  AND2X1 U17541 ( .IN1(P2_N3680), .IN2(n6820), .Q(n15830) );
  AND2X1 U17542 ( .IN1(P2_N4427), .IN2(n7485), .Q(n15831) );
  AND2X1 U17543 ( .IN1(n15833), .IN2(n6782), .Q(n15832) );
  AND2X1 U17544 ( .IN1(n15835), .IN2(n6781), .Q(n15834) );
  AND2X1 U17545 ( .IN1(P2_N392), .IN2(n14522), .Q(n15836) );
  AND2X1 U17546 ( .IN1(P2_N4690), .IN2(n6986), .Q(n15837) );
  AND2X1 U17547 ( .IN1(n15839), .IN2(n6932), .Q(n15838) );
  AND2X1 U17548 ( .IN1(n15841), .IN2(n6943), .Q(n15840) );
  AND2X1 U17549 ( .IN1(n15842), .IN2(n6966), .Q(n14584) );
  AND2X1 U17550 ( .IN1(n15843), .IN2(P2_N294), .Q(n14585) );
  AND2X1 U17551 ( .IN1(P2_N630), .IN2(n6836), .Q(n15844) );
  AND2X1 U17552 ( .IN1(P2_N976), .IN2(n6835), .Q(n15845) );
  AND2X1 U17553 ( .IN1(n6681), .IN2(n6836), .Q(n15846) );
  AND2X1 U17554 ( .IN1(P2_N1231), .IN2(n6835), .Q(n15847) );
  AND2X1 U17555 ( .IN1(n15849), .IN2(n6776), .Q(n15848) );
  AND2X1 U17556 ( .IN1(n15851), .IN2(n6775), .Q(n15850) );
  AND2X1 U17557 ( .IN1(P2_N1638), .IN2(n6818), .Q(n15852) );
  AND2X1 U17558 ( .IN1(P2_N2384), .IN2(P2_N292), .Q(n15853) );
  AND2X1 U17559 ( .IN1(P2_N2011), .IN2(n6836), .Q(n15854) );
  AND2X1 U17560 ( .IN1(P2_N2757), .IN2(n6835), .Q(n15855) );
  AND2X1 U17561 ( .IN1(n15857), .IN2(n6776), .Q(n15856) );
  AND2X1 U17562 ( .IN1(n15859), .IN2(n6775), .Q(n15858) );
  AND2X1 U17563 ( .IN1(n15861), .IN2(n6946), .Q(n15860) );
  AND2X1 U17564 ( .IN1(n15863), .IN2(n6937), .Q(n15862) );
  AND2X1 U17565 ( .IN1(P2_N3130), .IN2(n6818), .Q(n15864) );
  AND2X1 U17566 ( .IN1(P2_N3876), .IN2(P2_N292), .Q(n15865) );
  AND2X1 U17567 ( .IN1(P2_N3503), .IN2(n6818), .Q(n15866) );
  AND2X1 U17568 ( .IN1(P2_N4278), .IN2(P2_N292), .Q(n15867) );
  AND2X1 U17569 ( .IN1(n15869), .IN2(n6776), .Q(n15868) );
  AND2X1 U17570 ( .IN1(n15871), .IN2(n6775), .Q(n15870) );
  AND2X1 U17571 ( .IN1(P2_N4499), .IN2(n6941), .Q(n15872) );
  AND2X1 U17572 ( .IN1(n15874), .IN2(n6942), .Q(n15873) );
  AND2X1 U17573 ( .IN1(n15875), .IN2(n6974), .Q(n14586) );
  AND2X1 U17574 ( .IN1(n15876), .IN2(n6967), .Q(n14587) );
  AND2X1 U17575 ( .IN1(P2_N631), .IN2(n6836), .Q(n15877) );
  AND2X1 U17576 ( .IN1(P2_N977), .IN2(n6835), .Q(n15878) );
  AND2X1 U17577 ( .IN1(n6682), .IN2(n6836), .Q(n15879) );
  AND2X1 U17578 ( .IN1(P2_N1232), .IN2(n6835), .Q(n15880) );
  AND2X1 U17579 ( .IN1(n15882), .IN2(n6776), .Q(n15881) );
  AND2X1 U17580 ( .IN1(n15884), .IN2(n6775), .Q(n15883) );
  AND2X1 U17581 ( .IN1(P2_N1639), .IN2(n6818), .Q(n15885) );
  AND2X1 U17582 ( .IN1(P2_N2385), .IN2(P2_N292), .Q(n15886) );
  AND2X1 U17583 ( .IN1(P2_N2012), .IN2(n6836), .Q(n15887) );
  AND2X1 U17584 ( .IN1(P2_N2758), .IN2(n6835), .Q(n15888) );
  AND2X1 U17585 ( .IN1(n15890), .IN2(n6776), .Q(n15889) );
  AND2X1 U17586 ( .IN1(n15892), .IN2(n6775), .Q(n15891) );
  AND2X1 U17587 ( .IN1(n15894), .IN2(n6942), .Q(n15893) );
  AND2X1 U17588 ( .IN1(n15896), .IN2(n6941), .Q(n15895) );
  AND2X1 U17589 ( .IN1(P2_N3131), .IN2(n6818), .Q(n15897) );
  AND2X1 U17590 ( .IN1(P2_N3877), .IN2(P2_N292), .Q(n15898) );
  AND2X1 U17591 ( .IN1(P2_N3504), .IN2(n6818), .Q(n15899) );
  AND2X1 U17592 ( .IN1(P2_N4279), .IN2(P2_N292), .Q(n15900) );
  AND2X1 U17593 ( .IN1(n15902), .IN2(n6776), .Q(n15901) );
  AND2X1 U17594 ( .IN1(n15904), .IN2(n6775), .Q(n15903) );
  AND2X1 U17595 ( .IN1(P2_N4500), .IN2(n6941), .Q(n15905) );
  AND2X1 U17596 ( .IN1(n15907), .IN2(n6942), .Q(n15906) );
  AND2X1 U17597 ( .IN1(n15908), .IN2(n6974), .Q(n14588) );
  AND2X1 U17598 ( .IN1(n15909), .IN2(n6967), .Q(n14589) );
  AND2X1 U17599 ( .IN1(P2_N632), .IN2(n6836), .Q(n15910) );
  AND2X1 U17600 ( .IN1(P2_N978), .IN2(n6835), .Q(n15911) );
  AND2X1 U17601 ( .IN1(n6683), .IN2(n6836), .Q(n15912) );
  AND2X1 U17602 ( .IN1(P2_N1233), .IN2(n6835), .Q(n15913) );
  AND2X1 U17603 ( .IN1(n15915), .IN2(n6776), .Q(n15914) );
  AND2X1 U17604 ( .IN1(n15917), .IN2(n6775), .Q(n15916) );
  AND2X1 U17605 ( .IN1(P2_N1640), .IN2(n6852), .Q(n15918) );
  AND2X1 U17606 ( .IN1(P2_N2386), .IN2(P2_N292), .Q(n15919) );
  AND2X1 U17421 ( .IN1(P2_N837), .IN2(n6828), .Q(n15664) );
  AND2X1 U17422 ( .IN1(P2_N1183), .IN2(n6827), .Q(n15665) );
  AND2X1 U17423 ( .IN1(P2_N909), .IN2(n6828), .Q(n15666) );
  AND2X1 U17424 ( .IN1(P2_N1438), .IN2(n6827), .Q(n15667) );
  AND2X1 U17425 ( .IN1(n15669), .IN2(n6802), .Q(n15668) );
  AND2X1 U17426 ( .IN1(n15671), .IN2(P2_N291), .Q(n15670) );
  AND2X1 U17427 ( .IN1(P2_N1811), .IN2(n6812), .Q(n15672) );
  AND2X1 U17428 ( .IN1(P2_N2557), .IN2(n7486), .Q(n15673) );
  AND2X1 U17429 ( .IN1(P2_N2184), .IN2(n6812), .Q(n15674) );
  AND2X1 U17430 ( .IN1(P2_N2930), .IN2(n7486), .Q(n15675) );
  AND2X1 U17431 ( .IN1(n15677), .IN2(n6802), .Q(n15676) );
  AND2X1 U17432 ( .IN1(n15679), .IN2(n6781), .Q(n15678) );
  AND2X1 U17433 ( .IN1(n15681), .IN2(n6934), .Q(n15680) );
  AND2X1 U17434 ( .IN1(n15683), .IN2(n7460), .Q(n15682) );
  AND2X1 U17435 ( .IN1(P2_N3303), .IN2(n6812), .Q(n15684) );
  AND2X1 U17436 ( .IN1(P2_N4049), .IN2(n7486), .Q(n15685) );
  AND2X1 U17437 ( .IN1(P2_N3676), .IN2(n6812), .Q(n15686) );
  AND2X1 U17438 ( .IN1(P2_N4423), .IN2(n7486), .Q(n15687) );
  AND2X1 U17439 ( .IN1(n15689), .IN2(n6782), .Q(n15688) );
  AND2X1 U17440 ( .IN1(n15691), .IN2(n6781), .Q(n15690) );
  AND2X1 U17441 ( .IN1(P2_N388), .IN2(n14522), .Q(n15692) );
  AND2X1 U17442 ( .IN1(P2_N4686), .IN2(n6986), .Q(n15693) );
  AND2X1 U17443 ( .IN1(n15695), .IN2(n6934), .Q(n15694) );
  AND2X1 U17444 ( .IN1(n15697), .IN2(n7460), .Q(n15696) );
  AND2X1 U17445 ( .IN1(n15698), .IN2(n6966), .Q(n14576) );
  AND2X1 U17446 ( .IN1(n15699), .IN2(P2_N294), .Q(n14577) );
  AND2X1 U17447 ( .IN1(P2_N838), .IN2(n6828), .Q(n15700) );
  AND2X1 U17448 ( .IN1(P2_N1184), .IN2(n7486), .Q(n15701) );
  AND2X1 U17449 ( .IN1(P2_N910), .IN2(n6828), .Q(n15702) );
  AND2X1 U17450 ( .IN1(P2_N1439), .IN2(n6827), .Q(n15703) );
  AND2X1 U17451 ( .IN1(n15705), .IN2(n6802), .Q(n15704) );
  AND2X1 U17452 ( .IN1(n15707), .IN2(P2_N291), .Q(n15706) );
  AND2X1 U17453 ( .IN1(P2_N1812), .IN2(n6812), .Q(n15708) );
  AND2X1 U17454 ( .IN1(P2_N2558), .IN2(n7486), .Q(n15709) );
  AND2X1 U17455 ( .IN1(P2_N2185), .IN2(n6812), .Q(n15710) );
  AND2X1 U17456 ( .IN1(P2_N2931), .IN2(n7486), .Q(n15711) );
  AND2X1 U17457 ( .IN1(n15713), .IN2(n6782), .Q(n15712) );
  AND2X1 U17458 ( .IN1(n15715), .IN2(n6781), .Q(n15714) );
  AND2X1 U17459 ( .IN1(n15717), .IN2(n6934), .Q(n15716) );
  AND2X1 U17460 ( .IN1(n15719), .IN2(n7460), .Q(n15718) );
  AND2X1 U17461 ( .IN1(P2_N3304), .IN2(n6812), .Q(n15720) );
  AND2X1 U17462 ( .IN1(P2_N4050), .IN2(n7486), .Q(n15721) );
  AND2X1 U17463 ( .IN1(P2_N3677), .IN2(n6812), .Q(n15722) );
  AND2X1 U17464 ( .IN1(P2_N4424), .IN2(n7486), .Q(n15723) );
  AND2X1 U17465 ( .IN1(n15725), .IN2(n6782), .Q(n15724) );
  AND2X1 U17466 ( .IN1(n15727), .IN2(n6781), .Q(n15726) );
  AND2X1 U17467 ( .IN1(P2_N389), .IN2(n14522), .Q(n15728) );
  AND2X1 U17468 ( .IN1(P2_N4687), .IN2(n6986), .Q(n15729) );
  AND2X1 U17469 ( .IN1(n15731), .IN2(n6934), .Q(n15730) );
  AND2X1 U17470 ( .IN1(n15733), .IN2(n7460), .Q(n15732) );
  AND2X1 U17471 ( .IN1(n15734), .IN2(n6966), .Q(n14578) );
  AND2X1 U17472 ( .IN1(n15735), .IN2(P2_N294), .Q(n14579) );
  AND2X1 U17473 ( .IN1(P2_N839), .IN2(n6828), .Q(n15736) );
  AND2X1 U17474 ( .IN1(P2_N1185), .IN2(n7485), .Q(n15737) );
  AND2X1 U17475 ( .IN1(P2_N911), .IN2(n6812), .Q(n15738) );
  AND2X1 U17476 ( .IN1(P2_N1440), .IN2(n7485), .Q(n15739) );
  AND2X1 U17477 ( .IN1(n15741), .IN2(n6782), .Q(n15740) );
  AND2X1 U17478 ( .IN1(n15743), .IN2(n6781), .Q(n15742) );
  AND2X1 U17479 ( .IN1(P2_N1813), .IN2(n6812), .Q(n15744) );
  AND2X1 U17480 ( .IN1(P2_N2559), .IN2(n7486), .Q(n15745) );
  AND2X1 U17481 ( .IN1(P2_N2186), .IN2(n6812), .Q(n15746) );
  AND2X1 U17482 ( .IN1(P2_N2932), .IN2(n7486), .Q(n15747) );
  AND2X1 U17483 ( .IN1(n15749), .IN2(n6782), .Q(n15748) );
  AND2X1 U17484 ( .IN1(n15751), .IN2(n6781), .Q(n15750) );
  AND2X1 U17485 ( .IN1(n15753), .IN2(n6934), .Q(n15752) );
  AND2X1 U17486 ( .IN1(n15755), .IN2(n7460), .Q(n15754) );
  AND2X1 U17487 ( .IN1(P2_N3305), .IN2(n6812), .Q(n15756) );
  AND2X1 U17488 ( .IN1(P2_N4051), .IN2(n7486), .Q(n15757) );
  AND2X1 U17489 ( .IN1(P2_N3678), .IN2(n6812), .Q(n15758) );
  AND2X1 U17490 ( .IN1(P2_N4425), .IN2(n7486), .Q(n15759) );
  AND2X1 U17491 ( .IN1(n15761), .IN2(n6782), .Q(n15760) );
  AND2X1 U17492 ( .IN1(n15763), .IN2(n6781), .Q(n15762) );
  AND2X1 U17493 ( .IN1(P2_N390), .IN2(n14522), .Q(n15764) );
  AND2X1 U17494 ( .IN1(P2_N4688), .IN2(n6986), .Q(n15765) );
  AND2X1 U17495 ( .IN1(n15767), .IN2(n6934), .Q(n15766) );
  AND2X1 U17496 ( .IN1(n15769), .IN2(n6943), .Q(n15768) );
  AND2X1 U17497 ( .IN1(n15770), .IN2(n6966), .Q(n14580) );
  AND2X1 U17498 ( .IN1(n15771), .IN2(P2_N294), .Q(n14581) );
  AND2X1 U17499 ( .IN1(P2_N840), .IN2(n6820), .Q(n15772) );
  AND2X1 U17500 ( .IN1(P2_N1186), .IN2(n7485), .Q(n15773) );
  AND2X1 U17501 ( .IN1(P2_N912), .IN2(n6828), .Q(n15774) );
  AND2X1 U17502 ( .IN1(P2_N1441), .IN2(n7485), .Q(n15775) );
  AND2X1 U17503 ( .IN1(n15777), .IN2(n6782), .Q(n15776) );
  AND2X1 U17504 ( .IN1(n15779), .IN2(n6781), .Q(n15778) );
  AND2X1 U17505 ( .IN1(P2_N1814), .IN2(n6812), .Q(n15780) );
  AND2X1 U17506 ( .IN1(P2_N2560), .IN2(n7485), .Q(n15781) );
  AND2X1 U17507 ( .IN1(P2_N2187), .IN2(n6828), .Q(n15782) );
  AND2X1 U17508 ( .IN1(P2_N2933), .IN2(n7485), .Q(n15783) );
  AND2X1 U17509 ( .IN1(n15785), .IN2(n6782), .Q(n15784) );
  AND2X1 U17510 ( .IN1(n15787), .IN2(n6781), .Q(n15786) );
  AND2X1 U17511 ( .IN1(n15789), .IN2(n6934), .Q(n15788) );
  AND2X1 U17512 ( .IN1(n15791), .IN2(n6943), .Q(n15790) );
  AND2X1 U17513 ( .IN1(P2_N3306), .IN2(n6820), .Q(n15792) );
  AND2X1 U17328 ( .IN1(n15535), .IN2(n6793), .Q(n15534) );
  AND2X1 U17329 ( .IN1(n15537), .IN2(n6940), .Q(n15536) );
  AND2X1 U17330 ( .IN1(n15539), .IN2(n6931), .Q(n15538) );
  AND2X1 U17331 ( .IN1(P2_N3299), .IN2(n6842), .Q(n15540) );
  AND2X1 U17332 ( .IN1(P2_N4045), .IN2(n6813), .Q(n15541) );
  AND2X1 U17333 ( .IN1(P2_N3672), .IN2(n6842), .Q(n15542) );
  AND2X1 U17334 ( .IN1(P2_N4419), .IN2(n6813), .Q(n15543) );
  AND2X1 U17335 ( .IN1(n15545), .IN2(n6784), .Q(n15544) );
  AND2X1 U17336 ( .IN1(n15547), .IN2(n7488), .Q(n15546) );
  AND2X1 U17337 ( .IN1(P2_N384), .IN2(n14522), .Q(n15548) );
  AND2X1 U17338 ( .IN1(P2_N4682), .IN2(n6986), .Q(n15549) );
  AND2X1 U17339 ( .IN1(n15551), .IN2(n6940), .Q(n15550) );
  AND2X1 U17340 ( .IN1(n15553), .IN2(n6931), .Q(n15552) );
  AND2X1 U17341 ( .IN1(n15554), .IN2(n6972), .Q(n14568) );
  AND2X1 U17342 ( .IN1(n15555), .IN2(n6963), .Q(n14569) );
  AND2X1 U17343 ( .IN1(P2_N834), .IN2(n6828), .Q(n15556) );
  AND2X1 U17344 ( .IN1(P2_N1180), .IN2(n6813), .Q(n15557) );
  AND2X1 U17345 ( .IN1(P2_N906), .IN2(n6828), .Q(n15558) );
  AND2X1 U17346 ( .IN1(P2_N1435), .IN2(n6813), .Q(n15559) );
  AND2X1 U17347 ( .IN1(n15561), .IN2(n6784), .Q(n15560) );
  AND2X1 U17348 ( .IN1(n15563), .IN2(n7488), .Q(n15562) );
  AND2X1 U17349 ( .IN1(P2_N1808), .IN2(n6828), .Q(n15564) );
  AND2X1 U17350 ( .IN1(P2_N2554), .IN2(n6827), .Q(n15565) );
  AND2X1 U17351 ( .IN1(P2_N2181), .IN2(n6828), .Q(n15566) );
  AND2X1 U17352 ( .IN1(P2_N2927), .IN2(n6827), .Q(n15567) );
  AND2X1 U17353 ( .IN1(n15569), .IN2(n6802), .Q(n15568) );
  AND2X1 U17354 ( .IN1(n15571), .IN2(P2_N291), .Q(n15570) );
  AND2X1 U17355 ( .IN1(n15573), .IN2(n6934), .Q(n15572) );
  AND2X1 U17356 ( .IN1(n15575), .IN2(n7460), .Q(n15574) );
  AND2X1 U17357 ( .IN1(P2_N3300), .IN2(n6828), .Q(n15576) );
  AND2X1 U17358 ( .IN1(P2_N4046), .IN2(n6827), .Q(n15577) );
  AND2X1 U17359 ( .IN1(P2_N3673), .IN2(n6828), .Q(n15578) );
  AND2X1 U17360 ( .IN1(P2_N4420), .IN2(n6827), .Q(n15579) );
  AND2X1 U17361 ( .IN1(n15581), .IN2(n6802), .Q(n15580) );
  AND2X1 U17362 ( .IN1(n15583), .IN2(P2_N291), .Q(n15582) );
  AND2X1 U17363 ( .IN1(P2_N385), .IN2(n14522), .Q(n15584) );
  AND2X1 U17364 ( .IN1(P2_N4683), .IN2(n6986), .Q(n15585) );
  AND2X1 U17365 ( .IN1(n15587), .IN2(n6934), .Q(n15586) );
  AND2X1 U17366 ( .IN1(n15589), .IN2(n7460), .Q(n15588) );
  AND2X1 U17367 ( .IN1(n15590), .IN2(n6966), .Q(n14570) );
  AND2X1 U17368 ( .IN1(n15591), .IN2(P2_N294), .Q(n14571) );
  AND2X1 U17369 ( .IN1(P2_N835), .IN2(n6828), .Q(n15592) );
  AND2X1 U17370 ( .IN1(P2_N1181), .IN2(n6827), .Q(n15593) );
  AND2X1 U17371 ( .IN1(P2_N907), .IN2(n6828), .Q(n15594) );
  AND2X1 U17372 ( .IN1(P2_N1436), .IN2(n6827), .Q(n15595) );
  AND2X1 U17373 ( .IN1(n15597), .IN2(n6802), .Q(n15596) );
  AND2X1 U17374 ( .IN1(n15599), .IN2(P2_N291), .Q(n15598) );
  AND2X1 U17375 ( .IN1(P2_N1809), .IN2(n6828), .Q(n15600) );
  AND2X1 U17376 ( .IN1(P2_N2555), .IN2(n6827), .Q(n15601) );
  AND2X1 U17377 ( .IN1(P2_N2182), .IN2(n6828), .Q(n15602) );
  AND2X1 U17378 ( .IN1(P2_N2928), .IN2(n6827), .Q(n15603) );
  AND2X1 U17379 ( .IN1(n15605), .IN2(n6802), .Q(n15604) );
  AND2X1 U17380 ( .IN1(n15607), .IN2(P2_N291), .Q(n15606) );
  AND2X1 U17381 ( .IN1(n15609), .IN2(n6934), .Q(n15608) );
  AND2X1 U17382 ( .IN1(n15611), .IN2(n7460), .Q(n15610) );
  AND2X1 U17383 ( .IN1(P2_N3301), .IN2(n6828), .Q(n15612) );
  AND2X1 U17384 ( .IN1(P2_N4047), .IN2(n6827), .Q(n15613) );
  AND2X1 U17385 ( .IN1(P2_N3674), .IN2(n6812), .Q(n15614) );
  AND2X1 U17386 ( .IN1(P2_N4421), .IN2(n6827), .Q(n15615) );
  AND2X1 U17387 ( .IN1(n15617), .IN2(n6802), .Q(n15616) );
  AND2X1 U17388 ( .IN1(n15619), .IN2(P2_N291), .Q(n15618) );
  AND2X1 U17389 ( .IN1(P2_N386), .IN2(n14522), .Q(n15620) );
  AND2X1 U17390 ( .IN1(P2_N4684), .IN2(n6986), .Q(n15621) );
  AND2X1 U17391 ( .IN1(n15623), .IN2(n6934), .Q(n15622) );
  AND2X1 U17392 ( .IN1(n15625), .IN2(n7460), .Q(n15624) );
  AND2X1 U17393 ( .IN1(n15626), .IN2(n6966), .Q(n14572) );
  AND2X1 U17394 ( .IN1(n15627), .IN2(P2_N294), .Q(n14573) );
  AND2X1 U17395 ( .IN1(P2_N836), .IN2(n6828), .Q(n15628) );
  AND2X1 U17396 ( .IN1(P2_N1182), .IN2(n6827), .Q(n15629) );
  AND2X1 U17397 ( .IN1(P2_N908), .IN2(n6828), .Q(n15630) );
  AND2X1 U17398 ( .IN1(P2_N1437), .IN2(n6827), .Q(n15631) );
  AND2X1 U17399 ( .IN1(n15633), .IN2(n6802), .Q(n15632) );
  AND2X1 U17400 ( .IN1(n15635), .IN2(P2_N291), .Q(n15634) );
  AND2X1 U17401 ( .IN1(P2_N1810), .IN2(n6812), .Q(n15636) );
  AND2X1 U17402 ( .IN1(P2_N2556), .IN2(n7486), .Q(n15637) );
  AND2X1 U17403 ( .IN1(P2_N2183), .IN2(n6812), .Q(n15638) );
  AND2X1 U17404 ( .IN1(P2_N2929), .IN2(n7486), .Q(n15639) );
  AND2X1 U17405 ( .IN1(n15641), .IN2(n6802), .Q(n15640) );
  AND2X1 U17406 ( .IN1(n15643), .IN2(n6781), .Q(n15642) );
  AND2X1 U17407 ( .IN1(n15645), .IN2(n6934), .Q(n15644) );
  AND2X1 U17408 ( .IN1(n15647), .IN2(n7460), .Q(n15646) );
  AND2X1 U17409 ( .IN1(P2_N3302), .IN2(n6812), .Q(n15648) );
  AND2X1 U17410 ( .IN1(P2_N4048), .IN2(n7486), .Q(n15649) );
  AND2X1 U17411 ( .IN1(P2_N3675), .IN2(n6812), .Q(n15650) );
  AND2X1 U17412 ( .IN1(P2_N4422), .IN2(n7486), .Q(n15651) );
  AND2X1 U17413 ( .IN1(n15653), .IN2(n6802), .Q(n15652) );
  AND2X1 U17414 ( .IN1(n15655), .IN2(n6781), .Q(n15654) );
  AND2X1 U17415 ( .IN1(P2_N387), .IN2(n14522), .Q(n15656) );
  AND2X1 U17416 ( .IN1(P2_N4685), .IN2(n6986), .Q(n15657) );
  AND2X1 U17417 ( .IN1(n15659), .IN2(n6934), .Q(n15658) );
  AND2X1 U17418 ( .IN1(n15661), .IN2(n7460), .Q(n15660) );
  AND2X1 U17419 ( .IN1(n15662), .IN2(n6966), .Q(n14574) );
  AND2X1 U17420 ( .IN1(n15663), .IN2(P2_N294), .Q(n14575) );
  AND2X1 U17235 ( .IN1(n15407), .IN2(n6946), .Q(n15406) );
  AND2X1 U17236 ( .IN1(n15409), .IN2(n6937), .Q(n15408) );
  AND2X1 U17237 ( .IN1(n15410), .IN2(n6970), .Q(n14560) );
  AND2X1 U17238 ( .IN1(n15411), .IN2(n6969), .Q(n14561) );
  AND2X1 U17239 ( .IN1(P2_N830), .IN2(n6820), .Q(n15412) );
  AND2X1 U17240 ( .IN1(P2_N1176), .IN2(n6819), .Q(n15413) );
  AND2X1 U17241 ( .IN1(P2_N902), .IN2(n6820), .Q(n15414) );
  AND2X1 U17242 ( .IN1(P2_N1431), .IN2(n6819), .Q(n15415) );
  AND2X1 U17243 ( .IN1(n15417), .IN2(n6790), .Q(n15416) );
  AND2X1 U17244 ( .IN1(n15419), .IN2(n6789), .Q(n15418) );
  AND2X1 U17245 ( .IN1(P2_N1804), .IN2(n6820), .Q(n15420) );
  AND2X1 U17246 ( .IN1(P2_N2550), .IN2(n6819), .Q(n15421) );
  AND2X1 U17247 ( .IN1(P2_N2177), .IN2(n6820), .Q(n15422) );
  AND2X1 U17248 ( .IN1(P2_N2923), .IN2(n6819), .Q(n15423) );
  AND2X1 U17249 ( .IN1(n15425), .IN2(n6790), .Q(n15424) );
  AND2X1 U17250 ( .IN1(n15427), .IN2(n6789), .Q(n15426) );
  AND2X1 U17251 ( .IN1(n15429), .IN2(n6948), .Q(n15428) );
  AND2X1 U17252 ( .IN1(n15431), .IN2(n6937), .Q(n15430) );
  AND2X1 U17253 ( .IN1(P2_N3296), .IN2(n6820), .Q(n15432) );
  AND2X1 U17254 ( .IN1(P2_N4042), .IN2(n6819), .Q(n15433) );
  AND2X1 U17255 ( .IN1(P2_N3669), .IN2(n6820), .Q(n15434) );
  AND2X1 U17256 ( .IN1(P2_N4416), .IN2(n6819), .Q(n15435) );
  AND2X1 U17257 ( .IN1(n15437), .IN2(n6790), .Q(n15436) );
  AND2X1 U17258 ( .IN1(n15439), .IN2(n6789), .Q(n15438) );
  AND2X1 U17259 ( .IN1(P2_N381), .IN2(n14522), .Q(n15440) );
  AND2X1 U17260 ( .IN1(P2_N4679), .IN2(n6986), .Q(n15441) );
  AND2X1 U17261 ( .IN1(n15443), .IN2(n6942), .Q(n15442) );
  AND2X1 U17262 ( .IN1(n15445), .IN2(n6937), .Q(n15444) );
  AND2X1 U17263 ( .IN1(n15446), .IN2(n6970), .Q(n14562) );
  AND2X1 U17264 ( .IN1(n15447), .IN2(n6969), .Q(n14563) );
  AND2X1 U17265 ( .IN1(P2_N831), .IN2(n6820), .Q(n15448) );
  AND2X1 U17266 ( .IN1(P2_N1177), .IN2(n6819), .Q(n15449) );
  AND2X1 U17267 ( .IN1(P2_N903), .IN2(n6820), .Q(n15450) );
  AND2X1 U17268 ( .IN1(P2_N1432), .IN2(n6819), .Q(n15451) );
  AND2X1 U17269 ( .IN1(n15453), .IN2(n6784), .Q(n15452) );
  AND2X1 U17270 ( .IN1(n15455), .IN2(n7488), .Q(n15454) );
  AND2X1 U17271 ( .IN1(P2_N1805), .IN2(n6820), .Q(n15456) );
  AND2X1 U17272 ( .IN1(P2_N2551), .IN2(n6819), .Q(n15457) );
  AND2X1 U17273 ( .IN1(P2_N2178), .IN2(n6842), .Q(n15458) );
  AND2X1 U17274 ( .IN1(P2_N2924), .IN2(n6827), .Q(n15459) );
  AND2X1 U17275 ( .IN1(n15461), .IN2(n6784), .Q(n15460) );
  AND2X1 U17276 ( .IN1(n15463), .IN2(n7488), .Q(n15462) );
  AND2X1 U17277 ( .IN1(n15465), .IN2(n6940), .Q(n15464) );
  AND2X1 U17278 ( .IN1(n15467), .IN2(n6931), .Q(n15466) );
  AND2X1 U17279 ( .IN1(P2_N3297), .IN2(n6820), .Q(n15468) );
  AND2X1 U17280 ( .IN1(P2_N4043), .IN2(n6819), .Q(n15469) );
  AND2X1 U17281 ( .IN1(P2_N3670), .IN2(n6820), .Q(n15470) );
  AND2X1 U17282 ( .IN1(P2_N4417), .IN2(n6819), .Q(n15471) );
  AND2X1 U17283 ( .IN1(n15473), .IN2(n6784), .Q(n15472) );
  AND2X1 U17284 ( .IN1(n15475), .IN2(n7488), .Q(n15474) );
  AND2X1 U17285 ( .IN1(P2_N382), .IN2(n14522), .Q(n15476) );
  AND2X1 U17286 ( .IN1(P2_N4680), .IN2(n6986), .Q(n15477) );
  AND2X1 U17287 ( .IN1(n15479), .IN2(n6940), .Q(n15478) );
  AND2X1 U17288 ( .IN1(n15481), .IN2(n6931), .Q(n15480) );
  AND2X1 U17289 ( .IN1(n15482), .IN2(n6970), .Q(n14564) );
  AND2X1 U17290 ( .IN1(n15483), .IN2(n6969), .Q(n14565) );
  AND2X1 U17291 ( .IN1(P2_N832), .IN2(n6820), .Q(n15484) );
  AND2X1 U17292 ( .IN1(P2_N1178), .IN2(n6813), .Q(n15485) );
  AND2X1 U17293 ( .IN1(P2_N904), .IN2(n6820), .Q(n15486) );
  AND2X1 U17294 ( .IN1(P2_N1433), .IN2(n6813), .Q(n15487) );
  AND2X1 U17295 ( .IN1(n15489), .IN2(n6784), .Q(n15488) );
  AND2X1 U17296 ( .IN1(n15491), .IN2(n7488), .Q(n15490) );
  AND2X1 U17297 ( .IN1(P2_N1806), .IN2(n6842), .Q(n15492) );
  AND2X1 U17298 ( .IN1(P2_N2552), .IN2(n6827), .Q(n15493) );
  AND2X1 U17299 ( .IN1(P2_N2179), .IN2(n6842), .Q(n15494) );
  AND2X1 U17300 ( .IN1(P2_N2925), .IN2(n6827), .Q(n15495) );
  AND2X1 U17301 ( .IN1(n15497), .IN2(n6784), .Q(n15496) );
  AND2X1 U17302 ( .IN1(n15499), .IN2(n6793), .Q(n15498) );
  AND2X1 U17303 ( .IN1(n15501), .IN2(n6940), .Q(n15500) );
  AND2X1 U17304 ( .IN1(n15503), .IN2(n6931), .Q(n15502) );
  AND2X1 U17305 ( .IN1(P2_N3298), .IN2(n6842), .Q(n15504) );
  AND2X1 U17306 ( .IN1(P2_N4044), .IN2(n6813), .Q(n15505) );
  AND2X1 U17307 ( .IN1(P2_N3671), .IN2(n6842), .Q(n15506) );
  AND2X1 U17308 ( .IN1(P2_N4418), .IN2(n6813), .Q(n15507) );
  AND2X1 U17309 ( .IN1(n15509), .IN2(n6784), .Q(n15508) );
  AND2X1 U17310 ( .IN1(n15511), .IN2(n6793), .Q(n15510) );
  AND2X1 U17311 ( .IN1(P2_N383), .IN2(n14522), .Q(n15512) );
  AND2X1 U17312 ( .IN1(P2_N4681), .IN2(n6986), .Q(n15513) );
  AND2X1 U17313 ( .IN1(n15515), .IN2(n6940), .Q(n15514) );
  AND2X1 U17314 ( .IN1(n15517), .IN2(n6931), .Q(n15516) );
  AND2X1 U17315 ( .IN1(n15518), .IN2(n6972), .Q(n14566) );
  AND2X1 U17316 ( .IN1(n15519), .IN2(n6963), .Q(n14567) );
  AND2X1 U17317 ( .IN1(P2_N833), .IN2(n6828), .Q(n15520) );
  AND2X1 U17318 ( .IN1(P2_N1179), .IN2(n6813), .Q(n15521) );
  AND2X1 U17319 ( .IN1(P2_N905), .IN2(n6828), .Q(n15522) );
  AND2X1 U17320 ( .IN1(P2_N1434), .IN2(n6813), .Q(n15523) );
  AND2X1 U17321 ( .IN1(n15525), .IN2(n6784), .Q(n15524) );
  AND2X1 U17322 ( .IN1(n15527), .IN2(n7488), .Q(n15526) );
  AND2X1 U17323 ( .IN1(P2_N1807), .IN2(n6842), .Q(n15528) );
  AND2X1 U17324 ( .IN1(P2_N2553), .IN2(n6827), .Q(n15529) );
  AND2X1 U17325 ( .IN1(P2_N2180), .IN2(n6842), .Q(n15530) );
  AND2X1 U17326 ( .IN1(P2_N2926), .IN2(n6827), .Q(n15531) );
  AND2X1 U17327 ( .IN1(n15533), .IN2(n6784), .Q(n15532) );
  AND2X1 U17142 ( .IN1(P2_N2546), .IN2(n6825), .Q(n15277) );
  AND2X1 U17143 ( .IN1(P2_N2173), .IN2(n6816), .Q(n15278) );
  AND2X1 U17144 ( .IN1(P2_N2919), .IN2(n6825), .Q(n15279) );
  AND2X1 U17145 ( .IN1(n15281), .IN2(n6786), .Q(n15280) );
  AND2X1 U17146 ( .IN1(n15283), .IN2(n6775), .Q(n15282) );
  AND2X1 U17147 ( .IN1(n15285), .IN2(n6946), .Q(n15284) );
  AND2X1 U17148 ( .IN1(n15287), .IN2(n6937), .Q(n15286) );
  AND2X1 U17149 ( .IN1(P2_N3292), .IN2(n6816), .Q(n15288) );
  AND2X1 U17150 ( .IN1(P2_N4038), .IN2(n6825), .Q(n15289) );
  AND2X1 U17151 ( .IN1(P2_N3665), .IN2(n6812), .Q(n15290) );
  AND2X1 U17152 ( .IN1(P2_N4412), .IN2(n6825), .Q(n15291) );
  AND2X1 U17153 ( .IN1(n15293), .IN2(n6786), .Q(n15292) );
  AND2X1 U17154 ( .IN1(n15295), .IN2(n6787), .Q(n15294) );
  AND2X1 U17155 ( .IN1(P2_N377), .IN2(n14522), .Q(n15296) );
  AND2X1 U17156 ( .IN1(P2_N4675), .IN2(n6986), .Q(n15297) );
  AND2X1 U17157 ( .IN1(n15299), .IN2(n6946), .Q(n15298) );
  AND2X1 U17158 ( .IN1(n15301), .IN2(n6941), .Q(n15300) );
  AND2X1 U17159 ( .IN1(n15302), .IN2(n6974), .Q(n14554) );
  AND2X1 U17160 ( .IN1(n15303), .IN2(n6967), .Q(n14555) );
  AND2X1 U17161 ( .IN1(P2_N827), .IN2(n6822), .Q(n15304) );
  AND2X1 U17162 ( .IN1(P2_N1173), .IN2(n7486), .Q(n15305) );
  AND2X1 U17163 ( .IN1(P2_N899), .IN2(n6822), .Q(n15306) );
  AND2X1 U17164 ( .IN1(P2_N1428), .IN2(n6825), .Q(n15307) );
  AND2X1 U17165 ( .IN1(n15309), .IN2(n6790), .Q(n15308) );
  AND2X1 U17166 ( .IN1(n15311), .IN2(n6789), .Q(n15310) );
  AND2X1 U17167 ( .IN1(P2_N1801), .IN2(n6816), .Q(n15312) );
  AND2X1 U17168 ( .IN1(P2_N2547), .IN2(n6825), .Q(n15313) );
  AND2X1 U17169 ( .IN1(P2_N2174), .IN2(n6812), .Q(n15314) );
  AND2X1 U17170 ( .IN1(P2_N2920), .IN2(n6825), .Q(n15315) );
  AND2X1 U17171 ( .IN1(n15317), .IN2(n6786), .Q(n15316) );
  AND2X1 U17172 ( .IN1(n15319), .IN2(n6775), .Q(n15318) );
  AND2X1 U17173 ( .IN1(n15321), .IN2(n6946), .Q(n15320) );
  AND2X1 U17174 ( .IN1(n15323), .IN2(n6937), .Q(n15322) );
  AND2X1 U17175 ( .IN1(P2_N3293), .IN2(n6822), .Q(n15324) );
  AND2X1 U17176 ( .IN1(P2_N4039), .IN2(n6825), .Q(n15325) );
  AND2X1 U17177 ( .IN1(P2_N3666), .IN2(n6822), .Q(n15326) );
  AND2X1 U17178 ( .IN1(P2_N4413), .IN2(n7486), .Q(n15327) );
  AND2X1 U17179 ( .IN1(n15329), .IN2(n6790), .Q(n15328) );
  AND2X1 U17180 ( .IN1(n15331), .IN2(n6789), .Q(n15330) );
  AND2X1 U17181 ( .IN1(P2_N378), .IN2(n14522), .Q(n15332) );
  AND2X1 U17182 ( .IN1(P2_N4676), .IN2(n6986), .Q(n15333) );
  AND2X1 U17183 ( .IN1(n15335), .IN2(n6942), .Q(n15334) );
  AND2X1 U17184 ( .IN1(n15337), .IN2(n6937), .Q(n15336) );
  AND2X1 U17185 ( .IN1(n15338), .IN2(n6970), .Q(n14556) );
  AND2X1 U17186 ( .IN1(n15339), .IN2(n6969), .Q(n14557) );
  AND2X1 U17187 ( .IN1(P2_N828), .IN2(n6822), .Q(n15340) );
  AND2X1 U17188 ( .IN1(P2_N1174), .IN2(n7486), .Q(n15341) );
  AND2X1 U17189 ( .IN1(P2_N900), .IN2(n6822), .Q(n15342) );
  AND2X1 U17190 ( .IN1(P2_N1429), .IN2(n7486), .Q(n15343) );
  AND2X1 U17191 ( .IN1(n15345), .IN2(n6790), .Q(n15344) );
  AND2X1 U17192 ( .IN1(n15347), .IN2(n6789), .Q(n15346) );
  AND2X1 U17193 ( .IN1(P2_N1802), .IN2(n6822), .Q(n15348) );
  AND2X1 U17194 ( .IN1(P2_N2548), .IN2(n6825), .Q(n15349) );
  AND2X1 U17195 ( .IN1(P2_N2175), .IN2(n6822), .Q(n15350) );
  AND2X1 U17196 ( .IN1(P2_N2921), .IN2(n7486), .Q(n15351) );
  AND2X1 U17197 ( .IN1(n15353), .IN2(n6790), .Q(n15352) );
  AND2X1 U17198 ( .IN1(n15355), .IN2(n6789), .Q(n15354) );
  AND2X1 U17199 ( .IN1(n15357), .IN2(n6946), .Q(n15356) );
  AND2X1 U17200 ( .IN1(n15359), .IN2(n6937), .Q(n15358) );
  AND2X1 U17201 ( .IN1(P2_N3294), .IN2(n6822), .Q(n15360) );
  AND2X1 U17202 ( .IN1(P2_N4040), .IN2(n6825), .Q(n15361) );
  AND2X1 U17203 ( .IN1(P2_N3667), .IN2(n6822), .Q(n15362) );
  AND2X1 U17204 ( .IN1(P2_N4414), .IN2(n6825), .Q(n15363) );
  AND2X1 U17205 ( .IN1(n15365), .IN2(n6790), .Q(n15364) );
  AND2X1 U17206 ( .IN1(n15367), .IN2(n6789), .Q(n15366) );
  AND2X1 U17207 ( .IN1(P2_N379), .IN2(n14522), .Q(n15368) );
  AND2X1 U17208 ( .IN1(P2_N4677), .IN2(n6986), .Q(n15369) );
  AND2X1 U17209 ( .IN1(n15371), .IN2(n6948), .Q(n15370) );
  AND2X1 U17210 ( .IN1(n15373), .IN2(n6937), .Q(n15372) );
  AND2X1 U17211 ( .IN1(n15374), .IN2(n6970), .Q(n14558) );
  AND2X1 U17212 ( .IN1(n15375), .IN2(n6969), .Q(n14559) );
  AND2X1 U17213 ( .IN1(P2_N829), .IN2(n6820), .Q(n15376) );
  AND2X1 U17214 ( .IN1(P2_N1175), .IN2(n6819), .Q(n15377) );
  AND2X1 U17215 ( .IN1(P2_N901), .IN2(n6820), .Q(n15378) );
  AND2X1 U17216 ( .IN1(P2_N1430), .IN2(n6819), .Q(n15379) );
  AND2X1 U17217 ( .IN1(n15381), .IN2(n6790), .Q(n15380) );
  AND2X1 U17218 ( .IN1(n15383), .IN2(n6789), .Q(n15382) );
  AND2X1 U17219 ( .IN1(P2_N1803), .IN2(n6822), .Q(n15384) );
  AND2X1 U17220 ( .IN1(P2_N2549), .IN2(n6825), .Q(n15385) );
  AND2X1 U17221 ( .IN1(P2_N2176), .IN2(n6822), .Q(n15386) );
  AND2X1 U17222 ( .IN1(P2_N2922), .IN2(n6825), .Q(n15387) );
  AND2X1 U17223 ( .IN1(n15389), .IN2(n6790), .Q(n15388) );
  AND2X1 U17224 ( .IN1(n15391), .IN2(n6789), .Q(n15390) );
  AND2X1 U17225 ( .IN1(n15393), .IN2(n6946), .Q(n15392) );
  AND2X1 U17226 ( .IN1(n15395), .IN2(n6937), .Q(n15394) );
  AND2X1 U17227 ( .IN1(P2_N3295), .IN2(n6820), .Q(n15396) );
  AND2X1 U17228 ( .IN1(P2_N4041), .IN2(n6819), .Q(n15397) );
  AND2X1 U17229 ( .IN1(P2_N3668), .IN2(n6822), .Q(n15398) );
  AND2X1 U17230 ( .IN1(P2_N4415), .IN2(n6819), .Q(n15399) );
  AND2X1 U17231 ( .IN1(n15401), .IN2(n6790), .Q(n15400) );
  AND2X1 U17232 ( .IN1(n15403), .IN2(n6789), .Q(n15402) );
  AND2X1 U17233 ( .IN1(P2_N380), .IN2(n14522), .Q(n15404) );
  AND2X1 U17234 ( .IN1(P2_N4678), .IN2(n6986), .Q(n15405) );
  AND2X1 U17049 ( .IN1(n15149), .IN2(n6776), .Q(n15148) );
  AND2X1 U17050 ( .IN1(n15151), .IN2(n6787), .Q(n15150) );
  AND2X1 U17051 ( .IN1(P2_N373), .IN2(n14522), .Q(n15152) );
  AND2X1 U17052 ( .IN1(P2_N4671), .IN2(n6986), .Q(n15153) );
  AND2X1 U17053 ( .IN1(n15155), .IN2(n6948), .Q(n15154) );
  AND2X1 U17054 ( .IN1(n15157), .IN2(P2_N293), .Q(n15156) );
  AND2X1 U17055 ( .IN1(n15158), .IN2(n6970), .Q(n14546) );
  AND2X1 U17056 ( .IN1(n15159), .IN2(n6963), .Q(n14547) );
  AND2X1 U17057 ( .IN1(P2_N823), .IN2(n6816), .Q(n15160) );
  AND2X1 U17058 ( .IN1(P2_N1169), .IN2(n6815), .Q(n15161) );
  AND2X1 U17059 ( .IN1(P2_N895), .IN2(n6816), .Q(n15162) );
  AND2X1 U17060 ( .IN1(P2_N1424), .IN2(n6815), .Q(n15163) );
  AND2X1 U17061 ( .IN1(n15165), .IN2(n6776), .Q(n15164) );
  AND2X1 U17062 ( .IN1(n15167), .IN2(n6787), .Q(n15166) );
  AND2X1 U17063 ( .IN1(P2_N1797), .IN2(n6818), .Q(n15168) );
  AND2X1 U17064 ( .IN1(P2_N2543), .IN2(n6823), .Q(n15169) );
  AND2X1 U17065 ( .IN1(P2_N2170), .IN2(n6818), .Q(n15170) );
  AND2X1 U17066 ( .IN1(P2_N2916), .IN2(n6823), .Q(n15171) );
  AND2X1 U17067 ( .IN1(n15173), .IN2(n6786), .Q(n15172) );
  AND2X1 U17068 ( .IN1(n15175), .IN2(n6787), .Q(n15174) );
  AND2X1 U17069 ( .IN1(n15177), .IN2(n6948), .Q(n15176) );
  AND2X1 U17070 ( .IN1(n15179), .IN2(P2_N293), .Q(n15178) );
  AND2X1 U17071 ( .IN1(P2_N3289), .IN2(n6816), .Q(n15180) );
  AND2X1 U17072 ( .IN1(P2_N4035), .IN2(n6815), .Q(n15181) );
  AND2X1 U17073 ( .IN1(P2_N3662), .IN2(n6816), .Q(n15182) );
  AND2X1 U17074 ( .IN1(P2_N4409), .IN2(n6815), .Q(n15183) );
  AND2X1 U17075 ( .IN1(n15185), .IN2(n6786), .Q(n15184) );
  AND2X1 U17076 ( .IN1(n15187), .IN2(n6787), .Q(n15186) );
  AND2X1 U17077 ( .IN1(P2_N374), .IN2(n14522), .Q(n15188) );
  AND2X1 U17078 ( .IN1(P2_N4672), .IN2(n6986), .Q(n15189) );
  AND2X1 U17079 ( .IN1(n15191), .IN2(n6948), .Q(n15190) );
  AND2X1 U17080 ( .IN1(n15193), .IN2(n6941), .Q(n15192) );
  AND2X1 U17081 ( .IN1(n15194), .IN2(n6974), .Q(n14548) );
  AND2X1 U17082 ( .IN1(n15195), .IN2(n6963), .Q(n14549) );
  AND2X1 U17083 ( .IN1(P2_N824), .IN2(n6816), .Q(n15196) );
  AND2X1 U17084 ( .IN1(P2_N1170), .IN2(n6815), .Q(n15197) );
  AND2X1 U17085 ( .IN1(P2_N896), .IN2(n6816), .Q(n15198) );
  AND2X1 U17086 ( .IN1(P2_N1425), .IN2(n6815), .Q(n15199) );
  AND2X1 U17087 ( .IN1(n15201), .IN2(n6786), .Q(n15200) );
  AND2X1 U17088 ( .IN1(n15203), .IN2(n6775), .Q(n15202) );
  AND2X1 U17089 ( .IN1(P2_N1798), .IN2(n6816), .Q(n15204) );
  AND2X1 U17090 ( .IN1(P2_N2544), .IN2(n6815), .Q(n15205) );
  AND2X1 U17091 ( .IN1(P2_N2171), .IN2(n6816), .Q(n15206) );
  AND2X1 U17092 ( .IN1(P2_N2917), .IN2(n6815), .Q(n15207) );
  AND2X1 U17093 ( .IN1(n15209), .IN2(n6776), .Q(n15208) );
  AND2X1 U17094 ( .IN1(n15211), .IN2(n6787), .Q(n15210) );
  AND2X1 U17095 ( .IN1(n15213), .IN2(n6948), .Q(n15212) );
  AND2X1 U17096 ( .IN1(n15215), .IN2(P2_N293), .Q(n15214) );
  AND2X1 U17097 ( .IN1(P2_N3290), .IN2(n6816), .Q(n15216) );
  AND2X1 U17098 ( .IN1(P2_N4036), .IN2(n6815), .Q(n15217) );
  AND2X1 U17099 ( .IN1(P2_N3663), .IN2(n6816), .Q(n15218) );
  AND2X1 U17100 ( .IN1(P2_N4410), .IN2(n6815), .Q(n15219) );
  AND2X1 U17101 ( .IN1(n15221), .IN2(n6786), .Q(n15220) );
  AND2X1 U17102 ( .IN1(n15223), .IN2(n6787), .Q(n15222) );
  AND2X1 U17103 ( .IN1(P2_N375), .IN2(n14522), .Q(n15224) );
  AND2X1 U17104 ( .IN1(P2_N4673), .IN2(n6986), .Q(n15225) );
  AND2X1 U17105 ( .IN1(n15227), .IN2(n6946), .Q(n15226) );
  AND2X1 U17106 ( .IN1(n15229), .IN2(n6941), .Q(n15228) );
  AND2X1 U17107 ( .IN1(n15230), .IN2(n6970), .Q(n14550) );
  AND2X1 U17108 ( .IN1(n15231), .IN2(n6963), .Q(n14551) );
  AND2X1 U17109 ( .IN1(P2_N825), .IN2(n6816), .Q(n15232) );
  AND2X1 U17110 ( .IN1(P2_N1171), .IN2(n6815), .Q(n15233) );
  AND2X1 U17111 ( .IN1(P2_N897), .IN2(n6816), .Q(n15234) );
  AND2X1 U17112 ( .IN1(P2_N1426), .IN2(n6815), .Q(n15235) );
  AND2X1 U17113 ( .IN1(n15237), .IN2(n6786), .Q(n15236) );
  AND2X1 U17114 ( .IN1(n15239), .IN2(n6775), .Q(n15238) );
  AND2X1 U17115 ( .IN1(P2_N1799), .IN2(n6816), .Q(n15240) );
  AND2X1 U17116 ( .IN1(P2_N2545), .IN2(n6815), .Q(n15241) );
  AND2X1 U17117 ( .IN1(P2_N2172), .IN2(n6816), .Q(n15242) );
  AND2X1 U17118 ( .IN1(P2_N2918), .IN2(n6815), .Q(n15243) );
  AND2X1 U17119 ( .IN1(n15245), .IN2(n6786), .Q(n15244) );
  AND2X1 U17120 ( .IN1(n15247), .IN2(n6775), .Q(n15246) );
  AND2X1 U17121 ( .IN1(n15249), .IN2(n6946), .Q(n15248) );
  AND2X1 U17122 ( .IN1(n15251), .IN2(n6937), .Q(n15250) );
  AND2X1 U17123 ( .IN1(P2_N3291), .IN2(n6816), .Q(n15252) );
  AND2X1 U17124 ( .IN1(P2_N4037), .IN2(n6815), .Q(n15253) );
  AND2X1 U17125 ( .IN1(P2_N3664), .IN2(n6816), .Q(n15254) );
  AND2X1 U17126 ( .IN1(P2_N4411), .IN2(n6815), .Q(n15255) );
  AND2X1 U17127 ( .IN1(n15257), .IN2(n6786), .Q(n15256) );
  AND2X1 U17128 ( .IN1(n15259), .IN2(n6787), .Q(n15258) );
  AND2X1 U17129 ( .IN1(P2_N376), .IN2(n14522), .Q(n15260) );
  AND2X1 U17130 ( .IN1(P2_N4674), .IN2(n6986), .Q(n15261) );
  AND2X1 U17131 ( .IN1(n15263), .IN2(n6946), .Q(n15262) );
  AND2X1 U17132 ( .IN1(n15265), .IN2(n6941), .Q(n15264) );
  AND2X1 U17133 ( .IN1(n15266), .IN2(n6974), .Q(n14552) );
  AND2X1 U17134 ( .IN1(n15267), .IN2(n6967), .Q(n14553) );
  AND2X1 U17135 ( .IN1(P2_N826), .IN2(n6812), .Q(n15268) );
  AND2X1 U17136 ( .IN1(P2_N1172), .IN2(n6825), .Q(n15269) );
  AND2X1 U17137 ( .IN1(P2_N898), .IN2(n6812), .Q(n15270) );
  AND2X1 U17138 ( .IN1(P2_N1427), .IN2(n6825), .Q(n15271) );
  AND2X1 U17139 ( .IN1(n15273), .IN2(n6786), .Q(n15272) );
  AND2X1 U17140 ( .IN1(n15275), .IN2(n6789), .Q(n15274) );
  AND2X1 U17141 ( .IN1(P2_N1800), .IN2(n6812), .Q(n15276) );
  AND2X1 U16956 ( .IN1(P2_N1420), .IN2(n6843), .Q(n15019) );
  AND2X1 U16957 ( .IN1(n15021), .IN2(n6786), .Q(n15020) );
  AND2X1 U16958 ( .IN1(n15023), .IN2(n6787), .Q(n15022) );
  AND2X1 U16959 ( .IN1(P2_N1793), .IN2(n6852), .Q(n15024) );
  AND2X1 U16960 ( .IN1(P2_N2539), .IN2(n6843), .Q(n15025) );
  AND2X1 U16961 ( .IN1(P2_N2166), .IN2(n6836), .Q(n15026) );
  AND2X1 U16962 ( .IN1(P2_N2912), .IN2(n6843), .Q(n15027) );
  AND2X1 U16963 ( .IN1(n15029), .IN2(n6776), .Q(n15028) );
  AND2X1 U16964 ( .IN1(n15031), .IN2(n6787), .Q(n15030) );
  AND2X1 U16965 ( .IN1(n15033), .IN2(n6948), .Q(n15032) );
  AND2X1 U16966 ( .IN1(n15035), .IN2(P2_N293), .Q(n15034) );
  AND2X1 U16967 ( .IN1(P2_N3285), .IN2(n6818), .Q(n15036) );
  AND2X1 U16968 ( .IN1(P2_N4031), .IN2(n6843), .Q(n15037) );
  AND2X1 U16969 ( .IN1(P2_N3658), .IN2(n6852), .Q(n15038) );
  AND2X1 U16970 ( .IN1(P2_N4405), .IN2(n6843), .Q(n15039) );
  AND2X1 U16971 ( .IN1(n15041), .IN2(n6776), .Q(n15040) );
  AND2X1 U16972 ( .IN1(n15043), .IN2(n6787), .Q(n15042) );
  AND2X1 U16973 ( .IN1(P2_N370), .IN2(n14522), .Q(n15044) );
  AND2X1 U16974 ( .IN1(P2_N4668), .IN2(n6986), .Q(n15045) );
  AND2X1 U16975 ( .IN1(n15047), .IN2(n6948), .Q(n15046) );
  AND2X1 U16976 ( .IN1(n15049), .IN2(P2_N293), .Q(n15048) );
  AND2X1 U16977 ( .IN1(n15050), .IN2(n6970), .Q(n14540) );
  AND2X1 U16978 ( .IN1(n15051), .IN2(n6963), .Q(n14541) );
  AND2X1 U16979 ( .IN1(P2_N820), .IN2(n6824), .Q(n15052) );
  AND2X1 U16980 ( .IN1(P2_N1166), .IN2(n6843), .Q(n15053) );
  AND2X1 U16981 ( .IN1(P2_N892), .IN2(n6824), .Q(n15054) );
  AND2X1 U16982 ( .IN1(P2_N1421), .IN2(n6843), .Q(n15055) );
  AND2X1 U16983 ( .IN1(n15057), .IN2(n6776), .Q(n15056) );
  AND2X1 U16984 ( .IN1(n15059), .IN2(n6787), .Q(n15058) );
  AND2X1 U16985 ( .IN1(P2_N1794), .IN2(n6818), .Q(n15060) );
  AND2X1 U16986 ( .IN1(P2_N2540), .IN2(n6823), .Q(n15061) );
  AND2X1 U16987 ( .IN1(P2_N2167), .IN2(n6818), .Q(n15062) );
  AND2X1 U16988 ( .IN1(P2_N2913), .IN2(n6823), .Q(n15063) );
  AND2X1 U16989 ( .IN1(n15065), .IN2(n6786), .Q(n15064) );
  AND2X1 U16990 ( .IN1(n15067), .IN2(n6787), .Q(n15066) );
  AND2X1 U16991 ( .IN1(n15069), .IN2(n6948), .Q(n15068) );
  AND2X1 U16992 ( .IN1(n15071), .IN2(P2_N293), .Q(n15070) );
  AND2X1 U16993 ( .IN1(P2_N3286), .IN2(n6818), .Q(n15072) );
  AND2X1 U16994 ( .IN1(P2_N4032), .IN2(n6823), .Q(n15073) );
  AND2X1 U16995 ( .IN1(P2_N3659), .IN2(n6818), .Q(n15074) );
  AND2X1 U16996 ( .IN1(P2_N4406), .IN2(n6823), .Q(n15075) );
  AND2X1 U16997 ( .IN1(n15077), .IN2(n6786), .Q(n15076) );
  AND2X1 U16998 ( .IN1(n15079), .IN2(n6787), .Q(n15078) );
  AND2X1 U16999 ( .IN1(P2_N371), .IN2(n14522), .Q(n15080) );
  AND2X1 U17000 ( .IN1(P2_N4669), .IN2(n6986), .Q(n15081) );
  AND2X1 U17001 ( .IN1(n15083), .IN2(n6948), .Q(n15082) );
  AND2X1 U17002 ( .IN1(n15085), .IN2(P2_N293), .Q(n15084) );
  AND2X1 U17003 ( .IN1(n15086), .IN2(n6970), .Q(n14542) );
  AND2X1 U17004 ( .IN1(n15087), .IN2(n6963), .Q(n14543) );
  AND2X1 U17005 ( .IN1(P2_N821), .IN2(n6824), .Q(n15088) );
  AND2X1 U17006 ( .IN1(P2_N1167), .IN2(n6843), .Q(n15089) );
  AND2X1 U17007 ( .IN1(P2_N893), .IN2(n6824), .Q(n15090) );
  AND2X1 U17008 ( .IN1(P2_N1422), .IN2(n6843), .Q(n15091) );
  AND2X1 U17009 ( .IN1(n15093), .IN2(n6790), .Q(n15092) );
  AND2X1 U17010 ( .IN1(n15095), .IN2(n6787), .Q(n15094) );
  AND2X1 U17011 ( .IN1(P2_N1795), .IN2(n6818), .Q(n15096) );
  AND2X1 U17012 ( .IN1(P2_N2541), .IN2(n6823), .Q(n15097) );
  AND2X1 U17013 ( .IN1(P2_N2168), .IN2(n6818), .Q(n15098) );
  AND2X1 U17014 ( .IN1(P2_N2914), .IN2(n6823), .Q(n15099) );
  AND2X1 U17015 ( .IN1(n15101), .IN2(n6776), .Q(n15100) );
  AND2X1 U17016 ( .IN1(n15103), .IN2(n6787), .Q(n15102) );
  AND2X1 U17017 ( .IN1(n15105), .IN2(n6948), .Q(n15104) );
  AND2X1 U17018 ( .IN1(n15107), .IN2(P2_N293), .Q(n15106) );
  AND2X1 U17019 ( .IN1(P2_N3287), .IN2(n6818), .Q(n15108) );
  AND2X1 U17020 ( .IN1(P2_N4033), .IN2(n6823), .Q(n15109) );
  AND2X1 U17021 ( .IN1(P2_N3660), .IN2(n6818), .Q(n15110) );
  AND2X1 U17022 ( .IN1(P2_N4407), .IN2(n6823), .Q(n15111) );
  AND2X1 U17023 ( .IN1(n15113), .IN2(n6776), .Q(n15112) );
  AND2X1 U17024 ( .IN1(n15115), .IN2(n6787), .Q(n15114) );
  AND2X1 U17025 ( .IN1(P2_N372), .IN2(n14522), .Q(n15116) );
  AND2X1 U17026 ( .IN1(P2_N4670), .IN2(n6986), .Q(n15117) );
  AND2X1 U17027 ( .IN1(n15119), .IN2(n6948), .Q(n15118) );
  AND2X1 U17028 ( .IN1(n15121), .IN2(P2_N293), .Q(n15120) );
  AND2X1 U17029 ( .IN1(n15122), .IN2(n6974), .Q(n14544) );
  AND2X1 U17030 ( .IN1(n15123), .IN2(n6963), .Q(n14545) );
  AND2X1 U17031 ( .IN1(P2_N822), .IN2(n6852), .Q(n15124) );
  AND2X1 U17032 ( .IN1(P2_N1168), .IN2(n6823), .Q(n15125) );
  AND2X1 U17033 ( .IN1(P2_N894), .IN2(n6852), .Q(n15126) );
  AND2X1 U17034 ( .IN1(P2_N1423), .IN2(n6843), .Q(n15127) );
  AND2X1 U17035 ( .IN1(n15129), .IN2(n6776), .Q(n15128) );
  AND2X1 U17036 ( .IN1(n15131), .IN2(n6787), .Q(n15130) );
  AND2X1 U17037 ( .IN1(P2_N1796), .IN2(n6818), .Q(n15132) );
  AND2X1 U17038 ( .IN1(P2_N2542), .IN2(n6823), .Q(n15133) );
  AND2X1 U17039 ( .IN1(P2_N2169), .IN2(n6818), .Q(n15134) );
  AND2X1 U17040 ( .IN1(P2_N2915), .IN2(n6823), .Q(n15135) );
  AND2X1 U17041 ( .IN1(n15137), .IN2(n6776), .Q(n15136) );
  AND2X1 U17042 ( .IN1(n15139), .IN2(n6787), .Q(n15138) );
  AND2X1 U17043 ( .IN1(n15141), .IN2(n6948), .Q(n15140) );
  AND2X1 U17044 ( .IN1(n15143), .IN2(P2_N293), .Q(n15142) );
  AND2X1 U17045 ( .IN1(P2_N3288), .IN2(n6818), .Q(n15144) );
  AND2X1 U17046 ( .IN1(P2_N4034), .IN2(n6823), .Q(n15145) );
  AND2X1 U17047 ( .IN1(P2_N3661), .IN2(n6818), .Q(n15146) );
  AND2X1 U17048 ( .IN1(P2_N4408), .IN2(n6823), .Q(n15147) );
  AND2X1 U16863 ( .IN1(P2_N3281), .IN2(n6836), .Q(n14892) );
  AND2X1 U16864 ( .IN1(P2_N4027), .IN2(P2_N292), .Q(n14893) );
  AND2X1 U16865 ( .IN1(P2_N3654), .IN2(n6852), .Q(n14894) );
  AND2X1 U16866 ( .IN1(P2_N4401), .IN2(P2_N292), .Q(n14895) );
  AND2X1 U16867 ( .IN1(n14897), .IN2(n6776), .Q(n14896) );
  AND2X1 U16868 ( .IN1(n14899), .IN2(n6775), .Q(n14898) );
  AND2X1 U16869 ( .IN1(n6683), .IN2(n14522), .Q(n14900) );
  AND2X1 U16870 ( .IN1(P2_N4664), .IN2(n6986), .Q(n14901) );
  AND2X1 U16871 ( .IN1(n14903), .IN2(n6942), .Q(n14902) );
  AND2X1 U16872 ( .IN1(n14905), .IN2(n6941), .Q(n14904) );
  AND2X1 U16873 ( .IN1(n14906), .IN2(n6970), .Q(n14532) );
  AND2X1 U16874 ( .IN1(n14907), .IN2(n6963), .Q(n14533) );
  AND2X1 U16875 ( .IN1(P2_N816), .IN2(n6824), .Q(n14908) );
  AND2X1 U16876 ( .IN1(P2_N1162), .IN2(P2_N292), .Q(n14909) );
  AND2X1 U16877 ( .IN1(P2_N888), .IN2(n6818), .Q(n14910) );
  AND2X1 U16878 ( .IN1(P2_N1417), .IN2(P2_N292), .Q(n14911) );
  AND2X1 U16879 ( .IN1(n14913), .IN2(n6786), .Q(n14912) );
  AND2X1 U16880 ( .IN1(n14915), .IN2(n6775), .Q(n14914) );
  AND2X1 U16881 ( .IN1(P2_N1790), .IN2(n6852), .Q(n14916) );
  AND2X1 U16882 ( .IN1(P2_N2536), .IN2(n6851), .Q(n14917) );
  AND2X1 U16883 ( .IN1(P2_N2163), .IN2(n6818), .Q(n14918) );
  AND2X1 U16884 ( .IN1(P2_N2909), .IN2(P2_N292), .Q(n14919) );
  AND2X1 U16885 ( .IN1(n14921), .IN2(n6790), .Q(n14920) );
  AND2X1 U16886 ( .IN1(n14923), .IN2(n7487), .Q(n14922) );
  AND2X1 U16887 ( .IN1(n14925), .IN2(n6948), .Q(n14924) );
  AND2X1 U16888 ( .IN1(n14927), .IN2(P2_N293), .Q(n14926) );
  AND2X1 U16889 ( .IN1(P2_N3282), .IN2(n6852), .Q(n14928) );
  AND2X1 U16890 ( .IN1(P2_N4028), .IN2(n6851), .Q(n14929) );
  AND2X1 U16891 ( .IN1(P2_N3655), .IN2(n6852), .Q(n14930) );
  AND2X1 U16892 ( .IN1(P2_N4402), .IN2(n6851), .Q(n14931) );
  AND2X1 U16893 ( .IN1(n14933), .IN2(n6786), .Q(n14932) );
  AND2X1 U16894 ( .IN1(n14935), .IN2(n7487), .Q(n14934) );
  AND2X1 U16895 ( .IN1(n18813), .IN2(n14522), .Q(n14936) );
  AND2X1 U16896 ( .IN1(P2_N4665), .IN2(n6986), .Q(n14937) );
  AND2X1 U16897 ( .IN1(n14939), .IN2(n6948), .Q(n14938) );
  AND2X1 U16898 ( .IN1(n14941), .IN2(n6941), .Q(n14940) );
  AND2X1 U16899 ( .IN1(n14942), .IN2(n6974), .Q(n14534) );
  AND2X1 U16900 ( .IN1(n14943), .IN2(n6963), .Q(n14535) );
  AND2X1 U16901 ( .IN1(P2_N817), .IN2(n6852), .Q(n14944) );
  AND2X1 U16902 ( .IN1(P2_N1163), .IN2(P2_N292), .Q(n14945) );
  AND2X1 U16903 ( .IN1(P2_N889), .IN2(n6818), .Q(n14946) );
  AND2X1 U16904 ( .IN1(P2_N1418), .IN2(P2_N292), .Q(n14947) );
  AND2X1 U16905 ( .IN1(n14949), .IN2(n6786), .Q(n14948) );
  AND2X1 U16906 ( .IN1(n14951), .IN2(n7487), .Q(n14950) );
  AND2X1 U16907 ( .IN1(P2_N1791), .IN2(n6852), .Q(n14952) );
  AND2X1 U16908 ( .IN1(P2_N2537), .IN2(n6851), .Q(n14953) );
  AND2X1 U16909 ( .IN1(P2_N2164), .IN2(n6852), .Q(n14954) );
  AND2X1 U16910 ( .IN1(P2_N2910), .IN2(P2_N292), .Q(n14955) );
  AND2X1 U16911 ( .IN1(n14957), .IN2(n6790), .Q(n14956) );
  AND2X1 U16912 ( .IN1(n14959), .IN2(n7487), .Q(n14958) );
  AND2X1 U16913 ( .IN1(n14961), .IN2(n6948), .Q(n14960) );
  AND2X1 U16914 ( .IN1(n14963), .IN2(P2_N293), .Q(n14962) );
  AND2X1 U16915 ( .IN1(P2_N3283), .IN2(n6852), .Q(n14964) );
  AND2X1 U16916 ( .IN1(P2_N4029), .IN2(n6851), .Q(n14965) );
  AND2X1 U16917 ( .IN1(P2_N3656), .IN2(n6852), .Q(n14966) );
  AND2X1 U16918 ( .IN1(P2_N4403), .IN2(n6851), .Q(n14967) );
  AND2X1 U16919 ( .IN1(n14969), .IN2(n6790), .Q(n14968) );
  AND2X1 U16920 ( .IN1(n14971), .IN2(n7487), .Q(n14970) );
  AND2X1 U16921 ( .IN1(P2_N368), .IN2(n14522), .Q(n14972) );
  AND2X1 U16922 ( .IN1(P2_N4666), .IN2(n6986), .Q(n14973) );
  AND2X1 U16923 ( .IN1(n14975), .IN2(n6946), .Q(n14974) );
  AND2X1 U16924 ( .IN1(n14977), .IN2(P2_N293), .Q(n14976) );
  AND2X1 U16925 ( .IN1(n14978), .IN2(n6974), .Q(n14536) );
  AND2X1 U16926 ( .IN1(n14979), .IN2(n6963), .Q(n14537) );
  AND2X1 U16927 ( .IN1(P2_N818), .IN2(n6852), .Q(n14980) );
  AND2X1 U16928 ( .IN1(P2_N1164), .IN2(n6843), .Q(n14981) );
  AND2X1 U16929 ( .IN1(P2_N890), .IN2(n6824), .Q(n14982) );
  AND2X1 U16930 ( .IN1(P2_N1419), .IN2(n6843), .Q(n14983) );
  AND2X1 U16931 ( .IN1(n14985), .IN2(n6790), .Q(n14984) );
  AND2X1 U16932 ( .IN1(n14987), .IN2(n7487), .Q(n14986) );
  AND2X1 U16933 ( .IN1(P2_N1792), .IN2(n6824), .Q(n14988) );
  AND2X1 U16934 ( .IN1(P2_N2538), .IN2(n6843), .Q(n14989) );
  AND2X1 U16935 ( .IN1(P2_N2165), .IN2(n6852), .Q(n14990) );
  AND2X1 U16936 ( .IN1(P2_N2911), .IN2(n6843), .Q(n14991) );
  AND2X1 U16937 ( .IN1(n14993), .IN2(n6792), .Q(n14992) );
  AND2X1 U16938 ( .IN1(n14995), .IN2(n6787), .Q(n14994) );
  AND2X1 U16939 ( .IN1(n14997), .IN2(n6946), .Q(n14996) );
  AND2X1 U16940 ( .IN1(n14999), .IN2(P2_N293), .Q(n14998) );
  AND2X1 U16941 ( .IN1(P2_N3284), .IN2(n6852), .Q(n15000) );
  AND2X1 U16942 ( .IN1(P2_N4030), .IN2(n6843), .Q(n15001) );
  AND2X1 U16943 ( .IN1(P2_N3657), .IN2(n6836), .Q(n15002) );
  AND2X1 U16944 ( .IN1(P2_N4404), .IN2(n6843), .Q(n15003) );
  AND2X1 U16945 ( .IN1(n15005), .IN2(n6786), .Q(n15004) );
  AND2X1 U16946 ( .IN1(n15007), .IN2(n7487), .Q(n15006) );
  AND2X1 U16947 ( .IN1(P2_N369), .IN2(n14522), .Q(n15008) );
  AND2X1 U16948 ( .IN1(P2_N4667), .IN2(n6986), .Q(n15009) );
  AND2X1 U16949 ( .IN1(n15011), .IN2(n6948), .Q(n15010) );
  AND2X1 U16950 ( .IN1(n15013), .IN2(P2_N293), .Q(n15012) );
  AND2X1 U16951 ( .IN1(n15014), .IN2(n6974), .Q(n14538) );
  AND2X1 U16952 ( .IN1(n15015), .IN2(n6963), .Q(n14539) );
  AND2X1 U16953 ( .IN1(P2_N819), .IN2(n6852), .Q(n15016) );
  AND2X1 U16954 ( .IN1(P2_N1165), .IN2(n6843), .Q(n15017) );
  AND2X1 U16955 ( .IN1(P2_N891), .IN2(n6824), .Q(n15018) );
  AND2X1 U16770 ( .IN1(n6793), .IN2(n14763), .Q(n14762) );
  AND2X1 U16771 ( .IN1(n14523), .IN2(n6794), .Q(n14764) );
  AND2X1 U16772 ( .IN1(n17734), .IN2(n6838), .Q(n14765) );
  AND2X1 U16773 ( .IN1(P2_N5135), .IN2(n6837), .Q(n14766) );
  AND2X1 U16774 ( .IN1(P2_N5065), .IN2(n6838), .Q(n14767) );
  AND2X1 U16775 ( .IN1(P2_N5204), .IN2(n6837), .Q(n14768) );
  AND2X1 U16776 ( .IN1(n14770), .IN2(n6784), .Q(n14769) );
  AND2X1 U16777 ( .IN1(n14772), .IN2(n6793), .Q(n14771) );
  AND2X1 U16778 ( .IN1(n14774), .IN2(n6940), .Q(n14773) );
  AND2X1 U16779 ( .IN1(n6931), .IN2(n14776), .Q(n14775) );
  AND2X1 U16780 ( .IN1(P2_N5206), .IN2(n6838), .Q(n14777) );
  AND2X1 U16781 ( .IN1(P2_N5210), .IN2(n6837), .Q(n14778) );
  AND2X1 U16782 ( .IN1(P2_N5208), .IN2(n6838), .Q(n14779) );
  AND2X1 U16783 ( .IN1(P2_N5212), .IN2(n6837), .Q(n14780) );
  AND2X1 U16784 ( .IN1(n14782), .IN2(n6784), .Q(n14781) );
  AND2X1 U16785 ( .IN1(n14784), .IN2(n6793), .Q(n14783) );
  AND2X1 U16786 ( .IN1(P2_N5214), .IN2(n6838), .Q(n14785) );
  AND2X1 U16787 ( .IN1(P2_N5285), .IN2(n6837), .Q(n14786) );
  AND2X1 U16788 ( .IN1(P2_N5216), .IN2(n6838), .Q(n14787) );
  AND2X1 U16789 ( .IN1(P2_N5354), .IN2(n6837), .Q(n14788) );
  AND2X1 U16790 ( .IN1(n14790), .IN2(n6784), .Q(n14789) );
  AND2X1 U16791 ( .IN1(n14792), .IN2(n6793), .Q(n14791) );
  AND2X1 U16792 ( .IN1(n14794), .IN2(n6940), .Q(n14793) );
  AND2X1 U16793 ( .IN1(n14796), .IN2(n6931), .Q(n14795) );
  AND2X1 U16795 ( .IN1(n14798), .IN2(n6972), .Q(n14526) );
  AND2X1 U16796 ( .IN1(n6963), .IN2(n14799), .Q(n14527) );
  AND2X1 U16797 ( .IN1(P2_N813), .IN2(n6836), .Q(n14800) );
  AND2X1 U16798 ( .IN1(P2_N1159), .IN2(n6835), .Q(n14801) );
  AND2X1 U16799 ( .IN1(P2_N885), .IN2(n6836), .Q(n14802) );
  AND2X1 U16800 ( .IN1(P2_N1414), .IN2(n6835), .Q(n14803) );
  AND2X1 U16801 ( .IN1(n14805), .IN2(n6776), .Q(n14804) );
  AND2X1 U16802 ( .IN1(n14807), .IN2(n6775), .Q(n14806) );
  AND2X1 U16803 ( .IN1(P2_N1787), .IN2(n6852), .Q(n14808) );
  AND2X1 U16804 ( .IN1(P2_N2533), .IN2(P2_N292), .Q(n14809) );
  AND2X1 U16805 ( .IN1(P2_N2160), .IN2(n6836), .Q(n14810) );
  AND2X1 U16806 ( .IN1(P2_N2906), .IN2(n6835), .Q(n14811) );
  AND2X1 U16807 ( .IN1(n14813), .IN2(n6776), .Q(n14812) );
  AND2X1 U16808 ( .IN1(n14815), .IN2(n6775), .Q(n14814) );
  AND2X1 U16809 ( .IN1(n14817), .IN2(n6946), .Q(n14816) );
  AND2X1 U16810 ( .IN1(n14819), .IN2(n6937), .Q(n14818) );
  AND2X1 U16811 ( .IN1(P2_N3279), .IN2(n6824), .Q(n14820) );
  AND2X1 U16812 ( .IN1(P2_N4025), .IN2(P2_N292), .Q(n14821) );
  AND2X1 U16813 ( .IN1(P2_N3652), .IN2(n6824), .Q(n14822) );
  AND2X1 U16814 ( .IN1(P2_N4399), .IN2(P2_N292), .Q(n14823) );
  AND2X1 U16815 ( .IN1(n14825), .IN2(n6776), .Q(n14824) );
  AND2X1 U16816 ( .IN1(n14827), .IN2(n6775), .Q(n14826) );
  AND2X1 U16817 ( .IN1(n6681), .IN2(n14522), .Q(n14828) );
  AND2X1 U16818 ( .IN1(P2_N4662), .IN2(n6986), .Q(n14829) );
  AND2X1 U16819 ( .IN1(n14831), .IN2(n6946), .Q(n14830) );
  AND2X1 U16820 ( .IN1(n14833), .IN2(n6937), .Q(n14832) );
  AND2X1 U16821 ( .IN1(n14834), .IN2(n6974), .Q(n14528) );
  AND2X1 U16822 ( .IN1(n14835), .IN2(n6967), .Q(n14529) );
  AND2X1 U16823 ( .IN1(P2_N814), .IN2(n6836), .Q(n14836) );
  AND2X1 U16824 ( .IN1(P2_N1160), .IN2(n6835), .Q(n14837) );
  AND2X1 U16825 ( .IN1(P2_N886), .IN2(n6836), .Q(n14838) );
  AND2X1 U16826 ( .IN1(P2_N1415), .IN2(n6835), .Q(n14839) );
  AND2X1 U16827 ( .IN1(n14841), .IN2(n6776), .Q(n14840) );
  AND2X1 U16828 ( .IN1(n14843), .IN2(n6775), .Q(n14842) );
  AND2X1 U16829 ( .IN1(P2_N1788), .IN2(n6818), .Q(n14844) );
  AND2X1 U16830 ( .IN1(P2_N2534), .IN2(P2_N292), .Q(n14845) );
  AND2X1 U16831 ( .IN1(P2_N2161), .IN2(n6836), .Q(n14846) );
  AND2X1 U16832 ( .IN1(P2_N2907), .IN2(n6835), .Q(n14847) );
  AND2X1 U16833 ( .IN1(n14849), .IN2(n6776), .Q(n14848) );
  AND2X1 U16834 ( .IN1(n14851), .IN2(n6775), .Q(n14850) );
  AND2X1 U16835 ( .IN1(n14853), .IN2(n6942), .Q(n14852) );
  AND2X1 U16836 ( .IN1(n14855), .IN2(n6941), .Q(n14854) );
  AND2X1 U16837 ( .IN1(P2_N3280), .IN2(n6818), .Q(n14856) );
  AND2X1 U16838 ( .IN1(P2_N4026), .IN2(P2_N292), .Q(n14857) );
  AND2X1 U16839 ( .IN1(P2_N3653), .IN2(n6818), .Q(n14858) );
  AND2X1 U16840 ( .IN1(P2_N4400), .IN2(P2_N292), .Q(n14859) );
  AND2X1 U16841 ( .IN1(n14861), .IN2(n6776), .Q(n14860) );
  AND2X1 U16842 ( .IN1(n14863), .IN2(n6775), .Q(n14862) );
  AND2X1 U16843 ( .IN1(n6682), .IN2(n14522), .Q(n14864) );
  AND2X1 U16844 ( .IN1(P2_N4663), .IN2(n6986), .Q(n14865) );
  AND2X1 U16845 ( .IN1(n14867), .IN2(n6942), .Q(n14866) );
  AND2X1 U16846 ( .IN1(n14869), .IN2(n6937), .Q(n14868) );
  AND2X1 U16847 ( .IN1(n14870), .IN2(n6974), .Q(n14530) );
  AND2X1 U16848 ( .IN1(n14871), .IN2(n6967), .Q(n14531) );
  AND2X1 U16849 ( .IN1(P2_N815), .IN2(n6836), .Q(n14872) );
  AND2X1 U16850 ( .IN1(P2_N1161), .IN2(n6835), .Q(n14873) );
  AND2X1 U16851 ( .IN1(P2_N887), .IN2(n6836), .Q(n14874) );
  AND2X1 U16852 ( .IN1(P2_N1416), .IN2(n6835), .Q(n14875) );
  AND2X1 U16853 ( .IN1(n14877), .IN2(n6776), .Q(n14876) );
  AND2X1 U16854 ( .IN1(n14879), .IN2(n6775), .Q(n14878) );
  AND2X1 U16855 ( .IN1(P2_N1789), .IN2(n6818), .Q(n14880) );
  AND2X1 U16856 ( .IN1(P2_N2535), .IN2(P2_N292), .Q(n14881) );
  AND2X1 U16857 ( .IN1(P2_N2162), .IN2(n6818), .Q(n14882) );
  AND2X1 U16858 ( .IN1(P2_N2908), .IN2(n6835), .Q(n14883) );
  AND2X1 U16859 ( .IN1(n14885), .IN2(n6776), .Q(n14884) );
  AND2X1 U16860 ( .IN1(n14887), .IN2(n6775), .Q(n14886) );
  AND2X1 U16861 ( .IN1(n14889), .IN2(n6942), .Q(n14888) );
  AND2X1 U16862 ( .IN1(n14891), .IN2(n6941), .Q(n14890) );
  OR2X1 U16677 ( .IN2(n14585), .IN1(n14584), .Q(P2_N4838) );
  OR2X1 U16678 ( .IN2(n14587), .IN1(n14586), .Q(P2_N4778) );
  OR2X1 U16679 ( .IN2(n14589), .IN1(n14588), .Q(P2_N4779) );
  OR2X1 U16680 ( .IN2(n14591), .IN1(n14590), .Q(P2_N4780) );
  OR2X1 U16681 ( .IN2(n14593), .IN1(n14592), .Q(P2_N4781) );
  OR2X1 U16682 ( .IN2(n14595), .IN1(n14594), .Q(P2_N4782) );
  OR2X1 U16683 ( .IN2(n14597), .IN1(n14596), .Q(P2_N4783) );
  OR2X1 U16684 ( .IN2(n14599), .IN1(n14598), .Q(P2_N4784) );
  OR2X1 U16685 ( .IN2(n14601), .IN1(n14600), .Q(P2_N4785) );
  OR2X1 U16686 ( .IN2(n14603), .IN1(n14602), .Q(P2_N4786) );
  OR2X1 U16687 ( .IN2(n14605), .IN1(n14604), .Q(P2_N4787) );
  OR2X1 U16688 ( .IN2(n14607), .IN1(n14606), .Q(P2_N4788) );
  OR2X1 U16689 ( .IN2(n14609), .IN1(n14608), .Q(P2_N4789) );
  OR2X1 U16690 ( .IN2(n14611), .IN1(n14610), .Q(P2_N4790) );
  OR2X1 U16691 ( .IN2(n14613), .IN1(n14612), .Q(P2_N4791) );
  OR2X1 U16692 ( .IN2(n14615), .IN1(n14614), .Q(P2_N4792) );
  OR2X1 U16693 ( .IN2(n14617), .IN1(n14616), .Q(P2_N4793) );
  OR2X1 U16694 ( .IN2(n14619), .IN1(n14618), .Q(P2_N4794) );
  OR2X1 U16695 ( .IN2(n14621), .IN1(n14620), .Q(P2_N4795) );
  OR2X1 U16696 ( .IN2(n14623), .IN1(n14622), .Q(P2_N4796) );
  OR2X1 U16697 ( .IN2(n14625), .IN1(n14624), .Q(P2_N4797) );
  OR2X1 U16698 ( .IN2(n14627), .IN1(n14626), .Q(P2_N4798) );
  OR2X1 U16699 ( .IN2(n14629), .IN1(n14628), .Q(P2_N4799) );
  OR2X1 U16700 ( .IN2(n14631), .IN1(n14630), .Q(P2_N4800) );
  OR2X1 U16701 ( .IN2(n14633), .IN1(n14632), .Q(P2_N4801) );
  OR2X1 U16702 ( .IN2(n14635), .IN1(n14634), .Q(P2_N4802) );
  OR2X1 U16703 ( .IN2(n14637), .IN1(n14636), .Q(P2_N4803) );
  OR2X1 U16704 ( .IN2(n14639), .IN1(n14638), .Q(P2_N4804) );
  OR2X1 U16705 ( .IN2(n14641), .IN1(n14640), .Q(P2_N4805) );
  OR2X1 U16706 ( .IN2(n14643), .IN1(n14642), .Q(P2_N4806) );
  OR2X1 U16707 ( .IN2(n14645), .IN1(n14644), .Q(P2_N4807) );
  OR2X1 U16708 ( .IN2(n14647), .IN1(n14646), .Q(P2_N4745) );
  OR2X1 U16709 ( .IN2(n14649), .IN1(n14648), .Q(P2_N4746) );
  OR2X1 U16710 ( .IN2(n14651), .IN1(n14650), .Q(P2_N4747) );
  OR2X1 U16711 ( .IN2(n14653), .IN1(n14652), .Q(P2_N4748) );
  OR2X1 U16712 ( .IN2(n14655), .IN1(n14654), .Q(P2_N4749) );
  OR2X1 U16713 ( .IN2(n14657), .IN1(n14656), .Q(P2_N4750) );
  OR2X1 U16714 ( .IN2(n14659), .IN1(n14658), .Q(P2_N4751) );
  OR2X1 U16715 ( .IN2(n14661), .IN1(n14660), .Q(P2_N4752) );
  OR2X1 U16716 ( .IN2(n14663), .IN1(n14662), .Q(P2_N4753) );
  OR2X1 U16717 ( .IN2(n14665), .IN1(n14664), .Q(P2_N4754) );
  OR2X1 U16718 ( .IN2(n14667), .IN1(n14666), .Q(P2_N4755) );
  OR2X1 U16719 ( .IN2(n14669), .IN1(n14668), .Q(P2_N4756) );
  OR2X1 U16720 ( .IN2(n14671), .IN1(n14670), .Q(P2_N4757) );
  OR2X1 U16721 ( .IN2(n14673), .IN1(n14672), .Q(P2_N4758) );
  OR2X1 U16722 ( .IN2(n14675), .IN1(n14674), .Q(P2_N4759) );
  OR2X1 U16723 ( .IN2(n14677), .IN1(n14676), .Q(P2_N4760) );
  OR2X1 U16724 ( .IN2(n14679), .IN1(n14678), .Q(P2_N4761) );
  OR2X1 U16725 ( .IN2(n14681), .IN1(n14680), .Q(P2_N4762) );
  OR2X1 U16726 ( .IN2(n14683), .IN1(n14682), .Q(P2_N4763) );
  OR2X1 U16727 ( .IN2(n14685), .IN1(n14684), .Q(P2_N4764) );
  OR2X1 U16728 ( .IN2(n14687), .IN1(n14686), .Q(P2_N4765) );
  OR2X1 U16729 ( .IN2(n14689), .IN1(n14688), .Q(P2_N4766) );
  OR2X1 U16730 ( .IN2(n14691), .IN1(n14690), .Q(P2_N4767) );
  OR2X1 U16731 ( .IN2(n14693), .IN1(n14692), .Q(P2_N4768) );
  OR2X1 U16732 ( .IN2(n14695), .IN1(n14694), .Q(P2_N4769) );
  OR2X1 U16733 ( .IN2(n14697), .IN1(n14696), .Q(P2_N4770) );
  OR2X1 U16734 ( .IN2(n14699), .IN1(n14698), .Q(P2_N4771) );
  OR2X1 U16735 ( .IN2(n14701), .IN1(n14700), .Q(P2_N4772) );
  OR2X1 U16736 ( .IN2(n14703), .IN1(n14702), .Q(P2_N4773) );
  OR2X1 U16737 ( .IN2(n14705), .IN1(n14704), .Q(P2_N4774) );
  AND2X1 U16738 ( .IN1(P2_N4691), .IN2(n6986), .Q(n14706) );
  OR2X1 U16739 ( .IN2(n14709), .IN1(n14708), .Q(P2_N4777) );
  AND2X1 U16740 ( .IN1(n7402), .IN2(n6986), .Q(n14710) );
  AND2X1 U16741 ( .IN1(P2_N1444), .IN2(n6837), .Q(n14711) );
  OR2X1 U16742 ( .IN2(n14713), .IN1(n14712), .Q(P2_N4744) );
  AND2X1 U16743 ( .IN1(P2_N4661), .IN2(n6986), .Q(n14714) );
  AND2X1 U16744 ( .IN1(P2_N1443), .IN2(n6837), .Q(n14715) );
  OR2X1 U16745 ( .IN2(n14717), .IN1(n14716), .Q(P2_N4713) );
  OR2X1 U16746 ( .IN2(n14719), .IN1(n14718), .Q(P2_N4693) );
  OR2X1 U16747 ( .IN2(n14721), .IN1(n14720), .Q(P2_N4694) );
  OR2X1 U16748 ( .IN2(n14723), .IN1(n14722), .Q(P2_N4695) );
  OR2X1 U16749 ( .IN2(n14725), .IN1(n14724), .Q(P2_N4696) );
  OR2X1 U16750 ( .IN2(n14727), .IN1(n14726), .Q(P2_N4697) );
  OR2X1 U16751 ( .IN2(n14729), .IN1(n14728), .Q(P2_N4698) );
  OR2X1 U16752 ( .IN2(n14731), .IN1(n14730), .Q(P2_N4699) );
  OR2X1 U16753 ( .IN2(n14733), .IN1(n14732), .Q(P2_N4700) );
  OR2X1 U16754 ( .IN2(n14735), .IN1(n14734), .Q(P2_N4701) );
  OR2X1 U16755 ( .IN2(n14737), .IN1(n14736), .Q(P2_N4702) );
  OR2X1 U16756 ( .IN2(n14739), .IN1(n14738), .Q(P2_N4703) );
  OR2X1 U16757 ( .IN2(n14741), .IN1(n14740), .Q(P2_N4704) );
  OR2X1 U16758 ( .IN2(n14743), .IN1(n14742), .Q(P2_N4705) );
  OR2X1 U16759 ( .IN2(n14745), .IN1(n14744), .Q(P2_N4706) );
  OR2X1 U16760 ( .IN2(n14747), .IN1(n14746), .Q(P2_N4707) );
  OR2X1 U16761 ( .IN2(n14749), .IN1(n14748), .Q(P2_N4708) );
  OR2X1 U16762 ( .IN2(n14751), .IN1(n14750), .Q(P2_N4709) );
  OR2X1 U16763 ( .IN2(n14753), .IN1(n14752), .Q(P2_N4710) );
  OR2X1 U16764 ( .IN2(n14755), .IN1(n14754), .Q(P2_N4711) );
  OR2X1 U16765 ( .IN2(n14757), .IN1(n14756), .Q(P2_N4712) );
  AND2X1 U16766 ( .IN1(n14759), .IN2(n6940), .Q(n14758) );
  OR2X1 U16767 ( .IN2(n14761), .IN1(n14760), .Q(P2_N4692) );
  AND2X1 U16768 ( .IN1(P2_N5059), .IN2(n6838), .Q(n14524) );
  AND2X1 U16769 ( .IN1(P2_N5062), .IN2(n6837), .Q(n14525) );
  OR2X1 U16584 ( .IN2(n14348), .IN1(n14346), .Q(n14359) );
  OR2X1 U16585 ( .IN2(n14351), .IN1(n14350), .Q(n14355) );
  OR2X1 U16586 ( .IN2(n14353), .IN1(n14352), .Q(n14357) );
  OR2X1 U16587 ( .IN2(n14356), .IN1(n14354), .Q(n14361) );
  OR2X1 U16588 ( .IN2(n14360), .IN1(n14358), .Q(n14370) );
  OR2X1 U16589 ( .IN2(n14363), .IN1(n14362), .Q(n14367) );
  OR2X1 U16590 ( .IN2(n14365), .IN1(n14364), .Q(n14369) );
  OR2X1 U16591 ( .IN2(n14368), .IN1(n14366), .Q(n14371) );
  OR2X1 U16592 ( .IN2(n14373), .IN1(n14372), .Q(n14377) );
  OR2X1 U16593 ( .IN2(n14375), .IN1(n14374), .Q(n14379) );
  OR2X1 U16594 ( .IN2(n14378), .IN1(n14376), .Q(n14389) );
  OR2X1 U16595 ( .IN2(n14381), .IN1(n14380), .Q(n14385) );
  OR2X1 U16596 ( .IN2(n14383), .IN1(n14382), .Q(n14387) );
  OR2X1 U16597 ( .IN2(n14386), .IN1(n14384), .Q(n14391) );
  OR2X1 U16598 ( .IN2(n14390), .IN1(n14388), .Q(n14400) );
  OR2X1 U16599 ( .IN2(n14393), .IN1(n14392), .Q(n14397) );
  OR2X1 U16600 ( .IN2(n14395), .IN1(n14394), .Q(n14399) );
  OR2X1 U16601 ( .IN2(n14398), .IN1(n14396), .Q(n14401) );
  OR2X1 U16602 ( .IN2(n14403), .IN1(n14402), .Q(n14407) );
  OR2X1 U16603 ( .IN2(n14405), .IN1(n14404), .Q(n14409) );
  OR2X1 U16604 ( .IN2(n14408), .IN1(n14406), .Q(n14419) );
  OR2X1 U16605 ( .IN2(n14411), .IN1(n14410), .Q(n14415) );
  OR2X1 U16606 ( .IN2(n14413), .IN1(n14412), .Q(n14417) );
  OR2X1 U16607 ( .IN2(n14416), .IN1(n14414), .Q(n14421) );
  OR2X1 U16608 ( .IN2(n14420), .IN1(n14418), .Q(n14430) );
  OR2X1 U16609 ( .IN2(n14423), .IN1(n14422), .Q(n14427) );
  OR2X1 U16610 ( .IN2(n14425), .IN1(n14424), .Q(n14429) );
  OR2X1 U16611 ( .IN2(n14428), .IN1(n14426), .Q(n14431) );
  OR2X1 U16612 ( .IN2(n14433), .IN1(n14432), .Q(n14437) );
  OR2X1 U16613 ( .IN2(n14435), .IN1(n14434), .Q(n14439) );
  OR2X1 U16614 ( .IN2(n14438), .IN1(n14436), .Q(n14449) );
  OR2X1 U16615 ( .IN2(n14441), .IN1(n14440), .Q(n14445) );
  OR2X1 U16616 ( .IN2(n14443), .IN1(n14442), .Q(n14447) );
  OR2X1 U16617 ( .IN2(n14446), .IN1(n14444), .Q(n14451) );
  OR2X1 U16618 ( .IN2(n14450), .IN1(n14448), .Q(n14460) );
  OR2X1 U16619 ( .IN2(n14453), .IN1(n14452), .Q(n14457) );
  OR2X1 U16620 ( .IN2(n14455), .IN1(n14454), .Q(n14459) );
  OR2X1 U16621 ( .IN2(n14458), .IN1(n14456), .Q(n14461) );
  OR2X1 U16622 ( .IN2(n14463), .IN1(n14462), .Q(n14467) );
  OR2X1 U16623 ( .IN2(n14465), .IN1(n14464), .Q(n14469) );
  OR2X1 U16624 ( .IN2(n14468), .IN1(n14466), .Q(n14479) );
  OR2X1 U16625 ( .IN2(n14471), .IN1(n14470), .Q(n14475) );
  OR2X1 U16626 ( .IN2(n14473), .IN1(n14472), .Q(n14477) );
  OR2X1 U16627 ( .IN2(n14476), .IN1(n14474), .Q(n14481) );
  OR2X1 U16628 ( .IN2(n14480), .IN1(n14478), .Q(n14490) );
  OR2X1 U16629 ( .IN2(n14483), .IN1(n14482), .Q(n14487) );
  OR2X1 U16630 ( .IN2(n14485), .IN1(n14484), .Q(n14489) );
  OR2X1 U16631 ( .IN2(n14488), .IN1(n14486), .Q(n14491) );
  OR2X1 U16632 ( .IN2(n14493), .IN1(n14492), .Q(n14497) );
  OR2X1 U16633 ( .IN2(n14495), .IN1(n14494), .Q(n14499) );
  OR2X1 U16634 ( .IN2(n14498), .IN1(n14496), .Q(n14509) );
  OR2X1 U16635 ( .IN2(n14501), .IN1(n14500), .Q(n14505) );
  OR2X1 U16636 ( .IN2(n14503), .IN1(n14502), .Q(n14507) );
  OR2X1 U16637 ( .IN2(n14506), .IN1(n14504), .Q(n14511) );
  OR2X1 U16638 ( .IN2(n14510), .IN1(n14508), .Q(n14520) );
  OR2X1 U16639 ( .IN2(n7019), .IN1(n6895), .Q(n14514) );
  OR2X1 U16640 ( .IN2(n6896), .IN1(n7019), .Q(n14513) );
  OR2X1 U16641 ( .IN2(n7019), .IN1(n6895), .Q(n14517) );
  OR2X1 U16642 ( .IN2(n6896), .IN1(n7019), .Q(n14516) );
  OR2X1 U16643 ( .IN2(n14512), .IN1(n6869), .Q(n14519) );
  OR2X1 U16644 ( .IN2(n14515), .IN1(n6870), .Q(n14518) );
  OR2X1 U16646 ( .IN2(n6813), .IN1(n7488), .Q(n14522) );
  OR2X1 U16647 ( .IN2(n14525), .IN1(n14524), .Q(n14523) );
  OR2X1 U16648 ( .IN2(n14527), .IN1(n14526), .Q(P2_N5355) );
  OR2X1 U16649 ( .IN2(n14529), .IN1(n14528), .Q(P2_N4810) );
  OR2X1 U16650 ( .IN2(n14531), .IN1(n14530), .Q(P2_N4811) );
  OR2X1 U16651 ( .IN2(n14533), .IN1(n14532), .Q(P2_N4812) );
  OR2X1 U16652 ( .IN2(n14535), .IN1(n14534), .Q(P2_N4813) );
  OR2X1 U16653 ( .IN2(n14537), .IN1(n14536), .Q(P2_N4814) );
  OR2X1 U16654 ( .IN2(n14539), .IN1(n14538), .Q(P2_N4815) );
  OR2X1 U16655 ( .IN2(n14541), .IN1(n14540), .Q(P2_N4816) );
  OR2X1 U16656 ( .IN2(n14543), .IN1(n14542), .Q(P2_N4817) );
  OR2X1 U16657 ( .IN2(n14545), .IN1(n14544), .Q(P2_N4818) );
  OR2X1 U16658 ( .IN2(n14547), .IN1(n14546), .Q(P2_N4819) );
  OR2X1 U16659 ( .IN2(n14549), .IN1(n14548), .Q(P2_N4820) );
  OR2X1 U16660 ( .IN2(n14551), .IN1(n14550), .Q(P2_N4821) );
  OR2X1 U16661 ( .IN2(n14553), .IN1(n14552), .Q(P2_N4822) );
  OR2X1 U16662 ( .IN2(n14555), .IN1(n14554), .Q(P2_N4823) );
  OR2X1 U16663 ( .IN2(n14557), .IN1(n14556), .Q(P2_N4824) );
  OR2X1 U16664 ( .IN2(n14559), .IN1(n14558), .Q(P2_N4825) );
  OR2X1 U16665 ( .IN2(n14561), .IN1(n14560), .Q(P2_N4826) );
  OR2X1 U16666 ( .IN2(n14563), .IN1(n14562), .Q(P2_N4827) );
  OR2X1 U16667 ( .IN2(n14565), .IN1(n14564), .Q(P2_N4828) );
  OR2X1 U16668 ( .IN2(n14567), .IN1(n14566), .Q(P2_N4829) );
  OR2X1 U16669 ( .IN2(n14569), .IN1(n14568), .Q(P2_N4830) );
  OR2X1 U16670 ( .IN2(n14571), .IN1(n14570), .Q(P2_N4831) );
  OR2X1 U16671 ( .IN2(n14573), .IN1(n14572), .Q(P2_N4832) );
  OR2X1 U16672 ( .IN2(n14575), .IN1(n14574), .Q(P2_N4833) );
  OR2X1 U16673 ( .IN2(n14577), .IN1(n14576), .Q(P2_N4834) );
  OR2X1 U16674 ( .IN2(n14579), .IN1(n14578), .Q(P2_N4835) );
  OR2X1 U16675 ( .IN2(n14581), .IN1(n14580), .Q(P2_N4836) );
  OR2X1 U16676 ( .IN2(n14583), .IN1(n14582), .Q(P2_N4837) );
  OR2X1 U16491 ( .IN2(n14068), .IN1(n14066), .Q(n14071) );
  OR2X1 U16492 ( .IN2(n14073), .IN1(n14072), .Q(n14077) );
  OR2X1 U16493 ( .IN2(n14075), .IN1(n14074), .Q(n14079) );
  OR2X1 U16494 ( .IN2(n14078), .IN1(n14076), .Q(n14089) );
  OR2X1 U16495 ( .IN2(n14081), .IN1(n14080), .Q(n14085) );
  OR2X1 U16496 ( .IN2(n14083), .IN1(n14082), .Q(n14087) );
  OR2X1 U16497 ( .IN2(n14086), .IN1(n14084), .Q(n14091) );
  OR2X1 U16498 ( .IN2(n14090), .IN1(n14088), .Q(n14100) );
  OR2X1 U16499 ( .IN2(n14093), .IN1(n14092), .Q(n14097) );
  OR2X1 U16500 ( .IN2(n14095), .IN1(n14094), .Q(n14099) );
  OR2X1 U16501 ( .IN2(n14098), .IN1(n14096), .Q(n14101) );
  OR2X1 U16502 ( .IN2(n14103), .IN1(n14102), .Q(n14107) );
  OR2X1 U16503 ( .IN2(n14105), .IN1(n14104), .Q(n14109) );
  OR2X1 U16504 ( .IN2(n14108), .IN1(n14106), .Q(n14119) );
  OR2X1 U16505 ( .IN2(n14111), .IN1(n14110), .Q(n14115) );
  OR2X1 U16506 ( .IN2(n14113), .IN1(n14112), .Q(n14117) );
  OR2X1 U16507 ( .IN2(n14116), .IN1(n14114), .Q(n14121) );
  OR2X1 U16508 ( .IN2(n14120), .IN1(n14118), .Q(n14130) );
  OR2X1 U16509 ( .IN2(n14123), .IN1(n14122), .Q(n14127) );
  OR2X1 U16510 ( .IN2(n14125), .IN1(n14124), .Q(n14129) );
  OR2X1 U16511 ( .IN2(n14128), .IN1(n14126), .Q(n14131) );
  OR2X1 U16512 ( .IN2(n14133), .IN1(n14132), .Q(n14137) );
  OR2X1 U16513 ( .IN2(n14135), .IN1(n14134), .Q(n14139) );
  OR2X1 U16514 ( .IN2(n14138), .IN1(n14136), .Q(n14149) );
  OR2X1 U16515 ( .IN2(n14141), .IN1(n14140), .Q(n14145) );
  OR2X1 U16516 ( .IN2(n14143), .IN1(n14142), .Q(n14147) );
  OR2X1 U16517 ( .IN2(n14146), .IN1(n14144), .Q(n14151) );
  OR2X1 U16518 ( .IN2(n14150), .IN1(n14148), .Q(n14160) );
  OR2X1 U16519 ( .IN2(n14153), .IN1(n14152), .Q(n14157) );
  OR2X1 U16520 ( .IN2(n14155), .IN1(n14154), .Q(n14159) );
  OR2X1 U16521 ( .IN2(n14158), .IN1(n14156), .Q(n14161) );
  OR2X1 U16522 ( .IN2(n14163), .IN1(n14162), .Q(n14167) );
  OR2X1 U16523 ( .IN2(n14165), .IN1(n14164), .Q(n14169) );
  OR2X1 U16524 ( .IN2(n14168), .IN1(n14166), .Q(n14179) );
  OR2X1 U16525 ( .IN2(n14171), .IN1(n14170), .Q(n14175) );
  OR2X1 U16526 ( .IN2(n14173), .IN1(n14172), .Q(n14177) );
  OR2X1 U16527 ( .IN2(n14176), .IN1(n14174), .Q(n14181) );
  OR2X1 U16528 ( .IN2(n14180), .IN1(n14178), .Q(n14190) );
  OR2X1 U16529 ( .IN2(n14183), .IN1(n14182), .Q(n14187) );
  OR2X1 U16530 ( .IN2(n14185), .IN1(n14184), .Q(n14189) );
  OR2X1 U16531 ( .IN2(n14188), .IN1(n14186), .Q(n14191) );
  OR2X1 U16532 ( .IN2(n14193), .IN1(n14192), .Q(n14197) );
  OR2X1 U16533 ( .IN2(n14195), .IN1(n14194), .Q(n14199) );
  OR2X1 U16534 ( .IN2(n14198), .IN1(n14196), .Q(n14209) );
  OR2X1 U16535 ( .IN2(n14201), .IN1(n14200), .Q(n14205) );
  OR2X1 U16536 ( .IN2(n14203), .IN1(n14202), .Q(n14207) );
  OR2X1 U16537 ( .IN2(n14206), .IN1(n14204), .Q(n14211) );
  OR2X1 U16538 ( .IN2(n14210), .IN1(n14208), .Q(n14220) );
  OR2X1 U16539 ( .IN2(n14213), .IN1(n14212), .Q(n14217) );
  OR2X1 U16540 ( .IN2(n14215), .IN1(n14214), .Q(n14219) );
  OR2X1 U16541 ( .IN2(n14218), .IN1(n14216), .Q(n14221) );
  OR2X1 U16542 ( .IN2(n14223), .IN1(n14222), .Q(n14227) );
  OR2X1 U16543 ( .IN2(n14225), .IN1(n14224), .Q(n14229) );
  OR2X1 U16544 ( .IN2(n14228), .IN1(n14226), .Q(n14239) );
  OR2X1 U16545 ( .IN2(n14231), .IN1(n14230), .Q(n14235) );
  OR2X1 U16546 ( .IN2(n14233), .IN1(n14232), .Q(n14237) );
  OR2X1 U16547 ( .IN2(n14236), .IN1(n14234), .Q(n14241) );
  OR2X1 U16548 ( .IN2(n14240), .IN1(n14238), .Q(n14250) );
  OR2X1 U16549 ( .IN2(n14243), .IN1(n14242), .Q(n14247) );
  OR2X1 U16550 ( .IN2(n14245), .IN1(n14244), .Q(n14249) );
  OR2X1 U16551 ( .IN2(n14248), .IN1(n14246), .Q(n14251) );
  OR2X1 U16552 ( .IN2(n14253), .IN1(n14252), .Q(n14257) );
  OR2X1 U16553 ( .IN2(n14255), .IN1(n14254), .Q(n14259) );
  OR2X1 U16554 ( .IN2(n14258), .IN1(n14256), .Q(n14269) );
  OR2X1 U16555 ( .IN2(n14261), .IN1(n14260), .Q(n14265) );
  OR2X1 U16556 ( .IN2(n14263), .IN1(n14262), .Q(n14267) );
  OR2X1 U16557 ( .IN2(n14266), .IN1(n14264), .Q(n14271) );
  OR2X1 U16558 ( .IN2(n14270), .IN1(n14268), .Q(n14280) );
  OR2X1 U16559 ( .IN2(n14273), .IN1(n14272), .Q(n14277) );
  OR2X1 U16560 ( .IN2(n14275), .IN1(n14274), .Q(n14279) );
  OR2X1 U16561 ( .IN2(n14278), .IN1(n14276), .Q(n14281) );
  OR2X1 U16562 ( .IN2(n14283), .IN1(n14282), .Q(n14287) );
  OR2X1 U16563 ( .IN2(n14285), .IN1(n14284), .Q(n14289) );
  OR2X1 U16564 ( .IN2(n14288), .IN1(n14286), .Q(n14299) );
  OR2X1 U16565 ( .IN2(n14291), .IN1(n14290), .Q(n14295) );
  OR2X1 U16566 ( .IN2(n14293), .IN1(n14292), .Q(n14297) );
  OR2X1 U16567 ( .IN2(n14296), .IN1(n14294), .Q(n14301) );
  OR2X1 U16568 ( .IN2(n14300), .IN1(n14298), .Q(n14310) );
  OR2X1 U16569 ( .IN2(n14303), .IN1(n14302), .Q(n14307) );
  OR2X1 U16570 ( .IN2(n14305), .IN1(n14304), .Q(n14309) );
  OR2X1 U16571 ( .IN2(n14308), .IN1(n14306), .Q(n14311) );
  OR2X1 U16572 ( .IN2(n14313), .IN1(n14312), .Q(n14317) );
  OR2X1 U16573 ( .IN2(n14315), .IN1(n14314), .Q(n14319) );
  OR2X1 U16574 ( .IN2(n14318), .IN1(n14316), .Q(n14329) );
  OR2X1 U16575 ( .IN2(n14321), .IN1(n14320), .Q(n14325) );
  OR2X1 U16576 ( .IN2(n14323), .IN1(n14322), .Q(n14327) );
  OR2X1 U16577 ( .IN2(n14326), .IN1(n14324), .Q(n14331) );
  OR2X1 U16578 ( .IN2(n14330), .IN1(n14328), .Q(n14340) );
  OR2X1 U16579 ( .IN2(n14333), .IN1(n14332), .Q(n14337) );
  OR2X1 U16580 ( .IN2(n14335), .IN1(n14334), .Q(n14339) );
  OR2X1 U16581 ( .IN2(n14338), .IN1(n14336), .Q(n14341) );
  OR2X1 U16582 ( .IN2(n14343), .IN1(n14342), .Q(n14347) );
  OR2X1 U16583 ( .IN2(n14345), .IN1(n14344), .Q(n14349) );
  OR2X1 U16398 ( .IN2(n13790), .IN1(n13789), .Q(n13793) );
  OR2X1 U16399 ( .IN2(n13792), .IN1(n13791), .Q(n13794) );
  OR2X1 U16400 ( .IN2(n13796), .IN1(n13795), .Q(n13799) );
  OR2X1 U16401 ( .IN2(n13798), .IN1(n13797), .Q(n13800) );
  OR2X1 U16402 ( .IN2(n13802), .IN1(n13801), .Q(n13804) );
  OR2X1 U16403 ( .IN2(n13805), .IN1(n13803), .Q(n13816) );
  OR2X1 U16404 ( .IN2(n13808), .IN1(n13807), .Q(n13812) );
  OR2X1 U16405 ( .IN2(n13810), .IN1(n13809), .Q(n13814) );
  OR2X1 U16406 ( .IN2(n13813), .IN1(n13811), .Q(n13818) );
  OR2X1 U16407 ( .IN2(n13817), .IN1(n13815), .Q(n13830) );
  OR2X1 U16408 ( .IN2(n13820), .IN1(n13819), .Q(n13824) );
  OR2X1 U16409 ( .IN2(n13822), .IN1(n13821), .Q(n13826) );
  OR2X1 U16410 ( .IN2(n13825), .IN1(n13823), .Q(n13828) );
  OR2X1 U16411 ( .IN2(n13829), .IN1(n13827), .Q(n13831) );
  OR2X1 U16412 ( .IN2(n13833), .IN1(n13832), .Q(n13835) );
  OR2X1 U16413 ( .IN2(n13836), .IN1(n13834), .Q(n13846) );
  OR2X1 U16414 ( .IN2(n13838), .IN1(n13837), .Q(n13842) );
  OR2X1 U16415 ( .IN2(n13840), .IN1(n13839), .Q(n13844) );
  OR2X1 U16416 ( .IN2(n13843), .IN1(n13841), .Q(n13848) );
  OR2X1 U16417 ( .IN2(n13847), .IN1(n13845), .Q(n13860) );
  OR2X1 U16418 ( .IN2(n13850), .IN1(n13849), .Q(n13854) );
  OR2X1 U16419 ( .IN2(n13852), .IN1(n13851), .Q(n13856) );
  OR2X1 U16420 ( .IN2(n13855), .IN1(n13853), .Q(n13858) );
  OR2X1 U16421 ( .IN2(n13859), .IN1(n13857), .Q(n13861) );
  OR2X1 U16422 ( .IN2(n13863), .IN1(n13862), .Q(n13865) );
  OR2X1 U16423 ( .IN2(n13866), .IN1(n13864), .Q(n13876) );
  OR2X1 U16424 ( .IN2(n13868), .IN1(n13867), .Q(n13872) );
  OR2X1 U16425 ( .IN2(n13870), .IN1(n13869), .Q(n13874) );
  OR2X1 U16426 ( .IN2(n13873), .IN1(n13871), .Q(n13878) );
  OR2X1 U16427 ( .IN2(n13877), .IN1(n13875), .Q(n13890) );
  OR2X1 U16428 ( .IN2(n13880), .IN1(n13879), .Q(n13884) );
  OR2X1 U16429 ( .IN2(n13882), .IN1(n13881), .Q(n13886) );
  OR2X1 U16430 ( .IN2(n13885), .IN1(n13883), .Q(n13888) );
  OR2X1 U16431 ( .IN2(n13889), .IN1(n13887), .Q(n13891) );
  OR2X1 U16432 ( .IN2(n13893), .IN1(n13892), .Q(n13897) );
  OR2X1 U16433 ( .IN2(n13895), .IN1(n13894), .Q(n13899) );
  OR2X1 U16434 ( .IN2(n13898), .IN1(n13896), .Q(n13909) );
  OR2X1 U16435 ( .IN2(n13901), .IN1(n13900), .Q(n13905) );
  OR2X1 U16436 ( .IN2(n13903), .IN1(n13902), .Q(n13907) );
  OR2X1 U16437 ( .IN2(n13906), .IN1(n13904), .Q(n13911) );
  OR2X1 U16438 ( .IN2(n13910), .IN1(n13908), .Q(n13920) );
  OR2X1 U16439 ( .IN2(n13913), .IN1(n13912), .Q(n13917) );
  OR2X1 U16440 ( .IN2(n13915), .IN1(n13914), .Q(n13919) );
  OR2X1 U16441 ( .IN2(n13918), .IN1(n13916), .Q(n13921) );
  OR2X1 U16442 ( .IN2(n13923), .IN1(n13922), .Q(n13927) );
  OR2X1 U16443 ( .IN2(n13925), .IN1(n13924), .Q(n13929) );
  OR2X1 U16444 ( .IN2(n13928), .IN1(n13926), .Q(n13939) );
  OR2X1 U16445 ( .IN2(n13931), .IN1(n13930), .Q(n13935) );
  OR2X1 U16446 ( .IN2(n13933), .IN1(n13932), .Q(n13937) );
  OR2X1 U16447 ( .IN2(n13936), .IN1(n13934), .Q(n13941) );
  OR2X1 U16448 ( .IN2(n13940), .IN1(n13938), .Q(n13950) );
  OR2X1 U16449 ( .IN2(n13943), .IN1(n13942), .Q(n13947) );
  OR2X1 U16450 ( .IN2(n13945), .IN1(n13944), .Q(n13949) );
  OR2X1 U16451 ( .IN2(n13948), .IN1(n13946), .Q(n13951) );
  OR2X1 U16452 ( .IN2(n13953), .IN1(n13952), .Q(n13957) );
  OR2X1 U16453 ( .IN2(n13955), .IN1(n13954), .Q(n13959) );
  OR2X1 U16454 ( .IN2(n13958), .IN1(n13956), .Q(n13969) );
  OR2X1 U16455 ( .IN2(n13961), .IN1(n13960), .Q(n13965) );
  OR2X1 U16456 ( .IN2(n13963), .IN1(n13962), .Q(n13967) );
  OR2X1 U16457 ( .IN2(n13966), .IN1(n13964), .Q(n13971) );
  OR2X1 U16458 ( .IN2(n13970), .IN1(n13968), .Q(n13980) );
  OR2X1 U16459 ( .IN2(n13973), .IN1(n13972), .Q(n13977) );
  OR2X1 U16460 ( .IN2(n13975), .IN1(n13974), .Q(n13979) );
  OR2X1 U16461 ( .IN2(n13978), .IN1(n13976), .Q(n13981) );
  OR2X1 U16462 ( .IN2(n13983), .IN1(n13982), .Q(n13987) );
  OR2X1 U16463 ( .IN2(n13985), .IN1(n13984), .Q(n13989) );
  OR2X1 U16464 ( .IN2(n13988), .IN1(n13986), .Q(n13999) );
  OR2X1 U16465 ( .IN2(n13991), .IN1(n13990), .Q(n13995) );
  OR2X1 U16466 ( .IN2(n13993), .IN1(n13992), .Q(n13997) );
  OR2X1 U16467 ( .IN2(n13996), .IN1(n13994), .Q(n14001) );
  OR2X1 U16468 ( .IN2(n14000), .IN1(n13998), .Q(n14010) );
  OR2X1 U16469 ( .IN2(n14003), .IN1(n14002), .Q(n14007) );
  OR2X1 U16470 ( .IN2(n14005), .IN1(n14004), .Q(n14009) );
  OR2X1 U16471 ( .IN2(n14008), .IN1(n14006), .Q(n14011) );
  OR2X1 U16472 ( .IN2(n14013), .IN1(n14012), .Q(n14017) );
  OR2X1 U16473 ( .IN2(n14015), .IN1(n14014), .Q(n14019) );
  OR2X1 U16474 ( .IN2(n14018), .IN1(n14016), .Q(n14029) );
  OR2X1 U16475 ( .IN2(n14021), .IN1(n14020), .Q(n14025) );
  OR2X1 U16476 ( .IN2(n14023), .IN1(n14022), .Q(n14027) );
  OR2X1 U16477 ( .IN2(n14026), .IN1(n14024), .Q(n14031) );
  OR2X1 U16478 ( .IN2(n14030), .IN1(n14028), .Q(n14040) );
  OR2X1 U16479 ( .IN2(n14033), .IN1(n14032), .Q(n14037) );
  OR2X1 U16480 ( .IN2(n14035), .IN1(n14034), .Q(n14039) );
  OR2X1 U16481 ( .IN2(n14038), .IN1(n14036), .Q(n14041) );
  OR2X1 U16482 ( .IN2(n14043), .IN1(n14042), .Q(n14047) );
  OR2X1 U16483 ( .IN2(n14045), .IN1(n14044), .Q(n14049) );
  OR2X1 U16484 ( .IN2(n14048), .IN1(n14046), .Q(n14059) );
  OR2X1 U16485 ( .IN2(n14051), .IN1(n14050), .Q(n14055) );
  OR2X1 U16486 ( .IN2(n14053), .IN1(n14052), .Q(n14057) );
  OR2X1 U16487 ( .IN2(n14056), .IN1(n14054), .Q(n14061) );
  OR2X1 U16488 ( .IN2(n14060), .IN1(n14058), .Q(n14070) );
  OR2X1 U16489 ( .IN2(n14063), .IN1(n14062), .Q(n14067) );
  OR2X1 U16490 ( .IN2(n14065), .IN1(n14064), .Q(n14069) );
  OR2X1 U16305 ( .IN2(n13510), .IN1(n13509), .Q(n13514) );
  OR2X1 U16306 ( .IN2(n13512), .IN1(n13511), .Q(n13516) );
  OR2X1 U16307 ( .IN2(n13515), .IN1(n13513), .Q(n13519) );
  OR2X1 U16308 ( .IN2(n13518), .IN1(n13517), .Q(n13521) );
  OR2X1 U16309 ( .IN2(n13523), .IN1(n13522), .Q(n13527) );
  OR2X1 U16310 ( .IN2(n13525), .IN1(n13524), .Q(n13529) );
  OR2X1 U16311 ( .IN2(n13528), .IN1(n13526), .Q(n13539) );
  OR2X1 U16312 ( .IN2(n13531), .IN1(n13530), .Q(n13535) );
  OR2X1 U16313 ( .IN2(n13533), .IN1(n13532), .Q(n13537) );
  OR2X1 U16314 ( .IN2(n13536), .IN1(n13534), .Q(n13541) );
  OR2X1 U16315 ( .IN2(n13540), .IN1(n13538), .Q(n13553) );
  OR2X1 U16316 ( .IN2(n13543), .IN1(n13542), .Q(n13547) );
  OR2X1 U16317 ( .IN2(n13545), .IN1(n13544), .Q(n13549) );
  OR2X1 U16318 ( .IN2(n13548), .IN1(n13546), .Q(n13552) );
  OR2X1 U16319 ( .IN2(n13551), .IN1(n13550), .Q(n13554) );
  OR2X1 U16320 ( .IN2(n13556), .IN1(n13555), .Q(n13560) );
  OR2X1 U16321 ( .IN2(n13558), .IN1(n13557), .Q(n13562) );
  OR2X1 U16322 ( .IN2(n13561), .IN1(n13559), .Q(n13572) );
  OR2X1 U16323 ( .IN2(n13564), .IN1(n13563), .Q(n13568) );
  OR2X1 U16324 ( .IN2(n13566), .IN1(n13565), .Q(n13570) );
  OR2X1 U16325 ( .IN2(n13569), .IN1(n13567), .Q(n13574) );
  OR2X1 U16326 ( .IN2(n13573), .IN1(n13571), .Q(n13586) );
  OR2X1 U16327 ( .IN2(n13576), .IN1(n13575), .Q(n13580) );
  OR2X1 U16328 ( .IN2(n13578), .IN1(n13577), .Q(n13582) );
  OR2X1 U16329 ( .IN2(n13581), .IN1(n13579), .Q(n13585) );
  OR2X1 U16330 ( .IN2(n13584), .IN1(n13583), .Q(n13587) );
  OR2X1 U16331 ( .IN2(n13589), .IN1(n13588), .Q(n13593) );
  OR2X1 U16332 ( .IN2(n13591), .IN1(n13590), .Q(n13595) );
  OR2X1 U16333 ( .IN2(n13594), .IN1(n13592), .Q(n13605) );
  OR2X1 U16334 ( .IN2(n13597), .IN1(n13596), .Q(n13601) );
  OR2X1 U16335 ( .IN2(n13599), .IN1(n13598), .Q(n13603) );
  OR2X1 U16336 ( .IN2(n13602), .IN1(n13600), .Q(n13607) );
  OR2X1 U16337 ( .IN2(n13606), .IN1(n13604), .Q(n13619) );
  OR2X1 U16338 ( .IN2(n13609), .IN1(n13608), .Q(n13613) );
  OR2X1 U16339 ( .IN2(n13611), .IN1(n13610), .Q(n13615) );
  OR2X1 U16340 ( .IN2(n13614), .IN1(n13612), .Q(n13618) );
  OR2X1 U16341 ( .IN2(n13617), .IN1(n13616), .Q(n13620) );
  OR2X1 U16342 ( .IN2(n13622), .IN1(n13621), .Q(n13625) );
  OR2X1 U16343 ( .IN2(n13624), .IN1(n13623), .Q(n13626) );
  OR2X1 U16344 ( .IN2(n13628), .IN1(n13627), .Q(n13631) );
  OR2X1 U16345 ( .IN2(n13630), .IN1(n13629), .Q(n13632) );
  OR2X1 U16346 ( .IN2(n13634), .IN1(n13633), .Q(n13637) );
  OR2X1 U16347 ( .IN2(n13636), .IN1(n13635), .Q(n13638) );
  OR2X1 U16348 ( .IN2(n13640), .IN1(n13639), .Q(n13643) );
  OR2X1 U16349 ( .IN2(n13642), .IN1(n13641), .Q(n13644) );
  OR2X1 U16350 ( .IN2(n13646), .IN1(n13645), .Q(n13649) );
  OR2X1 U16351 ( .IN2(n13648), .IN1(n13647), .Q(n13650) );
  OR2X1 U16352 ( .IN2(n13652), .IN1(n13651), .Q(n13655) );
  OR2X1 U16353 ( .IN2(n13654), .IN1(n13653), .Q(n13656) );
  OR2X1 U16354 ( .IN2(n13658), .IN1(n13657), .Q(n13661) );
  OR2X1 U16355 ( .IN2(n13660), .IN1(n13659), .Q(n13662) );
  OR2X1 U16356 ( .IN2(n13664), .IN1(n13663), .Q(n13667) );
  OR2X1 U16357 ( .IN2(n13666), .IN1(n13665), .Q(n13668) );
  OR2X1 U16358 ( .IN2(n13670), .IN1(n13669), .Q(n13673) );
  OR2X1 U16359 ( .IN2(n13672), .IN1(n13671), .Q(n13674) );
  OR2X1 U16360 ( .IN2(n13676), .IN1(n13675), .Q(n13679) );
  OR2X1 U16361 ( .IN2(n13678), .IN1(n13677), .Q(n13680) );
  OR2X1 U16362 ( .IN2(n13682), .IN1(n13681), .Q(n13685) );
  OR2X1 U16363 ( .IN2(n13684), .IN1(n13683), .Q(n13686) );
  OR2X1 U16364 ( .IN2(n13688), .IN1(n13687), .Q(n13691) );
  OR2X1 U16365 ( .IN2(n13690), .IN1(n13689), .Q(n13692) );
  OR2X1 U16366 ( .IN2(n13694), .IN1(n13693), .Q(n13697) );
  OR2X1 U16367 ( .IN2(n13696), .IN1(n13695), .Q(n13698) );
  OR2X1 U16368 ( .IN2(n13700), .IN1(n13699), .Q(n13703) );
  OR2X1 U16369 ( .IN2(n13702), .IN1(n13701), .Q(n13704) );
  OR2X1 U16370 ( .IN2(n13706), .IN1(n13705), .Q(n13709) );
  OR2X1 U16371 ( .IN2(n13708), .IN1(n13707), .Q(n13710) );
  OR2X1 U16372 ( .IN2(n13712), .IN1(n13711), .Q(n13715) );
  OR2X1 U16373 ( .IN2(n13714), .IN1(n13713), .Q(n13716) );
  OR2X1 U16374 ( .IN2(n13718), .IN1(n13717), .Q(n13721) );
  OR2X1 U16375 ( .IN2(n13720), .IN1(n13719), .Q(n13722) );
  OR2X1 U16376 ( .IN2(n13724), .IN1(n13723), .Q(n13727) );
  OR2X1 U16377 ( .IN2(n13726), .IN1(n13725), .Q(n13728) );
  OR2X1 U16378 ( .IN2(n13730), .IN1(n13729), .Q(n13733) );
  OR2X1 U16379 ( .IN2(n13732), .IN1(n13731), .Q(n13734) );
  OR2X1 U16380 ( .IN2(n13736), .IN1(n13735), .Q(n13739) );
  OR2X1 U16381 ( .IN2(n13738), .IN1(n13737), .Q(n13740) );
  OR2X1 U16382 ( .IN2(n13742), .IN1(n13741), .Q(n13745) );
  OR2X1 U16383 ( .IN2(n13744), .IN1(n13743), .Q(n13746) );
  OR2X1 U16384 ( .IN2(n13748), .IN1(n13747), .Q(n13751) );
  OR2X1 U16385 ( .IN2(n13750), .IN1(n13749), .Q(n13752) );
  OR2X1 U16386 ( .IN2(n13754), .IN1(n13753), .Q(n13757) );
  OR2X1 U16387 ( .IN2(n13756), .IN1(n13755), .Q(n13758) );
  OR2X1 U16388 ( .IN2(n13760), .IN1(n13759), .Q(n13763) );
  OR2X1 U16389 ( .IN2(n13762), .IN1(n13761), .Q(n13764) );
  OR2X1 U16390 ( .IN2(n13766), .IN1(n13765), .Q(n13769) );
  OR2X1 U16391 ( .IN2(n13768), .IN1(n13767), .Q(n13770) );
  OR2X1 U16392 ( .IN2(n13772), .IN1(n13771), .Q(n13775) );
  OR2X1 U16393 ( .IN2(n13774), .IN1(n13773), .Q(n13776) );
  OR2X1 U16394 ( .IN2(n13778), .IN1(n13777), .Q(n13781) );
  OR2X1 U16395 ( .IN2(n13780), .IN1(n13779), .Q(n13782) );
  OR2X1 U16396 ( .IN2(n13784), .IN1(n13783), .Q(n13787) );
  OR2X1 U16397 ( .IN2(n13786), .IN1(n13785), .Q(n13788) );
  OR2X1 U16212 ( .IN2(n13231), .IN1(n13229), .Q(n13242) );
  OR2X1 U16213 ( .IN2(n13234), .IN1(n13233), .Q(n13238) );
  OR2X1 U16214 ( .IN2(n13236), .IN1(n13235), .Q(n13240) );
  OR2X1 U16215 ( .IN2(n13239), .IN1(n13237), .Q(n13244) );
  OR2X1 U16216 ( .IN2(n13243), .IN1(n13241), .Q(n13256) );
  OR2X1 U16217 ( .IN2(n13246), .IN1(n13245), .Q(n13250) );
  OR2X1 U16218 ( .IN2(n13248), .IN1(n13247), .Q(n13252) );
  OR2X1 U16219 ( .IN2(n13251), .IN1(n13249), .Q(n13255) );
  OR2X1 U16220 ( .IN2(n13254), .IN1(n13253), .Q(n13257) );
  OR2X1 U16221 ( .IN2(n13259), .IN1(n13258), .Q(n13263) );
  OR2X1 U16222 ( .IN2(n13261), .IN1(n13260), .Q(n13265) );
  OR2X1 U16223 ( .IN2(n13264), .IN1(n13262), .Q(n13275) );
  OR2X1 U16224 ( .IN2(n13267), .IN1(n13266), .Q(n13271) );
  OR2X1 U16225 ( .IN2(n13269), .IN1(n13268), .Q(n13273) );
  OR2X1 U16226 ( .IN2(n13272), .IN1(n13270), .Q(n13277) );
  OR2X1 U16227 ( .IN2(n13276), .IN1(n13274), .Q(n13289) );
  OR2X1 U16228 ( .IN2(n13279), .IN1(n13278), .Q(n13283) );
  OR2X1 U16229 ( .IN2(n13281), .IN1(n13280), .Q(n13285) );
  OR2X1 U16230 ( .IN2(n13284), .IN1(n13282), .Q(n13288) );
  OR2X1 U16231 ( .IN2(n13287), .IN1(n13286), .Q(n13290) );
  OR2X1 U16232 ( .IN2(n13292), .IN1(n13291), .Q(n13296) );
  OR2X1 U16233 ( .IN2(n13294), .IN1(n13293), .Q(n13298) );
  OR2X1 U16234 ( .IN2(n13297), .IN1(n13295), .Q(n13308) );
  OR2X1 U16235 ( .IN2(n13300), .IN1(n13299), .Q(n13304) );
  OR2X1 U16236 ( .IN2(n13302), .IN1(n13301), .Q(n13306) );
  OR2X1 U16237 ( .IN2(n13305), .IN1(n13303), .Q(n13310) );
  OR2X1 U16238 ( .IN2(n13309), .IN1(n13307), .Q(n13322) );
  OR2X1 U16239 ( .IN2(n13312), .IN1(n13311), .Q(n13316) );
  OR2X1 U16240 ( .IN2(n13314), .IN1(n13313), .Q(n13318) );
  OR2X1 U16241 ( .IN2(n13317), .IN1(n13315), .Q(n13321) );
  OR2X1 U16242 ( .IN2(n13320), .IN1(n13319), .Q(n13323) );
  OR2X1 U16243 ( .IN2(n13325), .IN1(n13324), .Q(n13329) );
  OR2X1 U16244 ( .IN2(n13327), .IN1(n13326), .Q(n13331) );
  OR2X1 U16245 ( .IN2(n13330), .IN1(n13328), .Q(n13341) );
  OR2X1 U16246 ( .IN2(n13333), .IN1(n13332), .Q(n13337) );
  OR2X1 U16247 ( .IN2(n13335), .IN1(n13334), .Q(n13339) );
  OR2X1 U16248 ( .IN2(n13338), .IN1(n13336), .Q(n13343) );
  OR2X1 U16249 ( .IN2(n13342), .IN1(n13340), .Q(n13355) );
  OR2X1 U16250 ( .IN2(n13345), .IN1(n13344), .Q(n13349) );
  OR2X1 U16251 ( .IN2(n13347), .IN1(n13346), .Q(n13351) );
  OR2X1 U16252 ( .IN2(n13350), .IN1(n13348), .Q(n13354) );
  OR2X1 U16253 ( .IN2(n13353), .IN1(n13352), .Q(n13356) );
  OR2X1 U16254 ( .IN2(n13358), .IN1(n13357), .Q(n13362) );
  OR2X1 U16255 ( .IN2(n13360), .IN1(n13359), .Q(n13364) );
  OR2X1 U16256 ( .IN2(n13363), .IN1(n13361), .Q(n13374) );
  OR2X1 U16257 ( .IN2(n13366), .IN1(n13365), .Q(n13370) );
  OR2X1 U16258 ( .IN2(n13368), .IN1(n13367), .Q(n13372) );
  OR2X1 U16259 ( .IN2(n13371), .IN1(n13369), .Q(n13376) );
  OR2X1 U16260 ( .IN2(n13375), .IN1(n13373), .Q(n13388) );
  OR2X1 U16261 ( .IN2(n13378), .IN1(n13377), .Q(n13382) );
  OR2X1 U16262 ( .IN2(n13380), .IN1(n13379), .Q(n13384) );
  OR2X1 U16263 ( .IN2(n13383), .IN1(n13381), .Q(n13387) );
  OR2X1 U16264 ( .IN2(n13386), .IN1(n13385), .Q(n13389) );
  OR2X1 U16265 ( .IN2(n13391), .IN1(n13390), .Q(n13395) );
  OR2X1 U16266 ( .IN2(n13393), .IN1(n13392), .Q(n13397) );
  OR2X1 U16267 ( .IN2(n13396), .IN1(n13394), .Q(n13407) );
  OR2X1 U16268 ( .IN2(n13399), .IN1(n13398), .Q(n13403) );
  OR2X1 U16269 ( .IN2(n13401), .IN1(n13400), .Q(n13405) );
  OR2X1 U16270 ( .IN2(n13404), .IN1(n13402), .Q(n13409) );
  OR2X1 U16271 ( .IN2(n13408), .IN1(n13406), .Q(n13421) );
  OR2X1 U16272 ( .IN2(n13411), .IN1(n13410), .Q(n13415) );
  OR2X1 U16273 ( .IN2(n13413), .IN1(n13412), .Q(n13417) );
  OR2X1 U16274 ( .IN2(n13416), .IN1(n13414), .Q(n13420) );
  OR2X1 U16275 ( .IN2(n13419), .IN1(n13418), .Q(n13422) );
  OR2X1 U16276 ( .IN2(n13424), .IN1(n13423), .Q(n13428) );
  OR2X1 U16277 ( .IN2(n13426), .IN1(n13425), .Q(n13430) );
  OR2X1 U16278 ( .IN2(n13429), .IN1(n13427), .Q(n13440) );
  OR2X1 U16279 ( .IN2(n13432), .IN1(n13431), .Q(n13436) );
  OR2X1 U16280 ( .IN2(n13434), .IN1(n13433), .Q(n13438) );
  OR2X1 U16281 ( .IN2(n13437), .IN1(n13435), .Q(n13442) );
  OR2X1 U16282 ( .IN2(n13441), .IN1(n13439), .Q(n13454) );
  OR2X1 U16283 ( .IN2(n13444), .IN1(n13443), .Q(n13448) );
  OR2X1 U16284 ( .IN2(n13446), .IN1(n13445), .Q(n13450) );
  OR2X1 U16285 ( .IN2(n13449), .IN1(n13447), .Q(n13453) );
  OR2X1 U16286 ( .IN2(n13452), .IN1(n13451), .Q(n13455) );
  OR2X1 U16287 ( .IN2(n13457), .IN1(n13456), .Q(n13461) );
  OR2X1 U16288 ( .IN2(n13459), .IN1(n13458), .Q(n13463) );
  OR2X1 U16289 ( .IN2(n13462), .IN1(n13460), .Q(n13473) );
  OR2X1 U16290 ( .IN2(n13465), .IN1(n13464), .Q(n13469) );
  OR2X1 U16291 ( .IN2(n13467), .IN1(n13466), .Q(n13471) );
  OR2X1 U16292 ( .IN2(n13470), .IN1(n13468), .Q(n13475) );
  OR2X1 U16293 ( .IN2(n13474), .IN1(n13472), .Q(n13487) );
  OR2X1 U16294 ( .IN2(n13477), .IN1(n13476), .Q(n13481) );
  OR2X1 U16295 ( .IN2(n13479), .IN1(n13478), .Q(n13483) );
  OR2X1 U16296 ( .IN2(n13482), .IN1(n13480), .Q(n13486) );
  OR2X1 U16297 ( .IN2(n13485), .IN1(n13484), .Q(n13488) );
  OR2X1 U16298 ( .IN2(n13490), .IN1(n13489), .Q(n13494) );
  OR2X1 U16299 ( .IN2(n13492), .IN1(n13491), .Q(n13496) );
  OR2X1 U16300 ( .IN2(n13495), .IN1(n13493), .Q(n13506) );
  OR2X1 U16301 ( .IN2(n13498), .IN1(n13497), .Q(n13502) );
  OR2X1 U16302 ( .IN2(n13500), .IN1(n13499), .Q(n13504) );
  OR2X1 U16303 ( .IN2(n13503), .IN1(n13501), .Q(n13508) );
  OR2X1 U16304 ( .IN2(n13507), .IN1(n13505), .Q(n13520) );
  OR2X1 U16119 ( .IN2(n12951), .IN1(n12950), .Q(n12955) );
  OR2X1 U16120 ( .IN2(n12954), .IN1(n12952), .Q(n12958) );
  OR2X1 U16121 ( .IN2(n12957), .IN1(n12956), .Q(n12960) );
  OR2X1 U16122 ( .IN2(n12962), .IN1(n12961), .Q(n12966) );
  OR2X1 U16123 ( .IN2(n12964), .IN1(n12963), .Q(n12968) );
  OR2X1 U16124 ( .IN2(n12967), .IN1(n12965), .Q(n12978) );
  OR2X1 U16125 ( .IN2(n12970), .IN1(n12969), .Q(n12974) );
  OR2X1 U16126 ( .IN2(n12972), .IN1(n12971), .Q(n12976) );
  OR2X1 U16127 ( .IN2(n12975), .IN1(n12973), .Q(n12980) );
  OR2X1 U16128 ( .IN2(n12979), .IN1(n12977), .Q(n12992) );
  OR2X1 U16129 ( .IN2(n12982), .IN1(n12981), .Q(n12986) );
  OR2X1 U16130 ( .IN2(n12984), .IN1(n12983), .Q(n12988) );
  OR2X1 U16131 ( .IN2(n12987), .IN1(n12985), .Q(n12991) );
  OR2X1 U16132 ( .IN2(n12990), .IN1(n12989), .Q(n12993) );
  OR2X1 U16133 ( .IN2(n12995), .IN1(n12994), .Q(n12999) );
  OR2X1 U16134 ( .IN2(n12997), .IN1(n12996), .Q(n13001) );
  OR2X1 U16135 ( .IN2(n13000), .IN1(n12998), .Q(n13011) );
  OR2X1 U16136 ( .IN2(n13003), .IN1(n13002), .Q(n13007) );
  OR2X1 U16137 ( .IN2(n13005), .IN1(n13004), .Q(n13009) );
  OR2X1 U16138 ( .IN2(n13008), .IN1(n13006), .Q(n13013) );
  OR2X1 U16139 ( .IN2(n13012), .IN1(n13010), .Q(n13025) );
  OR2X1 U16140 ( .IN2(n13015), .IN1(n13014), .Q(n13019) );
  OR2X1 U16141 ( .IN2(n13017), .IN1(n13016), .Q(n13021) );
  OR2X1 U16142 ( .IN2(n13020), .IN1(n13018), .Q(n13024) );
  OR2X1 U16143 ( .IN2(n13023), .IN1(n13022), .Q(n13026) );
  OR2X1 U16144 ( .IN2(n13028), .IN1(n13027), .Q(n13032) );
  OR2X1 U16145 ( .IN2(n13030), .IN1(n13029), .Q(n13034) );
  OR2X1 U16146 ( .IN2(n13033), .IN1(n13031), .Q(n13044) );
  OR2X1 U16147 ( .IN2(n13036), .IN1(n13035), .Q(n13040) );
  OR2X1 U16148 ( .IN2(n13038), .IN1(n13037), .Q(n13042) );
  OR2X1 U16149 ( .IN2(n13041), .IN1(n13039), .Q(n13046) );
  OR2X1 U16150 ( .IN2(n13045), .IN1(n13043), .Q(n13058) );
  OR2X1 U16151 ( .IN2(n13048), .IN1(n13047), .Q(n13052) );
  OR2X1 U16152 ( .IN2(n13050), .IN1(n13049), .Q(n13054) );
  OR2X1 U16153 ( .IN2(n13053), .IN1(n13051), .Q(n13057) );
  OR2X1 U16154 ( .IN2(n13056), .IN1(n13055), .Q(n13059) );
  OR2X1 U16155 ( .IN2(n13061), .IN1(n13060), .Q(n13065) );
  OR2X1 U16156 ( .IN2(n13063), .IN1(n13062), .Q(n13067) );
  OR2X1 U16157 ( .IN2(n13066), .IN1(n13064), .Q(n13077) );
  OR2X1 U16158 ( .IN2(n13069), .IN1(n13068), .Q(n13073) );
  OR2X1 U16159 ( .IN2(n13071), .IN1(n13070), .Q(n13075) );
  OR2X1 U16160 ( .IN2(n13074), .IN1(n13072), .Q(n13079) );
  OR2X1 U16161 ( .IN2(n13078), .IN1(n13076), .Q(n13091) );
  OR2X1 U16162 ( .IN2(n13081), .IN1(n13080), .Q(n13085) );
  OR2X1 U16163 ( .IN2(n13083), .IN1(n13082), .Q(n13087) );
  OR2X1 U16164 ( .IN2(n13086), .IN1(n13084), .Q(n13090) );
  OR2X1 U16165 ( .IN2(n13089), .IN1(n13088), .Q(n13092) );
  OR2X1 U16166 ( .IN2(n13094), .IN1(n13093), .Q(n13098) );
  OR2X1 U16167 ( .IN2(n13096), .IN1(n13095), .Q(n13100) );
  OR2X1 U16168 ( .IN2(n13099), .IN1(n13097), .Q(n13110) );
  OR2X1 U16169 ( .IN2(n13102), .IN1(n13101), .Q(n13106) );
  OR2X1 U16170 ( .IN2(n13104), .IN1(n13103), .Q(n13108) );
  OR2X1 U16171 ( .IN2(n13107), .IN1(n13105), .Q(n13112) );
  OR2X1 U16172 ( .IN2(n13111), .IN1(n13109), .Q(n13124) );
  OR2X1 U16173 ( .IN2(n13114), .IN1(n13113), .Q(n13118) );
  OR2X1 U16174 ( .IN2(n13116), .IN1(n13115), .Q(n13120) );
  OR2X1 U16175 ( .IN2(n13119), .IN1(n13117), .Q(n13123) );
  OR2X1 U16176 ( .IN2(n13122), .IN1(n13121), .Q(n13125) );
  OR2X1 U16177 ( .IN2(n13127), .IN1(n13126), .Q(n13131) );
  OR2X1 U16178 ( .IN2(n13129), .IN1(n13128), .Q(n13133) );
  OR2X1 U16179 ( .IN2(n13132), .IN1(n13130), .Q(n13143) );
  OR2X1 U16180 ( .IN2(n13135), .IN1(n13134), .Q(n13139) );
  OR2X1 U16181 ( .IN2(n13137), .IN1(n13136), .Q(n13141) );
  OR2X1 U16182 ( .IN2(n13140), .IN1(n13138), .Q(n13145) );
  OR2X1 U16183 ( .IN2(n13144), .IN1(n13142), .Q(n13157) );
  OR2X1 U16184 ( .IN2(n13147), .IN1(n13146), .Q(n13151) );
  OR2X1 U16185 ( .IN2(n13149), .IN1(n13148), .Q(n13153) );
  OR2X1 U16186 ( .IN2(n13152), .IN1(n13150), .Q(n13156) );
  OR2X1 U16187 ( .IN2(n13155), .IN1(n13154), .Q(n13158) );
  OR2X1 U16188 ( .IN2(n13160), .IN1(n13159), .Q(n13164) );
  OR2X1 U16189 ( .IN2(n13162), .IN1(n13161), .Q(n13166) );
  OR2X1 U16190 ( .IN2(n13165), .IN1(n13163), .Q(n13176) );
  OR2X1 U16191 ( .IN2(n13168), .IN1(n13167), .Q(n13172) );
  OR2X1 U16192 ( .IN2(n13170), .IN1(n13169), .Q(n13174) );
  OR2X1 U16193 ( .IN2(n13173), .IN1(n13171), .Q(n13178) );
  OR2X1 U16194 ( .IN2(n13177), .IN1(n13175), .Q(n13190) );
  OR2X1 U16195 ( .IN2(n13180), .IN1(n13179), .Q(n13184) );
  OR2X1 U16196 ( .IN2(n13182), .IN1(n13181), .Q(n13186) );
  OR2X1 U16197 ( .IN2(n13185), .IN1(n13183), .Q(n13189) );
  OR2X1 U16198 ( .IN2(n13188), .IN1(n13187), .Q(n13191) );
  OR2X1 U16199 ( .IN2(n13193), .IN1(n13192), .Q(n13197) );
  OR2X1 U16200 ( .IN2(n13195), .IN1(n13194), .Q(n13199) );
  OR2X1 U16201 ( .IN2(n13198), .IN1(n13196), .Q(n13209) );
  OR2X1 U16202 ( .IN2(n13201), .IN1(n13200), .Q(n13205) );
  OR2X1 U16203 ( .IN2(n13203), .IN1(n13202), .Q(n13207) );
  OR2X1 U16204 ( .IN2(n13206), .IN1(n13204), .Q(n13211) );
  OR2X1 U16205 ( .IN2(n13210), .IN1(n13208), .Q(n13223) );
  OR2X1 U16206 ( .IN2(n13213), .IN1(n13212), .Q(n13217) );
  OR2X1 U16207 ( .IN2(n13215), .IN1(n13214), .Q(n13219) );
  OR2X1 U16208 ( .IN2(n13218), .IN1(n13216), .Q(n13222) );
  OR2X1 U16209 ( .IN2(n13221), .IN1(n13220), .Q(n13224) );
  OR2X1 U16210 ( .IN2(n13226), .IN1(n13225), .Q(n13230) );
  OR2X1 U16211 ( .IN2(n13228), .IN1(n13227), .Q(n13232) );
  OR2X1 U16026 ( .IN2(n12673), .IN1(n12672), .Q(n12677) );
  OR2X1 U16027 ( .IN2(n12675), .IN1(n12674), .Q(n12679) );
  OR2X1 U16028 ( .IN2(n12678), .IN1(n12676), .Q(n12683) );
  OR2X1 U16029 ( .IN2(n12682), .IN1(n12680), .Q(n12695) );
  OR2X1 U16030 ( .IN2(n12685), .IN1(n12684), .Q(n12689) );
  OR2X1 U16031 ( .IN2(n12687), .IN1(n12686), .Q(n12691) );
  OR2X1 U16032 ( .IN2(n12690), .IN1(n12688), .Q(n12694) );
  OR2X1 U16033 ( .IN2(n12693), .IN1(n12692), .Q(n12696) );
  OR2X1 U16034 ( .IN2(n12698), .IN1(n12697), .Q(n12702) );
  OR2X1 U16035 ( .IN2(n12700), .IN1(n12699), .Q(n12704) );
  OR2X1 U16036 ( .IN2(n12703), .IN1(n12701), .Q(n12714) );
  OR2X1 U16037 ( .IN2(n12706), .IN1(n12705), .Q(n12710) );
  OR2X1 U16038 ( .IN2(n12708), .IN1(n12707), .Q(n12712) );
  OR2X1 U16039 ( .IN2(n12711), .IN1(n12709), .Q(n12716) );
  OR2X1 U16040 ( .IN2(n12715), .IN1(n12713), .Q(n12728) );
  OR2X1 U16041 ( .IN2(n12718), .IN1(n12717), .Q(n12722) );
  OR2X1 U16042 ( .IN2(n12720), .IN1(n12719), .Q(n12724) );
  OR2X1 U16043 ( .IN2(n12723), .IN1(n12721), .Q(n12727) );
  OR2X1 U16044 ( .IN2(n12726), .IN1(n12725), .Q(n12729) );
  OR2X1 U16045 ( .IN2(n12731), .IN1(n12730), .Q(n12735) );
  OR2X1 U16046 ( .IN2(n12733), .IN1(n12732), .Q(n12737) );
  OR2X1 U16047 ( .IN2(n12736), .IN1(n12734), .Q(n12747) );
  OR2X1 U16048 ( .IN2(n12739), .IN1(n12738), .Q(n12743) );
  OR2X1 U16049 ( .IN2(n12741), .IN1(n12740), .Q(n12745) );
  OR2X1 U16050 ( .IN2(n12744), .IN1(n12742), .Q(n12749) );
  OR2X1 U16051 ( .IN2(n12748), .IN1(n12746), .Q(n12761) );
  OR2X1 U16052 ( .IN2(n12751), .IN1(n12750), .Q(n12755) );
  OR2X1 U16053 ( .IN2(n12753), .IN1(n12752), .Q(n12757) );
  OR2X1 U16054 ( .IN2(n12756), .IN1(n12754), .Q(n12760) );
  OR2X1 U16055 ( .IN2(n12759), .IN1(n12758), .Q(n12762) );
  OR2X1 U16056 ( .IN2(n12764), .IN1(n12763), .Q(n12768) );
  OR2X1 U16057 ( .IN2(n12766), .IN1(n12765), .Q(n12770) );
  OR2X1 U16058 ( .IN2(n12769), .IN1(n12767), .Q(n12780) );
  OR2X1 U16059 ( .IN2(n12772), .IN1(n12771), .Q(n12776) );
  OR2X1 U16060 ( .IN2(n12774), .IN1(n12773), .Q(n12778) );
  OR2X1 U16061 ( .IN2(n12777), .IN1(n12775), .Q(n12782) );
  OR2X1 U16062 ( .IN2(n12781), .IN1(n12779), .Q(n12794) );
  OR2X1 U16063 ( .IN2(n12784), .IN1(n12783), .Q(n12788) );
  OR2X1 U16064 ( .IN2(n12786), .IN1(n12785), .Q(n12790) );
  OR2X1 U16065 ( .IN2(n12789), .IN1(n12787), .Q(n12793) );
  OR2X1 U16066 ( .IN2(n12792), .IN1(n12791), .Q(n12795) );
  OR2X1 U16067 ( .IN2(n12797), .IN1(n12796), .Q(n12801) );
  OR2X1 U16068 ( .IN2(n12799), .IN1(n12798), .Q(n12803) );
  OR2X1 U16069 ( .IN2(n12802), .IN1(n12800), .Q(n12813) );
  OR2X1 U16070 ( .IN2(n12805), .IN1(n12804), .Q(n12809) );
  OR2X1 U16071 ( .IN2(n12807), .IN1(n12806), .Q(n12811) );
  OR2X1 U16072 ( .IN2(n12810), .IN1(n12808), .Q(n12815) );
  OR2X1 U16073 ( .IN2(n12814), .IN1(n12812), .Q(n12827) );
  OR2X1 U16074 ( .IN2(n12817), .IN1(n12816), .Q(n12821) );
  OR2X1 U16075 ( .IN2(n12819), .IN1(n12818), .Q(n12823) );
  OR2X1 U16076 ( .IN2(n12822), .IN1(n12820), .Q(n12826) );
  OR2X1 U16077 ( .IN2(n12825), .IN1(n12824), .Q(n12828) );
  OR2X1 U16078 ( .IN2(n12830), .IN1(n12829), .Q(n12834) );
  OR2X1 U16079 ( .IN2(n12832), .IN1(n12831), .Q(n12836) );
  OR2X1 U16080 ( .IN2(n12835), .IN1(n12833), .Q(n12846) );
  OR2X1 U16081 ( .IN2(n12838), .IN1(n12837), .Q(n12842) );
  OR2X1 U16082 ( .IN2(n12840), .IN1(n12839), .Q(n12844) );
  OR2X1 U16083 ( .IN2(n12843), .IN1(n12841), .Q(n12848) );
  OR2X1 U16084 ( .IN2(n12847), .IN1(n12845), .Q(n12860) );
  OR2X1 U16085 ( .IN2(n12850), .IN1(n12849), .Q(n12854) );
  OR2X1 U16086 ( .IN2(n12852), .IN1(n12851), .Q(n12856) );
  OR2X1 U16087 ( .IN2(n12855), .IN1(n12853), .Q(n12859) );
  OR2X1 U16088 ( .IN2(n12858), .IN1(n12857), .Q(n12861) );
  OR2X1 U16089 ( .IN2(n12863), .IN1(n12862), .Q(n12867) );
  OR2X1 U16090 ( .IN2(n12865), .IN1(n12864), .Q(n12869) );
  OR2X1 U16091 ( .IN2(n12868), .IN1(n12866), .Q(n12879) );
  OR2X1 U16092 ( .IN2(n12871), .IN1(n12870), .Q(n12875) );
  OR2X1 U16093 ( .IN2(n12873), .IN1(n12872), .Q(n12877) );
  OR2X1 U16094 ( .IN2(n12876), .IN1(n12874), .Q(n12881) );
  OR2X1 U16095 ( .IN2(n12880), .IN1(n12878), .Q(n12893) );
  OR2X1 U16096 ( .IN2(n12883), .IN1(n12882), .Q(n12887) );
  OR2X1 U16097 ( .IN2(n12885), .IN1(n12884), .Q(n12889) );
  OR2X1 U16098 ( .IN2(n12888), .IN1(n12886), .Q(n12892) );
  OR2X1 U16099 ( .IN2(n12891), .IN1(n12890), .Q(n12894) );
  OR2X1 U16100 ( .IN2(n12896), .IN1(n12895), .Q(n12900) );
  OR2X1 U16101 ( .IN2(n12898), .IN1(n12897), .Q(n12902) );
  OR2X1 U16102 ( .IN2(n12901), .IN1(n12899), .Q(n12912) );
  OR2X1 U16103 ( .IN2(n12904), .IN1(n12903), .Q(n12908) );
  OR2X1 U16104 ( .IN2(n12906), .IN1(n12905), .Q(n12910) );
  OR2X1 U16105 ( .IN2(n12909), .IN1(n12907), .Q(n12914) );
  OR2X1 U16106 ( .IN2(n12913), .IN1(n12911), .Q(n12926) );
  OR2X1 U16107 ( .IN2(n12916), .IN1(n12915), .Q(n12920) );
  OR2X1 U16108 ( .IN2(n12918), .IN1(n12917), .Q(n12922) );
  OR2X1 U16109 ( .IN2(n12921), .IN1(n12919), .Q(n12925) );
  OR2X1 U16110 ( .IN2(n12924), .IN1(n12923), .Q(n12927) );
  OR2X1 U16111 ( .IN2(n12929), .IN1(n12928), .Q(n12933) );
  OR2X1 U16112 ( .IN2(n12931), .IN1(n12930), .Q(n12935) );
  OR2X1 U16113 ( .IN2(n12934), .IN1(n12932), .Q(n12945) );
  OR2X1 U16114 ( .IN2(n12937), .IN1(n12936), .Q(n12941) );
  OR2X1 U16115 ( .IN2(n12939), .IN1(n12938), .Q(n12943) );
  OR2X1 U16116 ( .IN2(n12942), .IN1(n12940), .Q(n12947) );
  OR2X1 U16117 ( .IN2(n12946), .IN1(n12944), .Q(n12959) );
  OR2X1 U16118 ( .IN2(n12949), .IN1(n12948), .Q(n12953) );
  OR2X1 U15933 ( .IN2(n12393), .IN1(n12391), .Q(n12398) );
  OR2X1 U15934 ( .IN2(n12397), .IN1(n12395), .Q(n12413) );
  OR2X1 U15935 ( .IN2(n12400), .IN1(n12399), .Q(n12404) );
  OR2X1 U15936 ( .IN2(n12402), .IN1(n12401), .Q(n12406) );
  OR2X1 U15937 ( .IN2(n12405), .IN1(n12403), .Q(n12410) );
  OR2X1 U15938 ( .IN2(n12408), .IN1(n12407), .Q(n12412) );
  OR2X1 U15939 ( .IN2(n12411), .IN1(n12409), .Q(n12414) );
  OR2X1 U15940 ( .IN2(n12416), .IN1(n12415), .Q(n12420) );
  OR2X1 U15941 ( .IN2(n12418), .IN1(n12417), .Q(n12422) );
  OR2X1 U15942 ( .IN2(n12421), .IN1(n12419), .Q(n12432) );
  OR2X1 U15943 ( .IN2(n12424), .IN1(n12423), .Q(n12428) );
  OR2X1 U15944 ( .IN2(n12426), .IN1(n12425), .Q(n12430) );
  OR2X1 U15945 ( .IN2(n12429), .IN1(n12427), .Q(n12434) );
  OR2X1 U15946 ( .IN2(n12433), .IN1(n12431), .Q(n12449) );
  OR2X1 U15947 ( .IN2(n12436), .IN1(n12435), .Q(n12440) );
  OR2X1 U15948 ( .IN2(n12438), .IN1(n12437), .Q(n12442) );
  OR2X1 U15949 ( .IN2(n12441), .IN1(n12439), .Q(n12446) );
  OR2X1 U15950 ( .IN2(n12444), .IN1(n12443), .Q(n12448) );
  OR2X1 U15951 ( .IN2(n12447), .IN1(n12445), .Q(n12450) );
  OR2X1 U15952 ( .IN2(n12452), .IN1(n12451), .Q(n12456) );
  OR2X1 U15953 ( .IN2(n12454), .IN1(n12453), .Q(n12458) );
  OR2X1 U15954 ( .IN2(n12457), .IN1(n12455), .Q(n12468) );
  OR2X1 U15955 ( .IN2(n12460), .IN1(n12459), .Q(n12464) );
  OR2X1 U15956 ( .IN2(n12462), .IN1(n12461), .Q(n12466) );
  OR2X1 U15957 ( .IN2(n12465), .IN1(n12463), .Q(n12470) );
  OR2X1 U15958 ( .IN2(n12469), .IN1(n12467), .Q(n12485) );
  OR2X1 U15959 ( .IN2(n12472), .IN1(n12471), .Q(n12476) );
  OR2X1 U15960 ( .IN2(n12474), .IN1(n12473), .Q(n12478) );
  OR2X1 U15961 ( .IN2(n12477), .IN1(n12475), .Q(n12482) );
  OR2X1 U15962 ( .IN2(n12480), .IN1(n12479), .Q(n12484) );
  OR2X1 U15963 ( .IN2(n12483), .IN1(n12481), .Q(n12486) );
  OR2X1 U15964 ( .IN2(n12488), .IN1(n12487), .Q(n12492) );
  OR2X1 U15965 ( .IN2(n12490), .IN1(n12489), .Q(n12494) );
  OR2X1 U15966 ( .IN2(n12493), .IN1(n12491), .Q(n12504) );
  OR2X1 U15967 ( .IN2(n12496), .IN1(n12495), .Q(n12500) );
  OR2X1 U15968 ( .IN2(n12498), .IN1(n12497), .Q(n12502) );
  OR2X1 U15969 ( .IN2(n12501), .IN1(n12499), .Q(n12506) );
  OR2X1 U15970 ( .IN2(n12505), .IN1(n12503), .Q(n12521) );
  OR2X1 U15971 ( .IN2(n12508), .IN1(n12507), .Q(n12512) );
  OR2X1 U15972 ( .IN2(n12510), .IN1(n12509), .Q(n12514) );
  OR2X1 U15973 ( .IN2(n12513), .IN1(n12511), .Q(n12518) );
  OR2X1 U15974 ( .IN2(n12516), .IN1(n12515), .Q(n12520) );
  OR2X1 U15975 ( .IN2(n12519), .IN1(n12517), .Q(n12522) );
  OR2X1 U15976 ( .IN2(n12524), .IN1(n12523), .Q(n12528) );
  OR2X1 U15977 ( .IN2(n12526), .IN1(n12525), .Q(n12530) );
  OR2X1 U15978 ( .IN2(n12529), .IN1(n12527), .Q(n12540) );
  OR2X1 U15979 ( .IN2(n12532), .IN1(n12531), .Q(n12536) );
  OR2X1 U15980 ( .IN2(n12534), .IN1(n12533), .Q(n12538) );
  OR2X1 U15981 ( .IN2(n12537), .IN1(n12535), .Q(n12542) );
  OR2X1 U15982 ( .IN2(n12541), .IN1(n12539), .Q(n12557) );
  OR2X1 U15983 ( .IN2(n12544), .IN1(n12543), .Q(n12548) );
  OR2X1 U15984 ( .IN2(n12546), .IN1(n12545), .Q(n12550) );
  OR2X1 U15985 ( .IN2(n12549), .IN1(n12547), .Q(n12554) );
  OR2X1 U15986 ( .IN2(n12552), .IN1(n12551), .Q(n12556) );
  OR2X1 U15987 ( .IN2(n12555), .IN1(n12553), .Q(n12558) );
  OR2X1 U15988 ( .IN2(n12560), .IN1(n12559), .Q(n12564) );
  OR2X1 U15989 ( .IN2(n12562), .IN1(n12561), .Q(n12566) );
  OR2X1 U15990 ( .IN2(n12565), .IN1(n12563), .Q(n12576) );
  OR2X1 U15991 ( .IN2(n12568), .IN1(n12567), .Q(n12572) );
  OR2X1 U15992 ( .IN2(n12570), .IN1(n12569), .Q(n12574) );
  OR2X1 U15993 ( .IN2(n12573), .IN1(n12571), .Q(n12578) );
  OR2X1 U15994 ( .IN2(n12577), .IN1(n12575), .Q(n12593) );
  OR2X1 U15995 ( .IN2(n12580), .IN1(n12579), .Q(n12584) );
  OR2X1 U15996 ( .IN2(n12582), .IN1(n12581), .Q(n12586) );
  OR2X1 U15997 ( .IN2(n12585), .IN1(n12583), .Q(n12590) );
  OR2X1 U15998 ( .IN2(n12588), .IN1(n12587), .Q(n12592) );
  OR2X1 U15999 ( .IN2(n12591), .IN1(n12589), .Q(n12594) );
  OR2X1 U16000 ( .IN2(n12596), .IN1(n12595), .Q(n12600) );
  OR2X1 U16001 ( .IN2(n12598), .IN1(n12597), .Q(n12602) );
  OR2X1 U16002 ( .IN2(n12601), .IN1(n12599), .Q(n12612) );
  OR2X1 U16003 ( .IN2(n12604), .IN1(n12603), .Q(n12608) );
  OR2X1 U16004 ( .IN2(n12606), .IN1(n12605), .Q(n12610) );
  OR2X1 U16005 ( .IN2(n12609), .IN1(n12607), .Q(n12614) );
  OR2X1 U16006 ( .IN2(n12613), .IN1(n12611), .Q(n12629) );
  OR2X1 U16007 ( .IN2(n12616), .IN1(n12615), .Q(n12620) );
  OR2X1 U16008 ( .IN2(n12618), .IN1(n12617), .Q(n12622) );
  OR2X1 U16009 ( .IN2(n12621), .IN1(n12619), .Q(n12626) );
  OR2X1 U16010 ( .IN2(n12624), .IN1(n12623), .Q(n12628) );
  OR2X1 U16011 ( .IN2(n12627), .IN1(n12625), .Q(n12630) );
  OR2X1 U16012 ( .IN2(n12632), .IN1(n12631), .Q(n12636) );
  OR2X1 U16013 ( .IN2(n12634), .IN1(n12633), .Q(n12638) );
  OR2X1 U16014 ( .IN2(n12637), .IN1(n12635), .Q(n12648) );
  OR2X1 U16015 ( .IN2(n12640), .IN1(n12639), .Q(n12644) );
  OR2X1 U16016 ( .IN2(n12642), .IN1(n12641), .Q(n12646) );
  OR2X1 U16017 ( .IN2(n12645), .IN1(n12643), .Q(n12650) );
  OR2X1 U16018 ( .IN2(n12649), .IN1(n12647), .Q(n12662) );
  OR2X1 U16019 ( .IN2(n12652), .IN1(n12651), .Q(n12656) );
  OR2X1 U16020 ( .IN2(n12654), .IN1(n12653), .Q(n12658) );
  OR2X1 U16021 ( .IN2(n12657), .IN1(n12655), .Q(n12661) );
  OR2X1 U16022 ( .IN2(n12660), .IN1(n12659), .Q(n12663) );
  OR2X1 U16023 ( .IN2(n12665), .IN1(n12664), .Q(n12669) );
  OR2X1 U16024 ( .IN2(n12667), .IN1(n12666), .Q(n12671) );
  OR2X1 U16025 ( .IN2(n12670), .IN1(n12668), .Q(n12681) );
  OR2X1 U15840 ( .IN2(n12114), .IN1(n12113), .Q(n12118) );
  OR2X1 U15841 ( .IN2(n12117), .IN1(n12115), .Q(n12122) );
  OR2X1 U15842 ( .IN2(n12120), .IN1(n12119), .Q(n12124) );
  OR2X1 U15843 ( .IN2(n12123), .IN1(n12121), .Q(n12126) );
  OR2X1 U15844 ( .IN2(n12128), .IN1(n12127), .Q(n12132) );
  OR2X1 U15845 ( .IN2(n12130), .IN1(n12129), .Q(n12134) );
  OR2X1 U15846 ( .IN2(n12133), .IN1(n12131), .Q(n12144) );
  OR2X1 U15847 ( .IN2(n12136), .IN1(n12135), .Q(n12140) );
  OR2X1 U15848 ( .IN2(n12138), .IN1(n12137), .Q(n12142) );
  OR2X1 U15849 ( .IN2(n12141), .IN1(n12139), .Q(n12146) );
  OR2X1 U15850 ( .IN2(n12145), .IN1(n12143), .Q(n12161) );
  OR2X1 U15851 ( .IN2(n12148), .IN1(n12147), .Q(n12152) );
  OR2X1 U15852 ( .IN2(n12150), .IN1(n12149), .Q(n12154) );
  OR2X1 U15853 ( .IN2(n12153), .IN1(n12151), .Q(n12158) );
  OR2X1 U15854 ( .IN2(n12156), .IN1(n12155), .Q(n12160) );
  OR2X1 U15855 ( .IN2(n12159), .IN1(n12157), .Q(n12162) );
  OR2X1 U15856 ( .IN2(n12164), .IN1(n12163), .Q(n12168) );
  OR2X1 U15857 ( .IN2(n12166), .IN1(n12165), .Q(n12170) );
  OR2X1 U15858 ( .IN2(n12169), .IN1(n12167), .Q(n12180) );
  OR2X1 U15859 ( .IN2(n12172), .IN1(n12171), .Q(n12176) );
  OR2X1 U15860 ( .IN2(n12174), .IN1(n12173), .Q(n12178) );
  OR2X1 U15861 ( .IN2(n12177), .IN1(n12175), .Q(n12182) );
  OR2X1 U15862 ( .IN2(n12181), .IN1(n12179), .Q(n12197) );
  OR2X1 U15863 ( .IN2(n12184), .IN1(n12183), .Q(n12188) );
  OR2X1 U15864 ( .IN2(n12186), .IN1(n12185), .Q(n12190) );
  OR2X1 U15865 ( .IN2(n12189), .IN1(n12187), .Q(n12194) );
  OR2X1 U15866 ( .IN2(n12192), .IN1(n12191), .Q(n12196) );
  OR2X1 U15867 ( .IN2(n12195), .IN1(n12193), .Q(n12198) );
  OR2X1 U15868 ( .IN2(n12200), .IN1(n12199), .Q(n12204) );
  OR2X1 U15869 ( .IN2(n12202), .IN1(n12201), .Q(n12206) );
  OR2X1 U15870 ( .IN2(n12205), .IN1(n12203), .Q(n12216) );
  OR2X1 U15871 ( .IN2(n12208), .IN1(n12207), .Q(n12212) );
  OR2X1 U15872 ( .IN2(n12210), .IN1(n12209), .Q(n12214) );
  OR2X1 U15873 ( .IN2(n12213), .IN1(n12211), .Q(n12218) );
  OR2X1 U15874 ( .IN2(n12217), .IN1(n12215), .Q(n12233) );
  OR2X1 U15875 ( .IN2(n12220), .IN1(n12219), .Q(n12224) );
  OR2X1 U15876 ( .IN2(n12222), .IN1(n12221), .Q(n12226) );
  OR2X1 U15877 ( .IN2(n12225), .IN1(n12223), .Q(n12230) );
  OR2X1 U15878 ( .IN2(n12228), .IN1(n12227), .Q(n12232) );
  OR2X1 U15879 ( .IN2(n12231), .IN1(n12229), .Q(n12234) );
  OR2X1 U15880 ( .IN2(n12236), .IN1(n12235), .Q(n12240) );
  OR2X1 U15881 ( .IN2(n12238), .IN1(n12237), .Q(n12242) );
  OR2X1 U15882 ( .IN2(n12241), .IN1(n12239), .Q(n12252) );
  OR2X1 U15883 ( .IN2(n12244), .IN1(n12243), .Q(n12248) );
  OR2X1 U15884 ( .IN2(n12246), .IN1(n12245), .Q(n12250) );
  OR2X1 U15885 ( .IN2(n12249), .IN1(n12247), .Q(n12254) );
  OR2X1 U15886 ( .IN2(n12253), .IN1(n12251), .Q(n12269) );
  OR2X1 U15887 ( .IN2(n12256), .IN1(n12255), .Q(n12260) );
  OR2X1 U15888 ( .IN2(n12258), .IN1(n12257), .Q(n12262) );
  OR2X1 U15889 ( .IN2(n12261), .IN1(n12259), .Q(n12266) );
  OR2X1 U15890 ( .IN2(n12264), .IN1(n12263), .Q(n12268) );
  OR2X1 U15891 ( .IN2(n12267), .IN1(n12265), .Q(n12270) );
  OR2X1 U15892 ( .IN2(n12272), .IN1(n12271), .Q(n12276) );
  OR2X1 U15893 ( .IN2(n12274), .IN1(n12273), .Q(n12278) );
  OR2X1 U15894 ( .IN2(n12277), .IN1(n12275), .Q(n12288) );
  OR2X1 U15895 ( .IN2(n12280), .IN1(n12279), .Q(n12284) );
  OR2X1 U15896 ( .IN2(n12282), .IN1(n12281), .Q(n12286) );
  OR2X1 U15897 ( .IN2(n12285), .IN1(n12283), .Q(n12290) );
  OR2X1 U15898 ( .IN2(n12289), .IN1(n12287), .Q(n12305) );
  OR2X1 U15899 ( .IN2(n12292), .IN1(n12291), .Q(n12296) );
  OR2X1 U15900 ( .IN2(n12294), .IN1(n12293), .Q(n12298) );
  OR2X1 U15901 ( .IN2(n12297), .IN1(n12295), .Q(n12302) );
  OR2X1 U15902 ( .IN2(n12300), .IN1(n12299), .Q(n12304) );
  OR2X1 U15903 ( .IN2(n12303), .IN1(n12301), .Q(n12306) );
  OR2X1 U15904 ( .IN2(n12308), .IN1(n12307), .Q(n12312) );
  OR2X1 U15905 ( .IN2(n12310), .IN1(n12309), .Q(n12314) );
  OR2X1 U15906 ( .IN2(n12313), .IN1(n12311), .Q(n12324) );
  OR2X1 U15907 ( .IN2(n12316), .IN1(n12315), .Q(n12320) );
  OR2X1 U15908 ( .IN2(n12318), .IN1(n12317), .Q(n12322) );
  OR2X1 U15909 ( .IN2(n12321), .IN1(n12319), .Q(n12326) );
  OR2X1 U15910 ( .IN2(n12325), .IN1(n12323), .Q(n12341) );
  OR2X1 U15911 ( .IN2(n12328), .IN1(n12327), .Q(n12332) );
  OR2X1 U15912 ( .IN2(n12330), .IN1(n12329), .Q(n12334) );
  OR2X1 U15913 ( .IN2(n12333), .IN1(n12331), .Q(n12338) );
  OR2X1 U15914 ( .IN2(n12336), .IN1(n12335), .Q(n12340) );
  OR2X1 U15915 ( .IN2(n12339), .IN1(n12337), .Q(n12342) );
  OR2X1 U15916 ( .IN2(n12344), .IN1(n12343), .Q(n12348) );
  OR2X1 U15917 ( .IN2(n12346), .IN1(n12345), .Q(n12350) );
  OR2X1 U15918 ( .IN2(n12349), .IN1(n12347), .Q(n12360) );
  OR2X1 U15919 ( .IN2(n12352), .IN1(n12351), .Q(n12356) );
  OR2X1 U15920 ( .IN2(n12354), .IN1(n12353), .Q(n12358) );
  OR2X1 U15921 ( .IN2(n12357), .IN1(n12355), .Q(n12362) );
  OR2X1 U15922 ( .IN2(n12361), .IN1(n12359), .Q(n12377) );
  OR2X1 U15923 ( .IN2(n12364), .IN1(n12363), .Q(n12368) );
  OR2X1 U15924 ( .IN2(n12366), .IN1(n12365), .Q(n12370) );
  OR2X1 U15925 ( .IN2(n12369), .IN1(n12367), .Q(n12374) );
  OR2X1 U15926 ( .IN2(n12372), .IN1(n12371), .Q(n12376) );
  OR2X1 U15927 ( .IN2(n12375), .IN1(n12373), .Q(n12378) );
  OR2X1 U15928 ( .IN2(n12380), .IN1(n12379), .Q(n12384) );
  OR2X1 U15929 ( .IN2(n12382), .IN1(n12381), .Q(n12386) );
  OR2X1 U15930 ( .IN2(n12385), .IN1(n12383), .Q(n12396) );
  OR2X1 U15931 ( .IN2(n12388), .IN1(n12387), .Q(n12392) );
  OR2X1 U15932 ( .IN2(n12390), .IN1(n12389), .Q(n12394) );
  OR2X1 U15747 ( .IN2(n11835), .IN1(n11833), .Q(n11838) );
  OR2X1 U15748 ( .IN2(n11840), .IN1(n11839), .Q(n11844) );
  OR2X1 U15749 ( .IN2(n11842), .IN1(n11841), .Q(n11846) );
  OR2X1 U15750 ( .IN2(n11845), .IN1(n11843), .Q(n11856) );
  OR2X1 U15751 ( .IN2(n11848), .IN1(n11847), .Q(n11852) );
  OR2X1 U15752 ( .IN2(n11850), .IN1(n11849), .Q(n11854) );
  OR2X1 U15753 ( .IN2(n11853), .IN1(n11851), .Q(n11858) );
  OR2X1 U15754 ( .IN2(n11857), .IN1(n11855), .Q(n11873) );
  OR2X1 U15755 ( .IN2(n11860), .IN1(n11859), .Q(n11864) );
  OR2X1 U15756 ( .IN2(n11862), .IN1(n11861), .Q(n11866) );
  OR2X1 U15757 ( .IN2(n11865), .IN1(n11863), .Q(n11870) );
  OR2X1 U15758 ( .IN2(n11868), .IN1(n11867), .Q(n11872) );
  OR2X1 U15759 ( .IN2(n11871), .IN1(n11869), .Q(n11874) );
  OR2X1 U15760 ( .IN2(n11876), .IN1(n11875), .Q(n11880) );
  OR2X1 U15761 ( .IN2(n11878), .IN1(n11877), .Q(n11882) );
  OR2X1 U15762 ( .IN2(n11881), .IN1(n11879), .Q(n11892) );
  OR2X1 U15763 ( .IN2(n11884), .IN1(n11883), .Q(n11888) );
  OR2X1 U15764 ( .IN2(n11886), .IN1(n11885), .Q(n11890) );
  OR2X1 U15765 ( .IN2(n11889), .IN1(n11887), .Q(n11894) );
  OR2X1 U15766 ( .IN2(n11893), .IN1(n11891), .Q(n11909) );
  OR2X1 U15767 ( .IN2(n11896), .IN1(n11895), .Q(n11900) );
  OR2X1 U15768 ( .IN2(n11898), .IN1(n11897), .Q(n11902) );
  OR2X1 U15769 ( .IN2(n11901), .IN1(n11899), .Q(n11906) );
  OR2X1 U15770 ( .IN2(n11904), .IN1(n11903), .Q(n11908) );
  OR2X1 U15771 ( .IN2(n11907), .IN1(n11905), .Q(n11910) );
  OR2X1 U15772 ( .IN2(n11912), .IN1(n11911), .Q(n11916) );
  OR2X1 U15773 ( .IN2(n11914), .IN1(n11913), .Q(n11918) );
  OR2X1 U15774 ( .IN2(n11917), .IN1(n11915), .Q(n11928) );
  OR2X1 U15775 ( .IN2(n11920), .IN1(n11919), .Q(n11924) );
  OR2X1 U15776 ( .IN2(n11922), .IN1(n11921), .Q(n11926) );
  OR2X1 U15777 ( .IN2(n11925), .IN1(n11923), .Q(n11930) );
  OR2X1 U15778 ( .IN2(n11929), .IN1(n11927), .Q(n11945) );
  OR2X1 U15779 ( .IN2(n11932), .IN1(n11931), .Q(n11936) );
  OR2X1 U15780 ( .IN2(n11934), .IN1(n11933), .Q(n11938) );
  OR2X1 U15781 ( .IN2(n11937), .IN1(n11935), .Q(n11942) );
  OR2X1 U15782 ( .IN2(n11940), .IN1(n11939), .Q(n11944) );
  OR2X1 U15783 ( .IN2(n11943), .IN1(n11941), .Q(n11946) );
  OR2X1 U15784 ( .IN2(n11948), .IN1(n11947), .Q(n11952) );
  OR2X1 U15785 ( .IN2(n11950), .IN1(n11949), .Q(n11954) );
  OR2X1 U15786 ( .IN2(n11953), .IN1(n11951), .Q(n11964) );
  OR2X1 U15787 ( .IN2(n11956), .IN1(n11955), .Q(n11960) );
  OR2X1 U15788 ( .IN2(n11958), .IN1(n11957), .Q(n11962) );
  OR2X1 U15789 ( .IN2(n11961), .IN1(n11959), .Q(n11966) );
  OR2X1 U15790 ( .IN2(n11965), .IN1(n11963), .Q(n11981) );
  OR2X1 U15791 ( .IN2(n11968), .IN1(n11967), .Q(n11972) );
  OR2X1 U15792 ( .IN2(n11970), .IN1(n11969), .Q(n11974) );
  OR2X1 U15793 ( .IN2(n11973), .IN1(n11971), .Q(n11978) );
  OR2X1 U15794 ( .IN2(n11976), .IN1(n11975), .Q(n11980) );
  OR2X1 U15795 ( .IN2(n11979), .IN1(n11977), .Q(n11982) );
  OR2X1 U15796 ( .IN2(n11984), .IN1(n11983), .Q(n11988) );
  OR2X1 U15797 ( .IN2(n11986), .IN1(n11985), .Q(n11990) );
  OR2X1 U15798 ( .IN2(n11989), .IN1(n11987), .Q(n12000) );
  OR2X1 U15799 ( .IN2(n11992), .IN1(n11991), .Q(n11996) );
  OR2X1 U15800 ( .IN2(n11994), .IN1(n11993), .Q(n11998) );
  OR2X1 U15801 ( .IN2(n11997), .IN1(n11995), .Q(n12002) );
  OR2X1 U15802 ( .IN2(n12001), .IN1(n11999), .Q(n12017) );
  OR2X1 U15803 ( .IN2(n12004), .IN1(n12003), .Q(n12008) );
  OR2X1 U15804 ( .IN2(n12006), .IN1(n12005), .Q(n12010) );
  OR2X1 U15805 ( .IN2(n12009), .IN1(n12007), .Q(n12014) );
  OR2X1 U15806 ( .IN2(n12012), .IN1(n12011), .Q(n12016) );
  OR2X1 U15807 ( .IN2(n12015), .IN1(n12013), .Q(n12018) );
  OR2X1 U15808 ( .IN2(n12020), .IN1(n12019), .Q(n12024) );
  OR2X1 U15809 ( .IN2(n12022), .IN1(n12021), .Q(n12026) );
  OR2X1 U15810 ( .IN2(n12025), .IN1(n12023), .Q(n12036) );
  OR2X1 U15811 ( .IN2(n12028), .IN1(n12027), .Q(n12032) );
  OR2X1 U15812 ( .IN2(n12030), .IN1(n12029), .Q(n12034) );
  OR2X1 U15813 ( .IN2(n12033), .IN1(n12031), .Q(n12038) );
  OR2X1 U15814 ( .IN2(n12037), .IN1(n12035), .Q(n12053) );
  OR2X1 U15815 ( .IN2(n12040), .IN1(n12039), .Q(n12044) );
  OR2X1 U15816 ( .IN2(n12042), .IN1(n12041), .Q(n12046) );
  OR2X1 U15817 ( .IN2(n12045), .IN1(n12043), .Q(n12050) );
  OR2X1 U15818 ( .IN2(n12048), .IN1(n12047), .Q(n12052) );
  OR2X1 U15819 ( .IN2(n12051), .IN1(n12049), .Q(n12054) );
  OR2X1 U15820 ( .IN2(n12056), .IN1(n12055), .Q(n12060) );
  OR2X1 U15821 ( .IN2(n12058), .IN1(n12057), .Q(n12062) );
  OR2X1 U15822 ( .IN2(n12061), .IN1(n12059), .Q(n12072) );
  OR2X1 U15823 ( .IN2(n12064), .IN1(n12063), .Q(n12068) );
  OR2X1 U15824 ( .IN2(n12066), .IN1(n12065), .Q(n12070) );
  OR2X1 U15825 ( .IN2(n12069), .IN1(n12067), .Q(n12074) );
  OR2X1 U15826 ( .IN2(n12073), .IN1(n12071), .Q(n12089) );
  OR2X1 U15827 ( .IN2(n12076), .IN1(n12075), .Q(n12080) );
  OR2X1 U15828 ( .IN2(n12078), .IN1(n12077), .Q(n12082) );
  OR2X1 U15829 ( .IN2(n12081), .IN1(n12079), .Q(n12086) );
  OR2X1 U15830 ( .IN2(n12084), .IN1(n12083), .Q(n12088) );
  OR2X1 U15831 ( .IN2(n12087), .IN1(n12085), .Q(n12090) );
  OR2X1 U15832 ( .IN2(n12092), .IN1(n12091), .Q(n12096) );
  OR2X1 U15833 ( .IN2(n12094), .IN1(n12093), .Q(n12098) );
  OR2X1 U15834 ( .IN2(n12097), .IN1(n12095), .Q(n12108) );
  OR2X1 U15835 ( .IN2(n12100), .IN1(n12099), .Q(n12104) );
  OR2X1 U15836 ( .IN2(n12102), .IN1(n12101), .Q(n12106) );
  OR2X1 U15837 ( .IN2(n12105), .IN1(n12103), .Q(n12110) );
  OR2X1 U15838 ( .IN2(n12109), .IN1(n12107), .Q(n12125) );
  OR2X1 U15839 ( .IN2(n12112), .IN1(n12111), .Q(n12116) );
  OR2X1 U15654 ( .IN2(n11555), .IN1(n11554), .Q(n11559) );
  OR2X1 U15655 ( .IN2(n11558), .IN1(n11556), .Q(n11563) );
  OR2X1 U15656 ( .IN2(n11562), .IN1(n11560), .Q(n11585) );
  OR2X1 U15657 ( .IN2(n11565), .IN1(n11564), .Q(n11569) );
  OR2X1 U15658 ( .IN2(n11567), .IN1(n11566), .Q(n11571) );
  OR2X1 U15659 ( .IN2(n11570), .IN1(n11568), .Q(n11581) );
  OR2X1 U15660 ( .IN2(n11573), .IN1(n11572), .Q(n11577) );
  OR2X1 U15661 ( .IN2(n11575), .IN1(n11574), .Q(n11579) );
  OR2X1 U15662 ( .IN2(n11578), .IN1(n11576), .Q(n11583) );
  OR2X1 U15663 ( .IN2(n11582), .IN1(n11580), .Q(n11586) );
  OR2X1 U15664 ( .IN2(n11588), .IN1(n11587), .Q(n11592) );
  OR2X1 U15665 ( .IN2(n11590), .IN1(n11589), .Q(n11594) );
  OR2X1 U15666 ( .IN2(n11593), .IN1(n11591), .Q(n11604) );
  OR2X1 U15667 ( .IN2(n11596), .IN1(n11595), .Q(n11600) );
  OR2X1 U15668 ( .IN2(n11598), .IN1(n11597), .Q(n11602) );
  OR2X1 U15669 ( .IN2(n11601), .IN1(n11599), .Q(n11606) );
  OR2X1 U15670 ( .IN2(n11605), .IN1(n11603), .Q(n11621) );
  OR2X1 U15671 ( .IN2(n11608), .IN1(n11607), .Q(n11612) );
  OR2X1 U15672 ( .IN2(n11610), .IN1(n11609), .Q(n11614) );
  OR2X1 U15673 ( .IN2(n11613), .IN1(n11611), .Q(n11618) );
  OR2X1 U15674 ( .IN2(n11616), .IN1(n11615), .Q(n11620) );
  OR2X1 U15675 ( .IN2(n11619), .IN1(n11617), .Q(n11622) );
  OR2X1 U15676 ( .IN2(n11624), .IN1(n11623), .Q(n11628) );
  OR2X1 U15677 ( .IN2(n11626), .IN1(n11625), .Q(n11630) );
  OR2X1 U15678 ( .IN2(n11629), .IN1(n11627), .Q(n11640) );
  OR2X1 U15679 ( .IN2(n11632), .IN1(n11631), .Q(n11636) );
  OR2X1 U15680 ( .IN2(n11634), .IN1(n11633), .Q(n11638) );
  OR2X1 U15681 ( .IN2(n11637), .IN1(n11635), .Q(n11642) );
  OR2X1 U15682 ( .IN2(n11641), .IN1(n11639), .Q(n11657) );
  OR2X1 U15683 ( .IN2(n11644), .IN1(n11643), .Q(n11648) );
  OR2X1 U15684 ( .IN2(n11646), .IN1(n11645), .Q(n11650) );
  OR2X1 U15685 ( .IN2(n11649), .IN1(n11647), .Q(n11654) );
  OR2X1 U15686 ( .IN2(n11652), .IN1(n11651), .Q(n11656) );
  OR2X1 U15687 ( .IN2(n11655), .IN1(n11653), .Q(n11658) );
  OR2X1 U15688 ( .IN2(n11660), .IN1(n11659), .Q(n11664) );
  OR2X1 U15689 ( .IN2(n11662), .IN1(n11661), .Q(n11666) );
  OR2X1 U15690 ( .IN2(n11665), .IN1(n11663), .Q(n11676) );
  OR2X1 U15691 ( .IN2(n11668), .IN1(n11667), .Q(n11672) );
  OR2X1 U15692 ( .IN2(n11670), .IN1(n11669), .Q(n11674) );
  OR2X1 U15693 ( .IN2(n11673), .IN1(n11671), .Q(n11678) );
  OR2X1 U15694 ( .IN2(n11677), .IN1(n11675), .Q(n11693) );
  OR2X1 U15695 ( .IN2(n11680), .IN1(n11679), .Q(n11684) );
  OR2X1 U15696 ( .IN2(n11682), .IN1(n11681), .Q(n11686) );
  OR2X1 U15697 ( .IN2(n11685), .IN1(n11683), .Q(n11690) );
  OR2X1 U15698 ( .IN2(n11688), .IN1(n11687), .Q(n11692) );
  OR2X1 U15699 ( .IN2(n11691), .IN1(n11689), .Q(n11694) );
  OR2X1 U15700 ( .IN2(n11696), .IN1(n11695), .Q(n11700) );
  OR2X1 U15701 ( .IN2(n11698), .IN1(n11697), .Q(n11702) );
  OR2X1 U15702 ( .IN2(n11701), .IN1(n11699), .Q(n11712) );
  OR2X1 U15703 ( .IN2(n11704), .IN1(n11703), .Q(n11708) );
  OR2X1 U15704 ( .IN2(n11706), .IN1(n11705), .Q(n11710) );
  OR2X1 U15705 ( .IN2(n11709), .IN1(n11707), .Q(n11714) );
  OR2X1 U15706 ( .IN2(n11713), .IN1(n11711), .Q(n11729) );
  OR2X1 U15707 ( .IN2(n11716), .IN1(n11715), .Q(n11720) );
  OR2X1 U15708 ( .IN2(n11718), .IN1(n11717), .Q(n11722) );
  OR2X1 U15709 ( .IN2(n11721), .IN1(n11719), .Q(n11726) );
  OR2X1 U15710 ( .IN2(n11724), .IN1(n11723), .Q(n11728) );
  OR2X1 U15711 ( .IN2(n11727), .IN1(n11725), .Q(n11730) );
  OR2X1 U15712 ( .IN2(n11732), .IN1(n11731), .Q(n11736) );
  OR2X1 U15713 ( .IN2(n11734), .IN1(n11733), .Q(n11738) );
  OR2X1 U15714 ( .IN2(n11737), .IN1(n11735), .Q(n11748) );
  OR2X1 U15715 ( .IN2(n11740), .IN1(n11739), .Q(n11744) );
  OR2X1 U15716 ( .IN2(n11742), .IN1(n11741), .Q(n11746) );
  OR2X1 U15717 ( .IN2(n11745), .IN1(n11743), .Q(n11750) );
  OR2X1 U15718 ( .IN2(n11749), .IN1(n11747), .Q(n11765) );
  OR2X1 U15719 ( .IN2(n11752), .IN1(n11751), .Q(n11756) );
  OR2X1 U15720 ( .IN2(n11754), .IN1(n11753), .Q(n11758) );
  OR2X1 U15721 ( .IN2(n11757), .IN1(n11755), .Q(n11762) );
  OR2X1 U15722 ( .IN2(n11760), .IN1(n11759), .Q(n11764) );
  OR2X1 U15723 ( .IN2(n11763), .IN1(n11761), .Q(n11766) );
  OR2X1 U15724 ( .IN2(n11768), .IN1(n11767), .Q(n11772) );
  OR2X1 U15725 ( .IN2(n11770), .IN1(n11769), .Q(n11774) );
  OR2X1 U15726 ( .IN2(n11773), .IN1(n11771), .Q(n11784) );
  OR2X1 U15727 ( .IN2(n11776), .IN1(n11775), .Q(n11780) );
  OR2X1 U15728 ( .IN2(n11778), .IN1(n11777), .Q(n11782) );
  OR2X1 U15729 ( .IN2(n11781), .IN1(n11779), .Q(n11786) );
  OR2X1 U15730 ( .IN2(n11785), .IN1(n11783), .Q(n11801) );
  OR2X1 U15731 ( .IN2(n11788), .IN1(n11787), .Q(n11792) );
  OR2X1 U15732 ( .IN2(n11790), .IN1(n11789), .Q(n11794) );
  OR2X1 U15733 ( .IN2(n11793), .IN1(n11791), .Q(n11798) );
  OR2X1 U15734 ( .IN2(n11796), .IN1(n11795), .Q(n11800) );
  OR2X1 U15735 ( .IN2(n11799), .IN1(n11797), .Q(n11802) );
  OR2X1 U15736 ( .IN2(n11804), .IN1(n11803), .Q(n11808) );
  OR2X1 U15737 ( .IN2(n11806), .IN1(n11805), .Q(n11810) );
  OR2X1 U15738 ( .IN2(n11809), .IN1(n11807), .Q(n11820) );
  OR2X1 U15739 ( .IN2(n11812), .IN1(n11811), .Q(n11816) );
  OR2X1 U15740 ( .IN2(n11814), .IN1(n11813), .Q(n11818) );
  OR2X1 U15741 ( .IN2(n11817), .IN1(n11815), .Q(n11822) );
  OR2X1 U15742 ( .IN2(n11821), .IN1(n11819), .Q(n11837) );
  OR2X1 U15743 ( .IN2(n11824), .IN1(n11823), .Q(n11828) );
  OR2X1 U15744 ( .IN2(n11826), .IN1(n11825), .Q(n11830) );
  OR2X1 U15745 ( .IN2(n11829), .IN1(n11827), .Q(n11834) );
  OR2X1 U15746 ( .IN2(n11832), .IN1(n11831), .Q(n11836) );
  AND2X1 U15561 ( .IN1(n14399), .IN2(n6869), .Q(n14398) );
  AND2X1 U15562 ( .IN1(n14400), .IN2(n6980), .Q(n11537) );
  AND2X1 U15563 ( .IN1(n14401), .IN2(n6979), .Q(n11538) );
  AND2X1 U15564 ( .IN1(P1_N680), .IN2(n6916), .Q(n14402) );
  AND2X1 U15565 ( .IN1(P1_N680), .IN2(n6915), .Q(n14403) );
  AND2X1 U15566 ( .IN1(P1_N680), .IN2(n6916), .Q(n14404) );
  AND2X1 U15567 ( .IN1(P1_N680), .IN2(n6915), .Q(n14405) );
  AND2X1 U15568 ( .IN1(n14407), .IN2(n6870), .Q(n14406) );
  AND2X1 U15569 ( .IN1(n14409), .IN2(n6869), .Q(n14408) );
  AND2X1 U15570 ( .IN1(P1_N680), .IN2(n6916), .Q(n14410) );
  AND2X1 U15571 ( .IN1(P1_N680), .IN2(n6915), .Q(n14411) );
  AND2X1 U15572 ( .IN1(P1_N680), .IN2(n6916), .Q(n14412) );
  AND2X1 U15573 ( .IN1(P1_N680), .IN2(n6915), .Q(n14413) );
  AND2X1 U15574 ( .IN1(n14415), .IN2(n6870), .Q(n14414) );
  AND2X1 U15575 ( .IN1(n14417), .IN2(n6869), .Q(n14416) );
  AND2X1 U15576 ( .IN1(n14419), .IN2(n6962), .Q(n14418) );
  AND2X1 U15577 ( .IN1(n14421), .IN2(n6949), .Q(n14420) );
  AND2X1 U15578 ( .IN1(P1_N680), .IN2(n6916), .Q(n14422) );
  AND2X1 U15579 ( .IN1(P1_N680), .IN2(n6915), .Q(n14423) );
  AND2X1 U15580 ( .IN1(P1_N680), .IN2(n6916), .Q(n14424) );
  AND2X1 U15581 ( .IN1(P1_N680), .IN2(n6915), .Q(n14425) );
  AND2X1 U15582 ( .IN1(n14427), .IN2(n6870), .Q(n14426) );
  AND2X1 U15583 ( .IN1(n14429), .IN2(n6869), .Q(n14428) );
  AND2X1 U15584 ( .IN1(n14430), .IN2(n6980), .Q(n11539) );
  AND2X1 U15585 ( .IN1(n14431), .IN2(n6979), .Q(n11540) );
  AND2X1 U15586 ( .IN1(P1_N681), .IN2(n6896), .Q(n14432) );
  AND2X1 U15587 ( .IN1(P1_N681), .IN2(n6895), .Q(n14433) );
  AND2X1 U15588 ( .IN1(P1_N681), .IN2(n6896), .Q(n14434) );
  AND2X1 U15589 ( .IN1(P1_N681), .IN2(n6895), .Q(n14435) );
  AND2X1 U15590 ( .IN1(n14437), .IN2(n6870), .Q(n14436) );
  AND2X1 U15591 ( .IN1(n14439), .IN2(n6869), .Q(n14438) );
  AND2X1 U15592 ( .IN1(P1_N681), .IN2(n6896), .Q(n14440) );
  AND2X1 U15593 ( .IN1(P1_N681), .IN2(n6895), .Q(n14441) );
  AND2X1 U15594 ( .IN1(P1_N681), .IN2(n6896), .Q(n14442) );
  AND2X1 U15595 ( .IN1(P1_N681), .IN2(n6895), .Q(n14443) );
  AND2X1 U15596 ( .IN1(n14445), .IN2(n6870), .Q(n14444) );
  AND2X1 U15597 ( .IN1(n14447), .IN2(n6869), .Q(n14446) );
  AND2X1 U15598 ( .IN1(n14449), .IN2(n6958), .Q(n14448) );
  AND2X1 U15599 ( .IN1(n14451), .IN2(n6949), .Q(n14450) );
  AND2X1 U15600 ( .IN1(P1_N681), .IN2(n6896), .Q(n14452) );
  AND2X1 U15601 ( .IN1(P1_N681), .IN2(n6895), .Q(n14453) );
  AND2X1 U15602 ( .IN1(P1_N681), .IN2(n6896), .Q(n14454) );
  AND2X1 U15603 ( .IN1(P1_N681), .IN2(n6895), .Q(n14455) );
  AND2X1 U15604 ( .IN1(n14457), .IN2(n6870), .Q(n14456) );
  AND2X1 U15605 ( .IN1(n14459), .IN2(n6869), .Q(n14458) );
  AND2X1 U15606 ( .IN1(n14460), .IN2(n6980), .Q(n11541) );
  AND2X1 U15607 ( .IN1(n14461), .IN2(n6979), .Q(n11542) );
  AND2X1 U15608 ( .IN1(P1_N682), .IN2(n6896), .Q(n14462) );
  AND2X1 U15609 ( .IN1(P1_N682), .IN2(n6895), .Q(n14463) );
  AND2X1 U15610 ( .IN1(P1_N682), .IN2(n6896), .Q(n14464) );
  AND2X1 U15611 ( .IN1(P1_N682), .IN2(n6895), .Q(n14465) );
  AND2X1 U15612 ( .IN1(n14467), .IN2(n6878), .Q(n14466) );
  AND2X1 U15613 ( .IN1(n14469), .IN2(n6857), .Q(n14468) );
  AND2X1 U15614 ( .IN1(P1_N682), .IN2(n6896), .Q(n14470) );
  AND2X1 U15615 ( .IN1(P1_N682), .IN2(n6895), .Q(n14471) );
  AND2X1 U15616 ( .IN1(P1_N682), .IN2(n6896), .Q(n14472) );
  AND2X1 U15617 ( .IN1(P1_N682), .IN2(n6895), .Q(n14473) );
  AND2X1 U15618 ( .IN1(n14475), .IN2(n6878), .Q(n14474) );
  AND2X1 U15619 ( .IN1(n14477), .IN2(n6857), .Q(n14476) );
  AND2X1 U15620 ( .IN1(n14479), .IN2(n6958), .Q(n14478) );
  AND2X1 U15621 ( .IN1(n14481), .IN2(n6949), .Q(n14480) );
  AND2X1 U15622 ( .IN1(P1_N682), .IN2(n6896), .Q(n14482) );
  AND2X1 U15623 ( .IN1(P1_N682), .IN2(n6895), .Q(n14483) );
  AND2X1 U15624 ( .IN1(P1_N682), .IN2(n6896), .Q(n14484) );
  AND2X1 U15625 ( .IN1(P1_N682), .IN2(n6895), .Q(n14485) );
  AND2X1 U15626 ( .IN1(n14487), .IN2(n6864), .Q(n14486) );
  AND2X1 U15627 ( .IN1(n14489), .IN2(n6857), .Q(n14488) );
  AND2X1 U15628 ( .IN1(n14490), .IN2(n6980), .Q(n11543) );
  AND2X1 U15629 ( .IN1(n14491), .IN2(n6979), .Q(n11544) );
  AND2X1 U15630 ( .IN1(n7019), .IN2(n6896), .Q(n14492) );
  AND2X1 U15631 ( .IN1(n7019), .IN2(n6895), .Q(n14493) );
  AND2X1 U15632 ( .IN1(n7019), .IN2(n6896), .Q(n14494) );
  AND2X1 U15633 ( .IN1(n7019), .IN2(n6895), .Q(n14495) );
  AND2X1 U15634 ( .IN1(n14497), .IN2(n6870), .Q(n14496) );
  AND2X1 U15635 ( .IN1(n14499), .IN2(n6869), .Q(n14498) );
  AND2X1 U15636 ( .IN1(n7028), .IN2(n6910), .Q(n14500) );
  AND2X1 U15637 ( .IN1(n7028), .IN2(n7483), .Q(n14501) );
  AND2X1 U15638 ( .IN1(n7019), .IN2(n6896), .Q(n14502) );
  AND2X1 U15639 ( .IN1(n7019), .IN2(n6895), .Q(n14503) );
  AND2X1 U15640 ( .IN1(n14505), .IN2(n6854), .Q(n14504) );
  AND2X1 U15641 ( .IN1(n14507), .IN2(n6869), .Q(n14506) );
  AND2X1 U15642 ( .IN1(n14509), .IN2(n6952), .Q(n14508) );
  AND2X1 U15643 ( .IN1(n14511), .IN2(n6949), .Q(n14510) );
  AND2X1 U15644 ( .IN1(n14513), .IN2(n14514), .Q(n14512) );
  AND2X1 U15645 ( .IN1(n14516), .IN2(n14517), .Q(n14515) );
  AND2X1 U15646 ( .IN1(n14518), .IN2(n14519), .Q(n11546) );
  AND2X1 U15647 ( .IN1(n14520), .IN2(n6980), .Q(n11547) );
  AND2X1 U15648 ( .IN1(n11545), .IN2(n6979), .Q(n11548) );
  OR2X1 U15650 ( .IN2(n6906), .IN1(P1_N1539), .Q(n13806) );
  OR2X1 U15652 ( .IN2(n11551), .IN1(n11549), .Q(n11561) );
  OR2X1 U15653 ( .IN2(n11553), .IN1(n11552), .Q(n11557) );
  AND2X1 U15468 ( .IN1(P1_N675), .IN2(n6900), .Q(n14272) );
  AND2X1 U15469 ( .IN1(P1_N675), .IN2(n6899), .Q(n14273) );
  AND2X1 U15470 ( .IN1(P1_N675), .IN2(n6900), .Q(n14274) );
  AND2X1 U15471 ( .IN1(P1_N675), .IN2(n6899), .Q(n14275) );
  AND2X1 U15472 ( .IN1(n14277), .IN2(n6856), .Q(n14276) );
  AND2X1 U15473 ( .IN1(n14279), .IN2(n6867), .Q(n14278) );
  AND2X1 U15474 ( .IN1(n14280), .IN2(n6982), .Q(n11529) );
  AND2X1 U15475 ( .IN1(n14281), .IN2(n6981), .Q(n11530) );
  AND2X1 U15476 ( .IN1(P1_N676), .IN2(n6898), .Q(n14282) );
  AND2X1 U15477 ( .IN1(P1_N676), .IN2(n6917), .Q(n14283) );
  AND2X1 U15478 ( .IN1(P1_N676), .IN2(n6916), .Q(n14284) );
  AND2X1 U15479 ( .IN1(P1_N676), .IN2(n6917), .Q(n14285) );
  AND2X1 U15480 ( .IN1(n14287), .IN2(n6862), .Q(n14286) );
  AND2X1 U15481 ( .IN1(n14289), .IN2(n6861), .Q(n14288) );
  AND2X1 U15482 ( .IN1(P1_N676), .IN2(n6894), .Q(n14290) );
  AND2X1 U15483 ( .IN1(P1_N676), .IN2(n6897), .Q(n14291) );
  AND2X1 U15484 ( .IN1(P1_N676), .IN2(n6898), .Q(n14292) );
  AND2X1 U15485 ( .IN1(P1_N676), .IN2(n6917), .Q(n14293) );
  AND2X1 U15486 ( .IN1(n14295), .IN2(n6862), .Q(n14294) );
  AND2X1 U15487 ( .IN1(n14297), .IN2(n6861), .Q(n14296) );
  AND2X1 U15488 ( .IN1(n14299), .IN2(n6956), .Q(n14298) );
  AND2X1 U15489 ( .IN1(n14301), .IN2(n6949), .Q(n14300) );
  AND2X1 U15490 ( .IN1(P1_N676), .IN2(n6916), .Q(n14302) );
  AND2X1 U15491 ( .IN1(P1_N676), .IN2(n6915), .Q(n14303) );
  AND2X1 U15492 ( .IN1(P1_N676), .IN2(n6916), .Q(n14304) );
  AND2X1 U15493 ( .IN1(P1_N676), .IN2(n6915), .Q(n14305) );
  AND2X1 U15494 ( .IN1(n14307), .IN2(n6862), .Q(n14306) );
  AND2X1 U15495 ( .IN1(n14309), .IN2(n6867), .Q(n14308) );
  AND2X1 U15496 ( .IN1(n14310), .IN2(n6982), .Q(n11531) );
  AND2X1 U15497 ( .IN1(n14311), .IN2(n6981), .Q(n11532) );
  AND2X1 U15498 ( .IN1(P1_N677), .IN2(n6916), .Q(n14312) );
  AND2X1 U15499 ( .IN1(P1_N677), .IN2(n6915), .Q(n14313) );
  AND2X1 U15500 ( .IN1(P1_N677), .IN2(n6916), .Q(n14314) );
  AND2X1 U15501 ( .IN1(P1_N677), .IN2(n6915), .Q(n14315) );
  AND2X1 U15502 ( .IN1(n14317), .IN2(n6862), .Q(n14316) );
  AND2X1 U15503 ( .IN1(n14319), .IN2(n6861), .Q(n14318) );
  AND2X1 U15504 ( .IN1(P1_N677), .IN2(n6916), .Q(n14320) );
  AND2X1 U15505 ( .IN1(P1_N677), .IN2(n6915), .Q(n14321) );
  AND2X1 U15506 ( .IN1(P1_N677), .IN2(n6916), .Q(n14322) );
  AND2X1 U15507 ( .IN1(P1_N677), .IN2(n6915), .Q(n14323) );
  AND2X1 U15508 ( .IN1(n14325), .IN2(n6878), .Q(n14324) );
  AND2X1 U15509 ( .IN1(n14327), .IN2(n6867), .Q(n14326) );
  AND2X1 U15510 ( .IN1(n14329), .IN2(n6956), .Q(n14328) );
  AND2X1 U15511 ( .IN1(n14331), .IN2(n6949), .Q(n14330) );
  AND2X1 U15512 ( .IN1(P1_N677), .IN2(n6916), .Q(n14332) );
  AND2X1 U15513 ( .IN1(P1_N677), .IN2(n6915), .Q(n14333) );
  AND2X1 U15514 ( .IN1(P1_N677), .IN2(n6916), .Q(n14334) );
  AND2X1 U15515 ( .IN1(P1_N677), .IN2(n6915), .Q(n14335) );
  AND2X1 U15516 ( .IN1(n14337), .IN2(n6862), .Q(n14336) );
  AND2X1 U15517 ( .IN1(n14339), .IN2(n6867), .Q(n14338) );
  AND2X1 U15518 ( .IN1(n14340), .IN2(n6982), .Q(n11533) );
  AND2X1 U15519 ( .IN1(n14341), .IN2(n6981), .Q(n11534) );
  AND2X1 U15520 ( .IN1(P1_N678), .IN2(n6916), .Q(n14342) );
  AND2X1 U15521 ( .IN1(P1_N678), .IN2(n6915), .Q(n14343) );
  AND2X1 U15522 ( .IN1(P1_N678), .IN2(n6916), .Q(n14344) );
  AND2X1 U15523 ( .IN1(P1_N678), .IN2(n6915), .Q(n14345) );
  AND2X1 U15524 ( .IN1(n14347), .IN2(n6878), .Q(n14346) );
  AND2X1 U15525 ( .IN1(n14349), .IN2(n6867), .Q(n14348) );
  AND2X1 U15526 ( .IN1(P1_N678), .IN2(n6916), .Q(n14350) );
  AND2X1 U15527 ( .IN1(P1_N678), .IN2(n6915), .Q(n14351) );
  AND2X1 U15528 ( .IN1(P1_N678), .IN2(n6916), .Q(n14352) );
  AND2X1 U15529 ( .IN1(P1_N678), .IN2(n6915), .Q(n14353) );
  AND2X1 U15530 ( .IN1(n14355), .IN2(n6878), .Q(n14354) );
  AND2X1 U15531 ( .IN1(n14357), .IN2(n6867), .Q(n14356) );
  AND2X1 U15532 ( .IN1(n14359), .IN2(n6956), .Q(n14358) );
  AND2X1 U15533 ( .IN1(n14361), .IN2(n6949), .Q(n14360) );
  AND2X1 U15534 ( .IN1(P1_N678), .IN2(n6916), .Q(n14362) );
  AND2X1 U15535 ( .IN1(P1_N678), .IN2(n6915), .Q(n14363) );
  AND2X1 U15536 ( .IN1(P1_N678), .IN2(n6916), .Q(n14364) );
  AND2X1 U15537 ( .IN1(P1_N678), .IN2(n6915), .Q(n14365) );
  AND2X1 U15538 ( .IN1(n14367), .IN2(n6878), .Q(n14366) );
  AND2X1 U15539 ( .IN1(n14369), .IN2(n6867), .Q(n14368) );
  AND2X1 U15540 ( .IN1(n14370), .IN2(n6982), .Q(n11535) );
  AND2X1 U15541 ( .IN1(n14371), .IN2(n6981), .Q(n11536) );
  AND2X1 U15542 ( .IN1(P1_N679), .IN2(n6916), .Q(n14372) );
  AND2X1 U15543 ( .IN1(P1_N679), .IN2(n6915), .Q(n14373) );
  AND2X1 U15544 ( .IN1(P1_N679), .IN2(n6916), .Q(n14374) );
  AND2X1 U15545 ( .IN1(P1_N679), .IN2(n6915), .Q(n14375) );
  AND2X1 U15546 ( .IN1(n14377), .IN2(n6870), .Q(n14376) );
  AND2X1 U15547 ( .IN1(n14379), .IN2(n6869), .Q(n14378) );
  AND2X1 U15548 ( .IN1(P1_N679), .IN2(n6916), .Q(n14380) );
  AND2X1 U15549 ( .IN1(P1_N679), .IN2(n6915), .Q(n14381) );
  AND2X1 U15550 ( .IN1(P1_N679), .IN2(n6916), .Q(n14382) );
  AND2X1 U15551 ( .IN1(P1_N679), .IN2(n6915), .Q(n14383) );
  AND2X1 U15552 ( .IN1(n14385), .IN2(n6870), .Q(n14384) );
  AND2X1 U15553 ( .IN1(n14387), .IN2(n6869), .Q(n14386) );
  AND2X1 U15554 ( .IN1(n14389), .IN2(n6962), .Q(n14388) );
  AND2X1 U15555 ( .IN1(n14391), .IN2(n6949), .Q(n14390) );
  AND2X1 U15556 ( .IN1(P1_N679), .IN2(n6916), .Q(n14392) );
  AND2X1 U15557 ( .IN1(P1_N679), .IN2(n6915), .Q(n14393) );
  AND2X1 U15558 ( .IN1(P1_N679), .IN2(n6916), .Q(n14394) );
  AND2X1 U15559 ( .IN1(P1_N679), .IN2(n6915), .Q(n14395) );
  AND2X1 U15560 ( .IN1(n14397), .IN2(n6870), .Q(n14396) );
  AND2X1 U15375 ( .IN1(P1_N671), .IN2(n6899), .Q(n14143) );
  AND2X1 U15376 ( .IN1(n14145), .IN2(n6862), .Q(n14144) );
  AND2X1 U15377 ( .IN1(n14147), .IN2(n6867), .Q(n14146) );
  AND2X1 U15378 ( .IN1(n14149), .IN2(n6962), .Q(n14148) );
  AND2X1 U15379 ( .IN1(n14151), .IN2(n6961), .Q(n14150) );
  AND2X1 U15380 ( .IN1(P1_N671), .IN2(n6884), .Q(n14152) );
  AND2X1 U15381 ( .IN1(P1_N671), .IN2(n6917), .Q(n14153) );
  AND2X1 U15382 ( .IN1(P1_N671), .IN2(n6884), .Q(n14154) );
  AND2X1 U15383 ( .IN1(P1_N671), .IN2(n6917), .Q(n14155) );
  AND2X1 U15384 ( .IN1(n14157), .IN2(n6856), .Q(n14156) );
  AND2X1 U15385 ( .IN1(n14159), .IN2(n6861), .Q(n14158) );
  AND2X1 U15386 ( .IN1(n14160), .IN2(n6982), .Q(n11521) );
  AND2X1 U15387 ( .IN1(n14161), .IN2(n6981), .Q(n11522) );
  AND2X1 U15388 ( .IN1(P1_N672), .IN2(n6900), .Q(n14162) );
  AND2X1 U15389 ( .IN1(P1_N672), .IN2(n6899), .Q(n14163) );
  AND2X1 U15390 ( .IN1(P1_N672), .IN2(n6900), .Q(n14164) );
  AND2X1 U15391 ( .IN1(P1_N672), .IN2(n6899), .Q(n14165) );
  AND2X1 U15392 ( .IN1(n14167), .IN2(n6878), .Q(n14166) );
  AND2X1 U15393 ( .IN1(n14169), .IN2(n6867), .Q(n14168) );
  AND2X1 U15394 ( .IN1(P1_N672), .IN2(n6900), .Q(n14170) );
  AND2X1 U15395 ( .IN1(P1_N672), .IN2(n6899), .Q(n14171) );
  AND2X1 U15396 ( .IN1(P1_N672), .IN2(n6900), .Q(n14172) );
  AND2X1 U15397 ( .IN1(P1_N672), .IN2(n6899), .Q(n14173) );
  AND2X1 U15398 ( .IN1(n14175), .IN2(n6878), .Q(n14174) );
  AND2X1 U15399 ( .IN1(n14177), .IN2(n6867), .Q(n14176) );
  AND2X1 U15400 ( .IN1(n14179), .IN2(n6962), .Q(n14178) );
  AND2X1 U15401 ( .IN1(n14181), .IN2(n6961), .Q(n14180) );
  AND2X1 U15402 ( .IN1(P1_N672), .IN2(n6900), .Q(n14182) );
  AND2X1 U15403 ( .IN1(P1_N672), .IN2(n6899), .Q(n14183) );
  AND2X1 U15404 ( .IN1(P1_N672), .IN2(n6900), .Q(n14184) );
  AND2X1 U15405 ( .IN1(P1_N672), .IN2(n6899), .Q(n14185) );
  AND2X1 U15406 ( .IN1(n14187), .IN2(n6856), .Q(n14186) );
  AND2X1 U15407 ( .IN1(n14189), .IN2(n6867), .Q(n14188) );
  AND2X1 U15408 ( .IN1(n14190), .IN2(n6982), .Q(n11523) );
  AND2X1 U15409 ( .IN1(n14191), .IN2(n6981), .Q(n11524) );
  AND2X1 U15410 ( .IN1(P1_N673), .IN2(n6900), .Q(n14192) );
  AND2X1 U15411 ( .IN1(P1_N673), .IN2(n6899), .Q(n14193) );
  AND2X1 U15412 ( .IN1(P1_N673), .IN2(n6900), .Q(n14194) );
  AND2X1 U15413 ( .IN1(P1_N673), .IN2(n6899), .Q(n14195) );
  AND2X1 U15414 ( .IN1(n14197), .IN2(n6862), .Q(n14196) );
  AND2X1 U15415 ( .IN1(n14199), .IN2(n6867), .Q(n14198) );
  AND2X1 U15416 ( .IN1(P1_N673), .IN2(n6900), .Q(n14200) );
  AND2X1 U15417 ( .IN1(P1_N673), .IN2(n6899), .Q(n14201) );
  AND2X1 U15418 ( .IN1(P1_N673), .IN2(n6900), .Q(n14202) );
  AND2X1 U15419 ( .IN1(P1_N673), .IN2(n6899), .Q(n14203) );
  AND2X1 U15420 ( .IN1(n14205), .IN2(n6862), .Q(n14204) );
  AND2X1 U15421 ( .IN1(n14207), .IN2(n6867), .Q(n14206) );
  AND2X1 U15422 ( .IN1(n14209), .IN2(n6962), .Q(n14208) );
  AND2X1 U15423 ( .IN1(n14211), .IN2(n6961), .Q(n14210) );
  AND2X1 U15424 ( .IN1(P1_N673), .IN2(n6900), .Q(n14212) );
  AND2X1 U15425 ( .IN1(P1_N673), .IN2(n6899), .Q(n14213) );
  AND2X1 U15426 ( .IN1(P1_N673), .IN2(n6900), .Q(n14214) );
  AND2X1 U15427 ( .IN1(P1_N673), .IN2(n6899), .Q(n14215) );
  AND2X1 U15428 ( .IN1(n14217), .IN2(n6862), .Q(n14216) );
  AND2X1 U15429 ( .IN1(n14219), .IN2(n6867), .Q(n14218) );
  AND2X1 U15430 ( .IN1(n14220), .IN2(n6982), .Q(n11525) );
  AND2X1 U15431 ( .IN1(n14221), .IN2(n6981), .Q(n11526) );
  AND2X1 U15432 ( .IN1(P1_N674), .IN2(n6900), .Q(n14222) );
  AND2X1 U15433 ( .IN1(P1_N674), .IN2(n6899), .Q(n14223) );
  AND2X1 U15434 ( .IN1(P1_N674), .IN2(n6900), .Q(n14224) );
  AND2X1 U15435 ( .IN1(P1_N674), .IN2(n6899), .Q(n14225) );
  AND2X1 U15436 ( .IN1(n14227), .IN2(n6862), .Q(n14226) );
  AND2X1 U15437 ( .IN1(n14229), .IN2(n6867), .Q(n14228) );
  AND2X1 U15438 ( .IN1(P1_N674), .IN2(n6900), .Q(n14230) );
  AND2X1 U15439 ( .IN1(P1_N674), .IN2(n6899), .Q(n14231) );
  AND2X1 U15440 ( .IN1(P1_N674), .IN2(n6900), .Q(n14232) );
  AND2X1 U15441 ( .IN1(P1_N674), .IN2(n6899), .Q(n14233) );
  AND2X1 U15442 ( .IN1(n14235), .IN2(n6862), .Q(n14234) );
  AND2X1 U15443 ( .IN1(n14237), .IN2(n6867), .Q(n14236) );
  AND2X1 U15444 ( .IN1(n14239), .IN2(n6962), .Q(n14238) );
  AND2X1 U15445 ( .IN1(n14241), .IN2(n6961), .Q(n14240) );
  AND2X1 U15446 ( .IN1(P1_N674), .IN2(n6900), .Q(n14242) );
  AND2X1 U15447 ( .IN1(P1_N674), .IN2(n6899), .Q(n14243) );
  AND2X1 U15448 ( .IN1(P1_N674), .IN2(n6900), .Q(n14244) );
  AND2X1 U15449 ( .IN1(P1_N674), .IN2(n6899), .Q(n14245) );
  AND2X1 U15450 ( .IN1(n14247), .IN2(n6862), .Q(n14246) );
  AND2X1 U15451 ( .IN1(n14249), .IN2(n6867), .Q(n14248) );
  AND2X1 U15452 ( .IN1(n14250), .IN2(n6982), .Q(n11527) );
  AND2X1 U15453 ( .IN1(n14251), .IN2(n6981), .Q(n11528) );
  AND2X1 U15454 ( .IN1(P1_N675), .IN2(n6900), .Q(n14252) );
  AND2X1 U15455 ( .IN1(P1_N675), .IN2(n6899), .Q(n14253) );
  AND2X1 U15456 ( .IN1(P1_N675), .IN2(n6900), .Q(n14254) );
  AND2X1 U15457 ( .IN1(P1_N675), .IN2(n6899), .Q(n14255) );
  AND2X1 U15458 ( .IN1(n14257), .IN2(n6878), .Q(n14256) );
  AND2X1 U15459 ( .IN1(n14259), .IN2(n6867), .Q(n14258) );
  AND2X1 U15460 ( .IN1(P1_N675), .IN2(n6900), .Q(n14260) );
  AND2X1 U15461 ( .IN1(P1_N675), .IN2(n6899), .Q(n14261) );
  AND2X1 U15462 ( .IN1(P1_N675), .IN2(n6900), .Q(n14262) );
  AND2X1 U15463 ( .IN1(P1_N675), .IN2(n6899), .Q(n14263) );
  AND2X1 U15464 ( .IN1(n14265), .IN2(n6862), .Q(n14264) );
  AND2X1 U15465 ( .IN1(n14267), .IN2(n6867), .Q(n14266) );
  AND2X1 U15466 ( .IN1(n14269), .IN2(n6962), .Q(n14268) );
  AND2X1 U15467 ( .IN1(n14271), .IN2(n6961), .Q(n14270) );
  AND2X1 U15282 ( .IN1(n14017), .IN2(n6862), .Q(n14016) );
  AND2X1 U15283 ( .IN1(n14019), .IN2(n6861), .Q(n14018) );
  AND2X1 U15284 ( .IN1(P1_N667), .IN2(n6898), .Q(n14020) );
  AND2X1 U15285 ( .IN1(P1_N667), .IN2(n6897), .Q(n14021) );
  AND2X1 U15286 ( .IN1(P1_N667), .IN2(n6898), .Q(n14022) );
  AND2X1 U15287 ( .IN1(P1_N667), .IN2(n6897), .Q(n14023) );
  AND2X1 U15288 ( .IN1(n14025), .IN2(n6862), .Q(n14024) );
  AND2X1 U15289 ( .IN1(n14027), .IN2(n6861), .Q(n14026) );
  AND2X1 U15290 ( .IN1(n14029), .IN2(n6962), .Q(n14028) );
  AND2X1 U15291 ( .IN1(n14031), .IN2(n6961), .Q(n14030) );
  AND2X1 U15292 ( .IN1(P1_N667), .IN2(n6884), .Q(n14032) );
  AND2X1 U15293 ( .IN1(P1_N667), .IN2(n6917), .Q(n14033) );
  AND2X1 U15294 ( .IN1(P1_N667), .IN2(n6884), .Q(n14034) );
  AND2X1 U15295 ( .IN1(P1_N667), .IN2(n6897), .Q(n14035) );
  AND2X1 U15296 ( .IN1(n14037), .IN2(n6862), .Q(n14036) );
  AND2X1 U15297 ( .IN1(n14039), .IN2(n6861), .Q(n14038) );
  AND2X1 U15298 ( .IN1(n14040), .IN2(n6982), .Q(n11513) );
  AND2X1 U15299 ( .IN1(n14041), .IN2(n6981), .Q(n11514) );
  AND2X1 U15300 ( .IN1(P1_N668), .IN2(n6900), .Q(n14042) );
  AND2X1 U15301 ( .IN1(P1_N668), .IN2(n6917), .Q(n14043) );
  AND2X1 U15302 ( .IN1(P1_N668), .IN2(n6898), .Q(n14044) );
  AND2X1 U15303 ( .IN1(P1_N668), .IN2(n6917), .Q(n14045) );
  AND2X1 U15304 ( .IN1(n14047), .IN2(n6862), .Q(n14046) );
  AND2X1 U15305 ( .IN1(n14049), .IN2(n6861), .Q(n14048) );
  AND2X1 U15306 ( .IN1(P1_N668), .IN2(n6900), .Q(n14050) );
  AND2X1 U15307 ( .IN1(P1_N668), .IN2(n6917), .Q(n14051) );
  AND2X1 U15308 ( .IN1(P1_N668), .IN2(n6916), .Q(n14052) );
  AND2X1 U15309 ( .IN1(P1_N668), .IN2(n6917), .Q(n14053) );
  AND2X1 U15310 ( .IN1(n14055), .IN2(n6862), .Q(n14054) );
  AND2X1 U15311 ( .IN1(n14057), .IN2(n6861), .Q(n14056) );
  AND2X1 U15312 ( .IN1(n14059), .IN2(n6962), .Q(n14058) );
  AND2X1 U15313 ( .IN1(n14061), .IN2(n6961), .Q(n14060) );
  AND2X1 U15314 ( .IN1(P1_N668), .IN2(n6884), .Q(n14062) );
  AND2X1 U15315 ( .IN1(P1_N668), .IN2(n6917), .Q(n14063) );
  AND2X1 U15316 ( .IN1(P1_N668), .IN2(n6884), .Q(n14064) );
  AND2X1 U15317 ( .IN1(P1_N668), .IN2(n6917), .Q(n14065) );
  AND2X1 U15318 ( .IN1(n14067), .IN2(n6862), .Q(n14066) );
  AND2X1 U15319 ( .IN1(n14069), .IN2(n6861), .Q(n14068) );
  AND2X1 U15320 ( .IN1(n14070), .IN2(n6982), .Q(n11515) );
  AND2X1 U15321 ( .IN1(n14071), .IN2(n6981), .Q(n11516) );
  AND2X1 U15322 ( .IN1(P1_N669), .IN2(n6900), .Q(n14072) );
  AND2X1 U15323 ( .IN1(P1_N669), .IN2(n6917), .Q(n14073) );
  AND2X1 U15324 ( .IN1(P1_N669), .IN2(n6894), .Q(n14074) );
  AND2X1 U15325 ( .IN1(P1_N669), .IN2(n6917), .Q(n14075) );
  AND2X1 U15326 ( .IN1(n14077), .IN2(n6862), .Q(n14076) );
  AND2X1 U15327 ( .IN1(n14079), .IN2(n6861), .Q(n14078) );
  AND2X1 U15328 ( .IN1(P1_N669), .IN2(n6916), .Q(n14080) );
  AND2X1 U15329 ( .IN1(P1_N669), .IN2(n6917), .Q(n14081) );
  AND2X1 U15330 ( .IN1(P1_N669), .IN2(n6916), .Q(n14082) );
  AND2X1 U15331 ( .IN1(P1_N669), .IN2(n6917), .Q(n14083) );
  AND2X1 U15332 ( .IN1(n14085), .IN2(n6862), .Q(n14084) );
  AND2X1 U15333 ( .IN1(n14087), .IN2(n6861), .Q(n14086) );
  AND2X1 U15334 ( .IN1(n14089), .IN2(n6962), .Q(n14088) );
  AND2X1 U15335 ( .IN1(n14091), .IN2(n6961), .Q(n14090) );
  AND2X1 U15336 ( .IN1(P1_N669), .IN2(n6884), .Q(n14092) );
  AND2X1 U15337 ( .IN1(P1_N669), .IN2(n6917), .Q(n14093) );
  AND2X1 U15338 ( .IN1(P1_N669), .IN2(n6884), .Q(n14094) );
  AND2X1 U15339 ( .IN1(P1_N669), .IN2(n6917), .Q(n14095) );
  AND2X1 U15340 ( .IN1(n14097), .IN2(n6862), .Q(n14096) );
  AND2X1 U15341 ( .IN1(n14099), .IN2(n6861), .Q(n14098) );
  AND2X1 U15342 ( .IN1(n14100), .IN2(n6982), .Q(n11517) );
  AND2X1 U15343 ( .IN1(n14101), .IN2(n6981), .Q(n11518) );
  AND2X1 U15344 ( .IN1(P1_N670), .IN2(n6916), .Q(n14102) );
  AND2X1 U15345 ( .IN1(P1_N670), .IN2(n6917), .Q(n14103) );
  AND2X1 U15346 ( .IN1(P1_N670), .IN2(n6898), .Q(n14104) );
  AND2X1 U15347 ( .IN1(P1_N670), .IN2(n6917), .Q(n14105) );
  AND2X1 U15348 ( .IN1(n14107), .IN2(n6862), .Q(n14106) );
  AND2X1 U15349 ( .IN1(n14109), .IN2(n6861), .Q(n14108) );
  AND2X1 U15350 ( .IN1(P1_N670), .IN2(n6900), .Q(n14110) );
  AND2X1 U15351 ( .IN1(P1_N670), .IN2(n6917), .Q(n14111) );
  AND2X1 U15352 ( .IN1(P1_N670), .IN2(n6900), .Q(n14112) );
  AND2X1 U15353 ( .IN1(P1_N670), .IN2(n6917), .Q(n14113) );
  AND2X1 U15354 ( .IN1(n14115), .IN2(n6862), .Q(n14114) );
  AND2X1 U15355 ( .IN1(n14117), .IN2(n6861), .Q(n14116) );
  AND2X1 U15356 ( .IN1(n14119), .IN2(n6962), .Q(n14118) );
  AND2X1 U15357 ( .IN1(n14121), .IN2(n6961), .Q(n14120) );
  AND2X1 U15358 ( .IN1(P1_N670), .IN2(n6884), .Q(n14122) );
  AND2X1 U15359 ( .IN1(P1_N670), .IN2(n6917), .Q(n14123) );
  AND2X1 U15360 ( .IN1(P1_N670), .IN2(n6884), .Q(n14124) );
  AND2X1 U15361 ( .IN1(P1_N670), .IN2(n6917), .Q(n14125) );
  AND2X1 U15362 ( .IN1(n14127), .IN2(n6862), .Q(n14126) );
  AND2X1 U15363 ( .IN1(n14129), .IN2(n6861), .Q(n14128) );
  AND2X1 U15364 ( .IN1(n14130), .IN2(n6982), .Q(n11519) );
  AND2X1 U15365 ( .IN1(n14131), .IN2(n6981), .Q(n11520) );
  AND2X1 U15366 ( .IN1(P1_N671), .IN2(n6916), .Q(n14132) );
  AND2X1 U15367 ( .IN1(P1_N671), .IN2(n6917), .Q(n14133) );
  AND2X1 U15368 ( .IN1(P1_N671), .IN2(n6916), .Q(n14134) );
  AND2X1 U15369 ( .IN1(P1_N671), .IN2(n6917), .Q(n14135) );
  AND2X1 U15370 ( .IN1(n14137), .IN2(n6862), .Q(n14136) );
  AND2X1 U15371 ( .IN1(n14139), .IN2(n6861), .Q(n14138) );
  AND2X1 U15372 ( .IN1(P1_N671), .IN2(n6900), .Q(n14140) );
  AND2X1 U15373 ( .IN1(P1_N671), .IN2(n6917), .Q(n14141) );
  AND2X1 U15374 ( .IN1(P1_N671), .IN2(n6900), .Q(n14142) );
  AND2X1 U15189 ( .IN1(n13891), .IN2(n6977), .Q(n11504) );
  AND2X1 U15190 ( .IN1(P1_N663), .IN2(n6898), .Q(n13892) );
  AND2X1 U15191 ( .IN1(P1_N663), .IN2(n6897), .Q(n13893) );
  AND2X1 U15192 ( .IN1(P1_N663), .IN2(n6898), .Q(n13894) );
  AND2X1 U15193 ( .IN1(P1_N663), .IN2(n6897), .Q(n13895) );
  AND2X1 U15194 ( .IN1(n13897), .IN2(n6862), .Q(n13896) );
  AND2X1 U15195 ( .IN1(n13899), .IN2(n6861), .Q(n13898) );
  AND2X1 U15196 ( .IN1(P1_N663), .IN2(n6898), .Q(n13900) );
  AND2X1 U15197 ( .IN1(P1_N663), .IN2(n6897), .Q(n13901) );
  AND2X1 U15198 ( .IN1(P1_N663), .IN2(n6898), .Q(n13902) );
  AND2X1 U15199 ( .IN1(P1_N663), .IN2(n6897), .Q(n13903) );
  AND2X1 U15200 ( .IN1(n13905), .IN2(n6862), .Q(n13904) );
  AND2X1 U15201 ( .IN1(n13907), .IN2(n6861), .Q(n13906) );
  AND2X1 U15202 ( .IN1(n13909), .IN2(n6956), .Q(n13908) );
  AND2X1 U15203 ( .IN1(n13911), .IN2(n6949), .Q(n13910) );
  AND2X1 U15204 ( .IN1(P1_N663), .IN2(n6898), .Q(n13912) );
  AND2X1 U15205 ( .IN1(P1_N663), .IN2(n6897), .Q(n13913) );
  AND2X1 U15206 ( .IN1(P1_N663), .IN2(n6898), .Q(n13914) );
  AND2X1 U15207 ( .IN1(P1_N663), .IN2(n6897), .Q(n13915) );
  AND2X1 U15208 ( .IN1(n13917), .IN2(n6862), .Q(n13916) );
  AND2X1 U15209 ( .IN1(n13919), .IN2(n6861), .Q(n13918) );
  AND2X1 U15210 ( .IN1(n13920), .IN2(n6980), .Q(n11505) );
  AND2X1 U15211 ( .IN1(n13921), .IN2(n6979), .Q(n11506) );
  AND2X1 U15212 ( .IN1(P1_N664), .IN2(n6898), .Q(n13922) );
  AND2X1 U15213 ( .IN1(P1_N664), .IN2(n6897), .Q(n13923) );
  AND2X1 U15214 ( .IN1(P1_N664), .IN2(n6898), .Q(n13924) );
  AND2X1 U15215 ( .IN1(P1_N664), .IN2(n6897), .Q(n13925) );
  AND2X1 U15216 ( .IN1(n13927), .IN2(n6862), .Q(n13926) );
  AND2X1 U15217 ( .IN1(n13929), .IN2(n6861), .Q(n13928) );
  AND2X1 U15218 ( .IN1(P1_N664), .IN2(n6898), .Q(n13930) );
  AND2X1 U15219 ( .IN1(P1_N664), .IN2(n6897), .Q(n13931) );
  AND2X1 U15220 ( .IN1(P1_N664), .IN2(n6898), .Q(n13932) );
  AND2X1 U15221 ( .IN1(P1_N664), .IN2(n6897), .Q(n13933) );
  AND2X1 U15222 ( .IN1(n13935), .IN2(n6862), .Q(n13934) );
  AND2X1 U15223 ( .IN1(n13937), .IN2(n6861), .Q(n13936) );
  AND2X1 U15224 ( .IN1(n13939), .IN2(n6956), .Q(n13938) );
  AND2X1 U15225 ( .IN1(n13941), .IN2(n6949), .Q(n13940) );
  AND2X1 U15226 ( .IN1(P1_N664), .IN2(n6898), .Q(n13942) );
  AND2X1 U15227 ( .IN1(P1_N664), .IN2(n6897), .Q(n13943) );
  AND2X1 U15228 ( .IN1(P1_N664), .IN2(n6898), .Q(n13944) );
  AND2X1 U15229 ( .IN1(P1_N664), .IN2(n6897), .Q(n13945) );
  AND2X1 U15230 ( .IN1(n13947), .IN2(n6862), .Q(n13946) );
  AND2X1 U15231 ( .IN1(n13949), .IN2(n6861), .Q(n13948) );
  AND2X1 U15232 ( .IN1(n13950), .IN2(n6980), .Q(n11507) );
  AND2X1 U15233 ( .IN1(n13951), .IN2(n6979), .Q(n11508) );
  AND2X1 U15234 ( .IN1(P1_N665), .IN2(n6898), .Q(n13952) );
  AND2X1 U15235 ( .IN1(P1_N665), .IN2(n6897), .Q(n13953) );
  AND2X1 U15236 ( .IN1(P1_N665), .IN2(n6898), .Q(n13954) );
  AND2X1 U15237 ( .IN1(P1_N665), .IN2(n6897), .Q(n13955) );
  AND2X1 U15238 ( .IN1(n13957), .IN2(n6862), .Q(n13956) );
  AND2X1 U15239 ( .IN1(n13959), .IN2(n6861), .Q(n13958) );
  AND2X1 U15240 ( .IN1(P1_N665), .IN2(n6898), .Q(n13960) );
  AND2X1 U15241 ( .IN1(P1_N665), .IN2(n6897), .Q(n13961) );
  AND2X1 U15242 ( .IN1(P1_N665), .IN2(n6898), .Q(n13962) );
  AND2X1 U15243 ( .IN1(P1_N665), .IN2(n6897), .Q(n13963) );
  AND2X1 U15244 ( .IN1(n13965), .IN2(n6862), .Q(n13964) );
  AND2X1 U15245 ( .IN1(n13967), .IN2(n6861), .Q(n13966) );
  AND2X1 U15246 ( .IN1(n13969), .IN2(n6962), .Q(n13968) );
  AND2X1 U15247 ( .IN1(n13971), .IN2(n6961), .Q(n13970) );
  AND2X1 U15248 ( .IN1(P1_N665), .IN2(n6898), .Q(n13972) );
  AND2X1 U15249 ( .IN1(P1_N665), .IN2(n6897), .Q(n13973) );
  AND2X1 U15250 ( .IN1(P1_N665), .IN2(n6898), .Q(n13974) );
  AND2X1 U15251 ( .IN1(P1_N665), .IN2(n6897), .Q(n13975) );
  AND2X1 U15252 ( .IN1(n13977), .IN2(n6862), .Q(n13976) );
  AND2X1 U15253 ( .IN1(n13979), .IN2(n6861), .Q(n13978) );
  AND2X1 U15254 ( .IN1(n13980), .IN2(n6982), .Q(n11509) );
  AND2X1 U15255 ( .IN1(n13981), .IN2(n6981), .Q(n11510) );
  AND2X1 U15256 ( .IN1(P1_N666), .IN2(n6898), .Q(n13982) );
  AND2X1 U15257 ( .IN1(P1_N666), .IN2(n6897), .Q(n13983) );
  AND2X1 U15258 ( .IN1(P1_N666), .IN2(n6898), .Q(n13984) );
  AND2X1 U15259 ( .IN1(P1_N666), .IN2(n6897), .Q(n13985) );
  AND2X1 U15260 ( .IN1(n13987), .IN2(n6862), .Q(n13986) );
  AND2X1 U15261 ( .IN1(n13989), .IN2(n6861), .Q(n13988) );
  AND2X1 U15262 ( .IN1(P1_N666), .IN2(n6898), .Q(n13990) );
  AND2X1 U15263 ( .IN1(P1_N666), .IN2(n6897), .Q(n13991) );
  AND2X1 U15264 ( .IN1(P1_N666), .IN2(n6898), .Q(n13992) );
  AND2X1 U15265 ( .IN1(P1_N666), .IN2(n6897), .Q(n13993) );
  AND2X1 U15266 ( .IN1(n13995), .IN2(n6862), .Q(n13994) );
  AND2X1 U15267 ( .IN1(n13997), .IN2(n6861), .Q(n13996) );
  AND2X1 U15268 ( .IN1(n13999), .IN2(n6962), .Q(n13998) );
  AND2X1 U15269 ( .IN1(n14001), .IN2(n6961), .Q(n14000) );
  AND2X1 U15270 ( .IN1(P1_N666), .IN2(n6898), .Q(n14002) );
  AND2X1 U15271 ( .IN1(P1_N666), .IN2(n6897), .Q(n14003) );
  AND2X1 U15272 ( .IN1(P1_N666), .IN2(n6898), .Q(n14004) );
  AND2X1 U15273 ( .IN1(P1_N666), .IN2(n6897), .Q(n14005) );
  AND2X1 U15274 ( .IN1(n14007), .IN2(n6862), .Q(n14006) );
  AND2X1 U15275 ( .IN1(n14009), .IN2(n6861), .Q(n14008) );
  AND2X1 U15276 ( .IN1(n14010), .IN2(n6982), .Q(n11511) );
  AND2X1 U15277 ( .IN1(n14011), .IN2(n6981), .Q(n11512) );
  AND2X1 U15278 ( .IN1(P1_N667), .IN2(n6898), .Q(n14012) );
  AND2X1 U15279 ( .IN1(P1_N667), .IN2(n6897), .Q(n14013) );
  AND2X1 U15280 ( .IN1(P1_N667), .IN2(n6898), .Q(n14014) );
  AND2X1 U15281 ( .IN1(P1_N667), .IN2(n6897), .Q(n14015) );
  AND2X1 U15096 ( .IN1(n13475), .IN2(n6957), .Q(n13773) );
  AND2X1 U15097 ( .IN1(n13775), .IN2(n6952), .Q(n13774) );
  AND2X1 U15098 ( .IN1(n13488), .IN2(n6977), .Q(n11483) );
  AND2X1 U15099 ( .IN1(n13776), .IN2(n6982), .Q(n11484) );
  AND2X1 U15100 ( .IN1(P1_N1383), .IN2(n6855), .Q(n13777) );
  AND2X1 U15101 ( .IN1(n13494), .IN2(n6856), .Q(n13778) );
  AND2X1 U15102 ( .IN1(n13508), .IN2(n6959), .Q(n13779) );
  AND2X1 U15103 ( .IN1(n13781), .IN2(n6952), .Q(n13780) );
  AND2X1 U15104 ( .IN1(n13521), .IN2(n6977), .Q(n11485) );
  AND2X1 U15105 ( .IN1(n13782), .IN2(n6980), .Q(n11486) );
  AND2X1 U15106 ( .IN1(P1_N1384), .IN2(n6855), .Q(n13783) );
  AND2X1 U15107 ( .IN1(n13527), .IN2(n6856), .Q(n13784) );
  AND2X1 U15108 ( .IN1(n13541), .IN2(n6959), .Q(n13785) );
  AND2X1 U15109 ( .IN1(n13787), .IN2(n6952), .Q(n13786) );
  AND2X1 U15110 ( .IN1(n13554), .IN2(n6977), .Q(n11487) );
  AND2X1 U15111 ( .IN1(n13788), .IN2(n6984), .Q(n11488) );
  AND2X1 U15112 ( .IN1(P1_N1385), .IN2(n6855), .Q(n13789) );
  AND2X1 U15113 ( .IN1(n13560), .IN2(n6866), .Q(n13790) );
  AND2X1 U15114 ( .IN1(n13574), .IN2(n6955), .Q(n13791) );
  AND2X1 U15115 ( .IN1(n13793), .IN2(n6952), .Q(n13792) );
  AND2X1 U15116 ( .IN1(n13587), .IN2(n6977), .Q(n11489) );
  AND2X1 U15117 ( .IN1(n13794), .IN2(n6976), .Q(n11490) );
  AND2X1 U15118 ( .IN1(P1_N1386), .IN2(n7458), .Q(n13795) );
  AND2X1 U15119 ( .IN1(n13593), .IN2(n6872), .Q(n13796) );
  AND2X1 U15120 ( .IN1(n13607), .IN2(n6957), .Q(n13797) );
  AND2X1 U15121 ( .IN1(n13799), .IN2(n6952), .Q(n13798) );
  AND2X1 U15122 ( .IN1(n13620), .IN2(n6977), .Q(n11491) );
  AND2X1 U15123 ( .IN1(n13800), .IN2(n6982), .Q(n11492) );
  AND2X1 U15124 ( .IN1(P1_N938), .IN2(n6906), .Q(n13801) );
  AND2X1 U15125 ( .IN1(P1_N1284), .IN2(n6923), .Q(n13802) );
  AND2X1 U15126 ( .IN1(n13804), .IN2(n6874), .Q(n13803) );
  AND2X1 U15127 ( .IN1(P1_N291), .IN2(n13806), .Q(n13805) );
  AND2X1 U15128 ( .IN1(P1_N1912), .IN2(n6906), .Q(n13807) );
  AND2X1 U15129 ( .IN1(P1_N2658), .IN2(n7481), .Q(n13808) );
  AND2X1 U15130 ( .IN1(P1_N2285), .IN2(n6906), .Q(n13809) );
  AND2X1 U15131 ( .IN1(P1_N3031), .IN2(n7481), .Q(n13810) );
  AND2X1 U15132 ( .IN1(n13812), .IN2(n6860), .Q(n13811) );
  AND2X1 U15133 ( .IN1(n13814), .IN2(n6865), .Q(n13813) );
  AND2X1 U15134 ( .IN1(n13816), .IN2(n6952), .Q(n13815) );
  AND2X1 U15135 ( .IN1(n13818), .IN2(n6957), .Q(n13817) );
  AND2X1 U15136 ( .IN1(P1_N3404), .IN2(n6906), .Q(n13819) );
  AND2X1 U15137 ( .IN1(P1_N4150), .IN2(n6923), .Q(n13820) );
  AND2X1 U15138 ( .IN1(P1_N3777), .IN2(n6906), .Q(n13821) );
  AND2X1 U15139 ( .IN1(P1_N4523), .IN2(n6923), .Q(n13822) );
  AND2X1 U15140 ( .IN1(n13824), .IN2(n6860), .Q(n13823) );
  AND2X1 U15141 ( .IN1(n13826), .IN2(n6865), .Q(n13825) );
  AND2X1 U15142 ( .IN1(n13828), .IN2(n6952), .Q(n13827) );
  AND2X1 U15143 ( .IN1(n11493), .IN2(n6961), .Q(n13829) );
  AND2X1 U15144 ( .IN1(n13830), .IN2(n6984), .Q(n11495) );
  AND2X1 U15145 ( .IN1(n13831), .IN2(n6977), .Q(n11496) );
  AND2X1 U15146 ( .IN1(P1_N969), .IN2(n6906), .Q(n13832) );
  AND2X1 U15147 ( .IN1(P1_N1315), .IN2(n6923), .Q(n13833) );
  AND2X1 U15148 ( .IN1(n13835), .IN2(n6874), .Q(n13834) );
  AND2X1 U15149 ( .IN1(n11498), .IN2(P1_N291), .Q(n13836) );
  AND2X1 U15150 ( .IN1(P1_N1943), .IN2(n6906), .Q(n13837) );
  AND2X1 U15151 ( .IN1(P1_N2689), .IN2(n7481), .Q(n13838) );
  AND2X1 U15152 ( .IN1(P1_N2316), .IN2(n6906), .Q(n13839) );
  AND2X1 U15153 ( .IN1(P1_N3062), .IN2(n7481), .Q(n13840) );
  AND2X1 U15154 ( .IN1(n13842), .IN2(n6860), .Q(n13841) );
  AND2X1 U15155 ( .IN1(n13844), .IN2(n6865), .Q(n13843) );
  AND2X1 U15156 ( .IN1(n13846), .IN2(n6952), .Q(n13845) );
  AND2X1 U15157 ( .IN1(n13848), .IN2(n6959), .Q(n13847) );
  AND2X1 U15158 ( .IN1(P1_N3435), .IN2(n6906), .Q(n13849) );
  AND2X1 U15159 ( .IN1(P1_N4181), .IN2(n7481), .Q(n13850) );
  AND2X1 U15160 ( .IN1(P1_N3808), .IN2(n6906), .Q(n13851) );
  AND2X1 U15161 ( .IN1(P1_N4554), .IN2(n6923), .Q(n13852) );
  AND2X1 U15162 ( .IN1(n13854), .IN2(n6860), .Q(n13853) );
  AND2X1 U15163 ( .IN1(n13856), .IN2(n6855), .Q(n13855) );
  AND2X1 U15164 ( .IN1(n13858), .IN2(n6952), .Q(n13857) );
  AND2X1 U15165 ( .IN1(n11497), .IN2(n6959), .Q(n13859) );
  AND2X1 U15166 ( .IN1(n13860), .IN2(n6976), .Q(n11499) );
  AND2X1 U15167 ( .IN1(n13861), .IN2(n6977), .Q(n11500) );
  AND2X1 U15168 ( .IN1(P1_N968), .IN2(n6906), .Q(n13862) );
  AND2X1 U15169 ( .IN1(P1_N1314), .IN2(n6923), .Q(n13863) );
  AND2X1 U15170 ( .IN1(n13865), .IN2(n6874), .Q(n13864) );
  AND2X1 U15171 ( .IN1(n11502), .IN2(n7458), .Q(n13866) );
  AND2X1 U15172 ( .IN1(P1_N1942), .IN2(n6906), .Q(n13867) );
  AND2X1 U15173 ( .IN1(P1_N2688), .IN2(n6921), .Q(n13868) );
  AND2X1 U15174 ( .IN1(P1_N2315), .IN2(n6906), .Q(n13869) );
  AND2X1 U15175 ( .IN1(P1_N3061), .IN2(n7481), .Q(n13870) );
  AND2X1 U15176 ( .IN1(n13872), .IN2(n6860), .Q(n13871) );
  AND2X1 U15177 ( .IN1(n13874), .IN2(n6871), .Q(n13873) );
  AND2X1 U15178 ( .IN1(n13876), .IN2(n6952), .Q(n13875) );
  AND2X1 U15179 ( .IN1(n13878), .IN2(n6955), .Q(n13877) );
  AND2X1 U15180 ( .IN1(P1_N3434), .IN2(n6906), .Q(n13879) );
  AND2X1 U15181 ( .IN1(P1_N4180), .IN2(n6881), .Q(n13880) );
  AND2X1 U15182 ( .IN1(P1_N3807), .IN2(n6906), .Q(n13881) );
  AND2X1 U15183 ( .IN1(P1_N4553), .IN2(n6923), .Q(n13882) );
  AND2X1 U15184 ( .IN1(n13884), .IN2(n6860), .Q(n13883) );
  AND2X1 U15185 ( .IN1(n13886), .IN2(n7458), .Q(n13885) );
  AND2X1 U15186 ( .IN1(n13888), .IN2(n6952), .Q(n13887) );
  AND2X1 U15187 ( .IN1(n11501), .IN2(n6959), .Q(n13889) );
  AND2X1 U15188 ( .IN1(n13890), .IN2(n6982), .Q(n11503) );
  AND2X1 U15003 ( .IN1(n13680), .IN2(n6982), .Q(n11452) );
  AND2X1 U15004 ( .IN1(P1_N1367), .IN2(n6871), .Q(n13681) );
  AND2X1 U15005 ( .IN1(n12966), .IN2(n6872), .Q(n13682) );
  AND2X1 U15006 ( .IN1(n12980), .IN2(n6957), .Q(n13683) );
  AND2X1 U15007 ( .IN1(n13685), .IN2(n6958), .Q(n13684) );
  AND2X1 U15008 ( .IN1(n12993), .IN2(n6975), .Q(n11453) );
  AND2X1 U15009 ( .IN1(n13686), .IN2(n6976), .Q(n11454) );
  AND2X1 U15010 ( .IN1(P1_N1368), .IN2(n6871), .Q(n13687) );
  AND2X1 U15011 ( .IN1(n12999), .IN2(n6872), .Q(n13688) );
  AND2X1 U15012 ( .IN1(n13013), .IN2(n6957), .Q(n13689) );
  AND2X1 U15013 ( .IN1(n13691), .IN2(n6958), .Q(n13690) );
  AND2X1 U15014 ( .IN1(n13026), .IN2(n6975), .Q(n11455) );
  AND2X1 U15015 ( .IN1(n13692), .IN2(n6976), .Q(n11456) );
  AND2X1 U15016 ( .IN1(P1_N1369), .IN2(n6865), .Q(n13693) );
  AND2X1 U15017 ( .IN1(n13032), .IN2(n6866), .Q(n13694) );
  AND2X1 U15018 ( .IN1(n13046), .IN2(n6957), .Q(n13695) );
  AND2X1 U15019 ( .IN1(n13697), .IN2(n6958), .Q(n13696) );
  AND2X1 U15020 ( .IN1(n13059), .IN2(n6975), .Q(n11457) );
  AND2X1 U15021 ( .IN1(n13698), .IN2(n6976), .Q(n11458) );
  AND2X1 U15022 ( .IN1(P1_N1370), .IN2(n6865), .Q(n13699) );
  AND2X1 U15023 ( .IN1(n13065), .IN2(n6866), .Q(n13700) );
  AND2X1 U15024 ( .IN1(n13079), .IN2(n6957), .Q(n13701) );
  AND2X1 U15025 ( .IN1(n13703), .IN2(n6958), .Q(n13702) );
  AND2X1 U15026 ( .IN1(n13092), .IN2(n6975), .Q(n11459) );
  AND2X1 U15027 ( .IN1(n13704), .IN2(n6976), .Q(n11460) );
  AND2X1 U15028 ( .IN1(P1_N1371), .IN2(n6865), .Q(n13705) );
  AND2X1 U15029 ( .IN1(n13098), .IN2(n6866), .Q(n13706) );
  AND2X1 U15030 ( .IN1(n13112), .IN2(n6955), .Q(n13707) );
  AND2X1 U15031 ( .IN1(n13709), .IN2(n6956), .Q(n13708) );
  AND2X1 U15032 ( .IN1(n13125), .IN2(n6975), .Q(n11461) );
  AND2X1 U15033 ( .IN1(n13710), .IN2(n6976), .Q(n11462) );
  AND2X1 U15034 ( .IN1(P1_N1372), .IN2(n6865), .Q(n13711) );
  AND2X1 U15035 ( .IN1(n13131), .IN2(n6866), .Q(n13712) );
  AND2X1 U15036 ( .IN1(n13145), .IN2(n6955), .Q(n13713) );
  AND2X1 U15037 ( .IN1(n13715), .IN2(n6956), .Q(n13714) );
  AND2X1 U15038 ( .IN1(n13158), .IN2(n6975), .Q(n11463) );
  AND2X1 U15039 ( .IN1(n13716), .IN2(n6976), .Q(n11464) );
  AND2X1 U15040 ( .IN1(P1_N1373), .IN2(n7459), .Q(n13717) );
  AND2X1 U15041 ( .IN1(n13164), .IN2(n6854), .Q(n13718) );
  AND2X1 U15042 ( .IN1(n13178), .IN2(n6955), .Q(n13719) );
  AND2X1 U15043 ( .IN1(n13721), .IN2(n6956), .Q(n13720) );
  AND2X1 U15044 ( .IN1(n13191), .IN2(n6975), .Q(n11465) );
  AND2X1 U15045 ( .IN1(n13722), .IN2(n6976), .Q(n11466) );
  AND2X1 U15046 ( .IN1(P1_N1374), .IN2(n7459), .Q(n13723) );
  AND2X1 U15047 ( .IN1(n13197), .IN2(n6854), .Q(n13724) );
  AND2X1 U15048 ( .IN1(n13211), .IN2(n6955), .Q(n13725) );
  AND2X1 U15049 ( .IN1(n13727), .IN2(n6956), .Q(n13726) );
  AND2X1 U15050 ( .IN1(n13224), .IN2(n6975), .Q(n11467) );
  AND2X1 U15051 ( .IN1(n13728), .IN2(n6976), .Q(n11468) );
  AND2X1 U15052 ( .IN1(P1_N1375), .IN2(n7459), .Q(n13729) );
  AND2X1 U15053 ( .IN1(n13230), .IN2(n6854), .Q(n13730) );
  AND2X1 U15054 ( .IN1(n13244), .IN2(n6955), .Q(n13731) );
  AND2X1 U15055 ( .IN1(n13733), .IN2(n6956), .Q(n13732) );
  AND2X1 U15056 ( .IN1(n13257), .IN2(n6975), .Q(n11469) );
  AND2X1 U15057 ( .IN1(n13734), .IN2(n6976), .Q(n11470) );
  AND2X1 U15058 ( .IN1(P1_N1376), .IN2(n6869), .Q(n13735) );
  AND2X1 U15059 ( .IN1(n13263), .IN2(n6870), .Q(n13736) );
  AND2X1 U15060 ( .IN1(n13277), .IN2(n6949), .Q(n13737) );
  AND2X1 U15061 ( .IN1(n13739), .IN2(n6956), .Q(n13738) );
  AND2X1 U15062 ( .IN1(n13290), .IN2(n6979), .Q(n11471) );
  AND2X1 U15063 ( .IN1(n13740), .IN2(n6980), .Q(n11472) );
  AND2X1 U15064 ( .IN1(P1_N1377), .IN2(n6869), .Q(n13741) );
  AND2X1 U15065 ( .IN1(n13296), .IN2(n6870), .Q(n13742) );
  AND2X1 U15066 ( .IN1(n13310), .IN2(n6949), .Q(n13743) );
  AND2X1 U15067 ( .IN1(n13745), .IN2(n6958), .Q(n13744) );
  AND2X1 U15068 ( .IN1(n13323), .IN2(n6979), .Q(n11473) );
  AND2X1 U15069 ( .IN1(n13746), .IN2(n6980), .Q(n11474) );
  AND2X1 U15070 ( .IN1(P1_N1378), .IN2(n6857), .Q(n13747) );
  AND2X1 U15071 ( .IN1(n13329), .IN2(n6856), .Q(n13748) );
  AND2X1 U15072 ( .IN1(n13343), .IN2(n6949), .Q(n13749) );
  AND2X1 U15073 ( .IN1(n13751), .IN2(n6958), .Q(n13750) );
  AND2X1 U15074 ( .IN1(n13356), .IN2(n6979), .Q(n11475) );
  AND2X1 U15075 ( .IN1(n13752), .IN2(n6980), .Q(n11476) );
  AND2X1 U15076 ( .IN1(P1_N1379), .IN2(n6857), .Q(n13753) );
  AND2X1 U15077 ( .IN1(n13362), .IN2(n6864), .Q(n13754) );
  AND2X1 U15078 ( .IN1(n13376), .IN2(n6959), .Q(n13755) );
  AND2X1 U15079 ( .IN1(n13757), .IN2(n6958), .Q(n13756) );
  AND2X1 U15080 ( .IN1(n13389), .IN2(n6979), .Q(n11477) );
  AND2X1 U15081 ( .IN1(n13758), .IN2(n6980), .Q(n11478) );
  AND2X1 U15082 ( .IN1(P1_N1380), .IN2(P1_N291), .Q(n13759) );
  AND2X1 U15083 ( .IN1(n13395), .IN2(n6878), .Q(n13760) );
  AND2X1 U15084 ( .IN1(n13409), .IN2(n6959), .Q(n13761) );
  AND2X1 U15085 ( .IN1(n13763), .IN2(n6962), .Q(n13762) );
  AND2X1 U15086 ( .IN1(n13422), .IN2(n6977), .Q(n11479) );
  AND2X1 U15087 ( .IN1(n13764), .IN2(n6976), .Q(n11480) );
  AND2X1 U15088 ( .IN1(P1_N1381), .IN2(P1_N291), .Q(n13765) );
  AND2X1 U15089 ( .IN1(n13428), .IN2(n6878), .Q(n13766) );
  AND2X1 U15090 ( .IN1(n13442), .IN2(n6959), .Q(n13767) );
  AND2X1 U15091 ( .IN1(n13769), .IN2(n6958), .Q(n13768) );
  AND2X1 U15092 ( .IN1(n13455), .IN2(n6977), .Q(n11481) );
  AND2X1 U15093 ( .IN1(n13770), .IN2(n6980), .Q(n11482) );
  AND2X1 U15094 ( .IN1(P1_N1382), .IN2(P1_N291), .Q(n13771) );
  AND2X1 U15095 ( .IN1(n13461), .IN2(n6878), .Q(n13772) );
  AND2X1 U14910 ( .IN1(P1_N3284), .IN2(n6882), .Q(n13575) );
  AND2X1 U14911 ( .IN1(P1_N4030), .IN2(n7481), .Q(n13576) );
  AND2X1 U14912 ( .IN1(P1_N3657), .IN2(n6906), .Q(n13577) );
  AND2X1 U14913 ( .IN1(P1_N4403), .IN2(n6881), .Q(n13578) );
  AND2X1 U14914 ( .IN1(n13580), .IN2(n6860), .Q(n13579) );
  AND2X1 U14915 ( .IN1(n13582), .IN2(n6865), .Q(n13581) );
  AND2X1 U14916 ( .IN1(P1_N4653), .IN2(n6955), .Q(n13583) );
  AND2X1 U14917 ( .IN1(n13585), .IN2(n6952), .Q(n13584) );
  AND2X1 U14918 ( .IN1(n13586), .IN2(n6982), .Q(n11429) );
  AND2X1 U14919 ( .IN1(n13587), .IN2(n6977), .Q(n11430) );
  AND2X1 U14920 ( .IN1(P1_N813), .IN2(n6882), .Q(n13588) );
  AND2X1 U14921 ( .IN1(P1_N1131), .IN2(n6923), .Q(n13589) );
  AND2X1 U14922 ( .IN1(P1_N393), .IN2(n6922), .Q(n13590) );
  AND2X1 U14923 ( .IN1(P1_N1386), .IN2(n6923), .Q(n13591) );
  AND2X1 U14924 ( .IN1(n13593), .IN2(n6866), .Q(n13592) );
  AND2X1 U14925 ( .IN1(n13595), .IN2(n7458), .Q(n13594) );
  AND2X1 U14926 ( .IN1(P1_N1793), .IN2(n6886), .Q(n13596) );
  AND2X1 U14927 ( .IN1(P1_N2539), .IN2(n7481), .Q(n13597) );
  AND2X1 U14928 ( .IN1(P1_N2166), .IN2(n6886), .Q(n13598) );
  AND2X1 U14929 ( .IN1(P1_N2912), .IN2(n7481), .Q(n13599) );
  AND2X1 U14930 ( .IN1(n13601), .IN2(n6860), .Q(n13600) );
  AND2X1 U14931 ( .IN1(n13603), .IN2(n6871), .Q(n13602) );
  AND2X1 U14932 ( .IN1(n13605), .IN2(n6952), .Q(n13604) );
  AND2X1 U14933 ( .IN1(n13607), .IN2(n6959), .Q(n13606) );
  AND2X1 U14934 ( .IN1(P1_N3285), .IN2(n6906), .Q(n13608) );
  AND2X1 U14935 ( .IN1(P1_N4031), .IN2(n7481), .Q(n13609) );
  AND2X1 U14936 ( .IN1(P1_N3658), .IN2(n6906), .Q(n13610) );
  AND2X1 U14937 ( .IN1(P1_N4404), .IN2(n6921), .Q(n13611) );
  AND2X1 U14938 ( .IN1(n13613), .IN2(n6860), .Q(n13612) );
  AND2X1 U14939 ( .IN1(n13615), .IN2(n6871), .Q(n13614) );
  AND2X1 U14940 ( .IN1(P1_N4654), .IN2(n6957), .Q(n13616) );
  AND2X1 U14941 ( .IN1(n13618), .IN2(n6952), .Q(n13617) );
  AND2X1 U14942 ( .IN1(n13619), .IN2(n6976), .Q(n11431) );
  AND2X1 U14943 ( .IN1(n13620), .IN2(n6977), .Q(n11432) );
  AND2X1 U14944 ( .IN1(P1_N1357), .IN2(n7458), .Q(n13621) );
  AND2X1 U14945 ( .IN1(n12636), .IN2(n6872), .Q(n13622) );
  AND2X1 U14946 ( .IN1(n12650), .IN2(n7461), .Q(n13623) );
  AND2X1 U14947 ( .IN1(n13625), .IN2(n6954), .Q(n13624) );
  AND2X1 U14948 ( .IN1(n12663), .IN2(P1_N294), .Q(n11433) );
  AND2X1 U14949 ( .IN1(n13626), .IN2(n6984), .Q(n11434) );
  AND2X1 U14950 ( .IN1(P1_N1358), .IN2(n7458), .Q(n13627) );
  AND2X1 U14951 ( .IN1(n12669), .IN2(n6866), .Q(n13628) );
  AND2X1 U14952 ( .IN1(n12683), .IN2(n7461), .Q(n13629) );
  AND2X1 U14953 ( .IN1(n13631), .IN2(n6954), .Q(n13630) );
  AND2X1 U14954 ( .IN1(n12696), .IN2(P1_N294), .Q(n11435) );
  AND2X1 U14955 ( .IN1(n13632), .IN2(n6984), .Q(n11436) );
  AND2X1 U14956 ( .IN1(P1_N1359), .IN2(n7458), .Q(n13633) );
  AND2X1 U14957 ( .IN1(n12702), .IN2(n6872), .Q(n13634) );
  AND2X1 U14958 ( .IN1(n12716), .IN2(n7461), .Q(n13635) );
  AND2X1 U14959 ( .IN1(n13637), .IN2(n6954), .Q(n13636) );
  AND2X1 U14960 ( .IN1(n12729), .IN2(P1_N294), .Q(n11437) );
  AND2X1 U14961 ( .IN1(n13638), .IN2(n6984), .Q(n11438) );
  AND2X1 U14962 ( .IN1(P1_N1360), .IN2(n7458), .Q(n13639) );
  AND2X1 U14963 ( .IN1(n12735), .IN2(n6866), .Q(n13640) );
  AND2X1 U14964 ( .IN1(n12749), .IN2(n7461), .Q(n13641) );
  AND2X1 U14965 ( .IN1(n13643), .IN2(n6954), .Q(n13642) );
  AND2X1 U14966 ( .IN1(n12762), .IN2(P1_N294), .Q(n11439) );
  AND2X1 U14967 ( .IN1(n13644), .IN2(n6984), .Q(n11440) );
  AND2X1 U14968 ( .IN1(P1_N1361), .IN2(n7458), .Q(n13645) );
  AND2X1 U14969 ( .IN1(n12768), .IN2(n6874), .Q(n13646) );
  AND2X1 U14970 ( .IN1(n12782), .IN2(n7461), .Q(n13647) );
  AND2X1 U14971 ( .IN1(n13649), .IN2(n6954), .Q(n13648) );
  AND2X1 U14972 ( .IN1(n12795), .IN2(P1_N294), .Q(n11441) );
  AND2X1 U14973 ( .IN1(n13650), .IN2(n6984), .Q(n11442) );
  AND2X1 U14974 ( .IN1(P1_N1362), .IN2(n7458), .Q(n13651) );
  AND2X1 U14975 ( .IN1(n12801), .IN2(n6874), .Q(n13652) );
  AND2X1 U14976 ( .IN1(n12815), .IN2(n7461), .Q(n13653) );
  AND2X1 U14977 ( .IN1(n13655), .IN2(n6954), .Q(n13654) );
  AND2X1 U14978 ( .IN1(n12828), .IN2(P1_N294), .Q(n11443) );
  AND2X1 U14979 ( .IN1(n13656), .IN2(n6984), .Q(n11444) );
  AND2X1 U14980 ( .IN1(P1_N1363), .IN2(n6857), .Q(n13657) );
  AND2X1 U14981 ( .IN1(n12834), .IN2(n6864), .Q(n13658) );
  AND2X1 U14982 ( .IN1(n12848), .IN2(n6961), .Q(n13659) );
  AND2X1 U14983 ( .IN1(n13661), .IN2(n6962), .Q(n13660) );
  AND2X1 U14984 ( .IN1(n12861), .IN2(n6981), .Q(n11445) );
  AND2X1 U14985 ( .IN1(n13662), .IN2(n6982), .Q(n11446) );
  AND2X1 U14986 ( .IN1(P1_N1364), .IN2(n6857), .Q(n13663) );
  AND2X1 U14987 ( .IN1(n12867), .IN2(n6864), .Q(n13664) );
  AND2X1 U14988 ( .IN1(n12881), .IN2(n6961), .Q(n13665) );
  AND2X1 U14989 ( .IN1(n13667), .IN2(n6962), .Q(n13666) );
  AND2X1 U14990 ( .IN1(n12894), .IN2(n6981), .Q(n11447) );
  AND2X1 U14991 ( .IN1(n13668), .IN2(n6982), .Q(n11448) );
  AND2X1 U14992 ( .IN1(P1_N1365), .IN2(n6867), .Q(n13669) );
  AND2X1 U14993 ( .IN1(n12900), .IN2(n6864), .Q(n13670) );
  AND2X1 U14994 ( .IN1(n12914), .IN2(n6961), .Q(n13671) );
  AND2X1 U14995 ( .IN1(n13673), .IN2(n6962), .Q(n13672) );
  AND2X1 U14996 ( .IN1(n12927), .IN2(n6981), .Q(n11449) );
  AND2X1 U14997 ( .IN1(n13674), .IN2(n6982), .Q(n11450) );
  AND2X1 U14998 ( .IN1(P1_N1366), .IN2(n6857), .Q(n13675) );
  AND2X1 U14999 ( .IN1(n12933), .IN2(n6864), .Q(n13676) );
  AND2X1 U15000 ( .IN1(n12947), .IN2(n6957), .Q(n13677) );
  AND2X1 U15001 ( .IN1(n13679), .IN2(n6958), .Q(n13678) );
  AND2X1 U15002 ( .IN1(n12960), .IN2(n6981), .Q(n11451) );
  AND2X1 U14817 ( .IN1(P1_N4399), .IN2(n7483), .Q(n13446) );
  AND2X1 U14818 ( .IN1(n13448), .IN2(n6856), .Q(n13447) );
  AND2X1 U14819 ( .IN1(n13450), .IN2(n6855), .Q(n13449) );
  AND2X1 U14820 ( .IN1(P1_N4649), .IN2(n6959), .Q(n13451) );
  AND2X1 U14821 ( .IN1(n13453), .IN2(n6952), .Q(n13452) );
  AND2X1 U14822 ( .IN1(n13454), .IN2(n6982), .Q(n11421) );
  AND2X1 U14823 ( .IN1(n13455), .IN2(n6977), .Q(n11422) );
  AND2X1 U14824 ( .IN1(P1_N809), .IN2(n6882), .Q(n13456) );
  AND2X1 U14825 ( .IN1(P1_N1127), .IN2(n6881), .Q(n13457) );
  AND2X1 U14826 ( .IN1(P1_N389), .IN2(n6882), .Q(n13458) );
  AND2X1 U14827 ( .IN1(P1_N1382), .IN2(n6907), .Q(n13459) );
  AND2X1 U14828 ( .IN1(n13461), .IN2(n6878), .Q(n13460) );
  AND2X1 U14829 ( .IN1(n13463), .IN2(P1_N291), .Q(n13462) );
  AND2X1 U14830 ( .IN1(P1_N1789), .IN2(n6910), .Q(n13464) );
  AND2X1 U14831 ( .IN1(P1_N2535), .IN2(n7483), .Q(n13465) );
  AND2X1 U14832 ( .IN1(P1_N2162), .IN2(n6910), .Q(n13466) );
  AND2X1 U14833 ( .IN1(P1_N2908), .IN2(n7483), .Q(n13467) );
  AND2X1 U14834 ( .IN1(n13469), .IN2(n6856), .Q(n13468) );
  AND2X1 U14835 ( .IN1(n13471), .IN2(n6855), .Q(n13470) );
  AND2X1 U14836 ( .IN1(n13473), .IN2(n6952), .Q(n13472) );
  AND2X1 U14837 ( .IN1(n13475), .IN2(n6955), .Q(n13474) );
  AND2X1 U14838 ( .IN1(P1_N3281), .IN2(n6910), .Q(n13476) );
  AND2X1 U14839 ( .IN1(P1_N4027), .IN2(n7483), .Q(n13477) );
  AND2X1 U14840 ( .IN1(P1_N3654), .IN2(n6910), .Q(n13478) );
  AND2X1 U14841 ( .IN1(P1_N4400), .IN2(n7483), .Q(n13479) );
  AND2X1 U14842 ( .IN1(n13481), .IN2(n6856), .Q(n13480) );
  AND2X1 U14843 ( .IN1(n13483), .IN2(n6855), .Q(n13482) );
  AND2X1 U14844 ( .IN1(P1_N4650), .IN2(n6959), .Q(n13484) );
  AND2X1 U14845 ( .IN1(n13486), .IN2(n6952), .Q(n13485) );
  AND2X1 U14846 ( .IN1(n13487), .IN2(n6980), .Q(n11423) );
  AND2X1 U14847 ( .IN1(n13488), .IN2(n6977), .Q(n11424) );
  AND2X1 U14848 ( .IN1(P1_N810), .IN2(n6882), .Q(n13489) );
  AND2X1 U14849 ( .IN1(P1_N1128), .IN2(n6881), .Q(n13490) );
  AND2X1 U14850 ( .IN1(P1_N390), .IN2(n6882), .Q(n13491) );
  AND2X1 U14851 ( .IN1(P1_N1383), .IN2(n6881), .Q(n13492) );
  AND2X1 U14852 ( .IN1(n13494), .IN2(n6856), .Q(n13493) );
  AND2X1 U14853 ( .IN1(n13496), .IN2(n6855), .Q(n13495) );
  AND2X1 U14854 ( .IN1(P1_N1790), .IN2(n6910), .Q(n13497) );
  AND2X1 U14855 ( .IN1(P1_N2536), .IN2(n7483), .Q(n13498) );
  AND2X1 U14856 ( .IN1(P1_N2163), .IN2(n6910), .Q(n13499) );
  AND2X1 U14857 ( .IN1(P1_N2909), .IN2(n7483), .Q(n13500) );
  AND2X1 U14858 ( .IN1(n13502), .IN2(n6856), .Q(n13501) );
  AND2X1 U14859 ( .IN1(n13504), .IN2(n6855), .Q(n13503) );
  AND2X1 U14860 ( .IN1(n13506), .IN2(n6952), .Q(n13505) );
  AND2X1 U14861 ( .IN1(n13508), .IN2(n6959), .Q(n13507) );
  AND2X1 U14862 ( .IN1(P1_N3282), .IN2(n6882), .Q(n13509) );
  AND2X1 U14863 ( .IN1(P1_N4028), .IN2(n6881), .Q(n13510) );
  AND2X1 U14864 ( .IN1(P1_N3655), .IN2(n6882), .Q(n13511) );
  AND2X1 U14865 ( .IN1(P1_N4401), .IN2(n6881), .Q(n13512) );
  AND2X1 U14866 ( .IN1(n13514), .IN2(n6856), .Q(n13513) );
  AND2X1 U14867 ( .IN1(n13516), .IN2(n6855), .Q(n13515) );
  AND2X1 U14868 ( .IN1(P1_N4651), .IN2(n6959), .Q(n13517) );
  AND2X1 U14869 ( .IN1(n13519), .IN2(n6952), .Q(n13518) );
  AND2X1 U14870 ( .IN1(n13520), .IN2(n6980), .Q(n11425) );
  AND2X1 U14871 ( .IN1(n13521), .IN2(n6977), .Q(n11426) );
  AND2X1 U14872 ( .IN1(P1_N811), .IN2(n6882), .Q(n13522) );
  AND2X1 U14873 ( .IN1(P1_N1129), .IN2(n6923), .Q(n13523) );
  AND2X1 U14874 ( .IN1(P1_N391), .IN2(n6882), .Q(n13524) );
  AND2X1 U14875 ( .IN1(P1_N1384), .IN2(n6923), .Q(n13525) );
  AND2X1 U14876 ( .IN1(n13527), .IN2(n6856), .Q(n13526) );
  AND2X1 U14877 ( .IN1(n13529), .IN2(n6855), .Q(n13528) );
  AND2X1 U14878 ( .IN1(P1_N1791), .IN2(n6886), .Q(n13530) );
  AND2X1 U14879 ( .IN1(P1_N2537), .IN2(n7481), .Q(n13531) );
  AND2X1 U14880 ( .IN1(P1_N2164), .IN2(n6886), .Q(n13532) );
  AND2X1 U14881 ( .IN1(P1_N2910), .IN2(n7481), .Q(n13533) );
  AND2X1 U14882 ( .IN1(n13535), .IN2(n6856), .Q(n13534) );
  AND2X1 U14883 ( .IN1(n13537), .IN2(n6855), .Q(n13536) );
  AND2X1 U14884 ( .IN1(n13539), .IN2(n6952), .Q(n13538) );
  AND2X1 U14885 ( .IN1(n13541), .IN2(n6957), .Q(n13540) );
  AND2X1 U14886 ( .IN1(P1_N3283), .IN2(n6882), .Q(n13542) );
  AND2X1 U14887 ( .IN1(P1_N4029), .IN2(n7481), .Q(n13543) );
  AND2X1 U14888 ( .IN1(P1_N3656), .IN2(n6882), .Q(n13544) );
  AND2X1 U14889 ( .IN1(P1_N4402), .IN2(n7481), .Q(n13545) );
  AND2X1 U14890 ( .IN1(n13547), .IN2(n6856), .Q(n13546) );
  AND2X1 U14891 ( .IN1(n13549), .IN2(n6855), .Q(n13548) );
  AND2X1 U14892 ( .IN1(P1_N4652), .IN2(n6957), .Q(n13550) );
  AND2X1 U14893 ( .IN1(n13552), .IN2(n6952), .Q(n13551) );
  AND2X1 U14894 ( .IN1(n13553), .IN2(n6984), .Q(n11427) );
  AND2X1 U14895 ( .IN1(n13554), .IN2(n6977), .Q(n11428) );
  AND2X1 U14896 ( .IN1(P1_N812), .IN2(n6882), .Q(n13555) );
  AND2X1 U14897 ( .IN1(P1_N1130), .IN2(n6923), .Q(n13556) );
  AND2X1 U14898 ( .IN1(P1_N392), .IN2(n6922), .Q(n13557) );
  AND2X1 U14899 ( .IN1(P1_N1385), .IN2(n6923), .Q(n13558) );
  AND2X1 U14900 ( .IN1(n13560), .IN2(n6872), .Q(n13559) );
  AND2X1 U14901 ( .IN1(n13562), .IN2(n6855), .Q(n13561) );
  AND2X1 U14902 ( .IN1(P1_N1792), .IN2(n6886), .Q(n13563) );
  AND2X1 U14903 ( .IN1(P1_N2538), .IN2(n7481), .Q(n13564) );
  AND2X1 U14904 ( .IN1(P1_N2165), .IN2(n6882), .Q(n13565) );
  AND2X1 U14905 ( .IN1(P1_N2911), .IN2(n7481), .Q(n13566) );
  AND2X1 U14906 ( .IN1(n13568), .IN2(n6860), .Q(n13567) );
  AND2X1 U14907 ( .IN1(n13570), .IN2(n6865), .Q(n13569) );
  AND2X1 U14908 ( .IN1(n13572), .IN2(n6952), .Q(n13571) );
  AND2X1 U14909 ( .IN1(n13574), .IN2(n6955), .Q(n13573) );
  AND2X1 U14724 ( .IN1(P1_N4645), .IN2(n6949), .Q(n13319) );
  AND2X1 U14725 ( .IN1(n13321), .IN2(n6956), .Q(n13320) );
  AND2X1 U14726 ( .IN1(n13322), .IN2(n6980), .Q(n11413) );
  AND2X1 U14727 ( .IN1(n13323), .IN2(n6979), .Q(n11414) );
  AND2X1 U14728 ( .IN1(P1_N805), .IN2(n6884), .Q(n13324) );
  AND2X1 U14729 ( .IN1(P1_N1123), .IN2(n6883), .Q(n13325) );
  AND2X1 U14730 ( .IN1(P1_N385), .IN2(n6884), .Q(n13326) );
  AND2X1 U14731 ( .IN1(P1_N1378), .IN2(n6883), .Q(n13327) );
  AND2X1 U14732 ( .IN1(n13329), .IN2(n6864), .Q(n13328) );
  AND2X1 U14733 ( .IN1(n13331), .IN2(n6857), .Q(n13330) );
  AND2X1 U14734 ( .IN1(P1_N1785), .IN2(n6884), .Q(n13332) );
  AND2X1 U14735 ( .IN1(P1_N2531), .IN2(n6883), .Q(n13333) );
  AND2X1 U14736 ( .IN1(P1_N2158), .IN2(n6884), .Q(n13334) );
  AND2X1 U14737 ( .IN1(P1_N2904), .IN2(n6883), .Q(n13335) );
  AND2X1 U14738 ( .IN1(n13337), .IN2(n6864), .Q(n13336) );
  AND2X1 U14739 ( .IN1(n13339), .IN2(n6857), .Q(n13338) );
  AND2X1 U14740 ( .IN1(n13341), .IN2(n6958), .Q(n13340) );
  AND2X1 U14741 ( .IN1(n13343), .IN2(n6949), .Q(n13342) );
  AND2X1 U14742 ( .IN1(P1_N3277), .IN2(n6884), .Q(n13344) );
  AND2X1 U14743 ( .IN1(P1_N4023), .IN2(n6883), .Q(n13345) );
  AND2X1 U14744 ( .IN1(P1_N3650), .IN2(n6884), .Q(n13346) );
  AND2X1 U14745 ( .IN1(P1_N4396), .IN2(n6883), .Q(n13347) );
  AND2X1 U14746 ( .IN1(n13349), .IN2(n6856), .Q(n13348) );
  AND2X1 U14747 ( .IN1(n13351), .IN2(n6857), .Q(n13350) );
  AND2X1 U14748 ( .IN1(P1_N4646), .IN2(n6949), .Q(n13352) );
  AND2X1 U14749 ( .IN1(n13354), .IN2(n6956), .Q(n13353) );
  AND2X1 U14750 ( .IN1(n13355), .IN2(n6980), .Q(n11415) );
  AND2X1 U14751 ( .IN1(n13356), .IN2(n6979), .Q(n11416) );
  AND2X1 U14752 ( .IN1(P1_N806), .IN2(n6884), .Q(n13357) );
  AND2X1 U14753 ( .IN1(P1_N1124), .IN2(n6883), .Q(n13358) );
  AND2X1 U14754 ( .IN1(P1_N386), .IN2(n6884), .Q(n13359) );
  AND2X1 U14755 ( .IN1(P1_N1379), .IN2(n6883), .Q(n13360) );
  AND2X1 U14756 ( .IN1(n13362), .IN2(n6856), .Q(n13361) );
  AND2X1 U14757 ( .IN1(n13364), .IN2(n6857), .Q(n13363) );
  AND2X1 U14758 ( .IN1(P1_N1786), .IN2(n6884), .Q(n13365) );
  AND2X1 U14759 ( .IN1(P1_N2532), .IN2(n6883), .Q(n13366) );
  AND2X1 U14760 ( .IN1(P1_N2159), .IN2(n6888), .Q(n13367) );
  AND2X1 U14761 ( .IN1(P1_N2905), .IN2(n6907), .Q(n13368) );
  AND2X1 U14762 ( .IN1(n13370), .IN2(n6878), .Q(n13369) );
  AND2X1 U14763 ( .IN1(n13372), .IN2(P1_N291), .Q(n13371) );
  AND2X1 U14764 ( .IN1(n13374), .IN2(n6962), .Q(n13373) );
  AND2X1 U14765 ( .IN1(n13376), .IN2(n6959), .Q(n13375) );
  AND2X1 U14766 ( .IN1(P1_N3278), .IN2(n6888), .Q(n13377) );
  AND2X1 U14767 ( .IN1(P1_N4024), .IN2(n6907), .Q(n13378) );
  AND2X1 U14768 ( .IN1(P1_N3651), .IN2(n6888), .Q(n13379) );
  AND2X1 U14769 ( .IN1(P1_N4397), .IN2(n6907), .Q(n13380) );
  AND2X1 U14770 ( .IN1(n13382), .IN2(n6878), .Q(n13381) );
  AND2X1 U14771 ( .IN1(n13384), .IN2(P1_N291), .Q(n13383) );
  AND2X1 U14772 ( .IN1(P1_N4647), .IN2(n6959), .Q(n13385) );
  AND2X1 U14773 ( .IN1(n13387), .IN2(n6958), .Q(n13386) );
  AND2X1 U14774 ( .IN1(n13388), .IN2(n6980), .Q(n11417) );
  AND2X1 U14775 ( .IN1(n13389), .IN2(n6979), .Q(n11418) );
  AND2X1 U14776 ( .IN1(P1_N807), .IN2(n6888), .Q(n13390) );
  AND2X1 U14777 ( .IN1(P1_N1125), .IN2(n6907), .Q(n13391) );
  AND2X1 U14778 ( .IN1(P1_N387), .IN2(n6888), .Q(n13392) );
  AND2X1 U14779 ( .IN1(P1_N1380), .IN2(n6907), .Q(n13393) );
  AND2X1 U14780 ( .IN1(n13395), .IN2(n6878), .Q(n13394) );
  AND2X1 U14781 ( .IN1(n13397), .IN2(P1_N291), .Q(n13396) );
  AND2X1 U14782 ( .IN1(P1_N1787), .IN2(n6904), .Q(n13398) );
  AND2X1 U14783 ( .IN1(P1_N2533), .IN2(n6907), .Q(n13399) );
  AND2X1 U14784 ( .IN1(P1_N2160), .IN2(n6910), .Q(n13400) );
  AND2X1 U14785 ( .IN1(P1_N2906), .IN2(n6907), .Q(n13401) );
  AND2X1 U14786 ( .IN1(n13403), .IN2(n6878), .Q(n13402) );
  AND2X1 U14787 ( .IN1(n13405), .IN2(P1_N291), .Q(n13404) );
  AND2X1 U14788 ( .IN1(n13407), .IN2(n6962), .Q(n13406) );
  AND2X1 U14789 ( .IN1(n13409), .IN2(n6959), .Q(n13408) );
  AND2X1 U14790 ( .IN1(P1_N3279), .IN2(n6888), .Q(n13410) );
  AND2X1 U14791 ( .IN1(P1_N4025), .IN2(n6907), .Q(n13411) );
  AND2X1 U14792 ( .IN1(P1_N3652), .IN2(n6910), .Q(n13412) );
  AND2X1 U14793 ( .IN1(P1_N4398), .IN2(n7483), .Q(n13413) );
  AND2X1 U14794 ( .IN1(n13415), .IN2(n6878), .Q(n13414) );
  AND2X1 U14795 ( .IN1(n13417), .IN2(P1_N291), .Q(n13416) );
  AND2X1 U14796 ( .IN1(P1_N4648), .IN2(n6959), .Q(n13418) );
  AND2X1 U14797 ( .IN1(n13420), .IN2(n6962), .Q(n13419) );
  AND2X1 U14798 ( .IN1(n13421), .IN2(n6984), .Q(n11419) );
  AND2X1 U14799 ( .IN1(n13422), .IN2(n6977), .Q(n11420) );
  AND2X1 U14800 ( .IN1(P1_N808), .IN2(n6888), .Q(n13423) );
  AND2X1 U14801 ( .IN1(P1_N1126), .IN2(n6907), .Q(n13424) );
  AND2X1 U14802 ( .IN1(P1_N388), .IN2(n6904), .Q(n13425) );
  AND2X1 U14803 ( .IN1(P1_N1381), .IN2(n6907), .Q(n13426) );
  AND2X1 U14804 ( .IN1(n13428), .IN2(n6878), .Q(n13427) );
  AND2X1 U14805 ( .IN1(n13430), .IN2(P1_N291), .Q(n13429) );
  AND2X1 U14806 ( .IN1(P1_N1788), .IN2(n6910), .Q(n13431) );
  AND2X1 U14807 ( .IN1(P1_N2534), .IN2(n7483), .Q(n13432) );
  AND2X1 U14808 ( .IN1(P1_N2161), .IN2(n6910), .Q(n13433) );
  AND2X1 U14809 ( .IN1(P1_N2907), .IN2(n7483), .Q(n13434) );
  AND2X1 U14810 ( .IN1(n13436), .IN2(n6856), .Q(n13435) );
  AND2X1 U14811 ( .IN1(n13438), .IN2(n6855), .Q(n13437) );
  AND2X1 U14812 ( .IN1(n13440), .IN2(n6962), .Q(n13439) );
  AND2X1 U14813 ( .IN1(n13442), .IN2(n6959), .Q(n13441) );
  AND2X1 U14814 ( .IN1(P1_N3280), .IN2(n6910), .Q(n13443) );
  AND2X1 U14815 ( .IN1(P1_N4026), .IN2(n7483), .Q(n13444) );
  AND2X1 U14816 ( .IN1(P1_N3653), .IN2(n6910), .Q(n13445) );
  AND2X1 U14631 ( .IN1(n13191), .IN2(n6975), .Q(n11406) );
  AND2X1 U14632 ( .IN1(P1_N801), .IN2(n6904), .Q(n13192) );
  AND2X1 U14633 ( .IN1(P1_N1119), .IN2(n6887), .Q(n13193) );
  AND2X1 U14634 ( .IN1(P1_N381), .IN2(n6920), .Q(n13194) );
  AND2X1 U14635 ( .IN1(P1_N1374), .IN2(n6887), .Q(n13195) );
  AND2X1 U14636 ( .IN1(n13197), .IN2(n6854), .Q(n13196) );
  AND2X1 U14637 ( .IN1(n13199), .IN2(n7459), .Q(n13198) );
  AND2X1 U14638 ( .IN1(P1_N1781), .IN2(n6920), .Q(n13200) );
  AND2X1 U14639 ( .IN1(P1_N2527), .IN2(n6919), .Q(n13201) );
  AND2X1 U14640 ( .IN1(P1_N2154), .IN2(n6926), .Q(n13202) );
  AND2X1 U14641 ( .IN1(P1_N2900), .IN2(n6919), .Q(n13203) );
  AND2X1 U14642 ( .IN1(n13205), .IN2(n6854), .Q(n13204) );
  AND2X1 U14643 ( .IN1(n13207), .IN2(n7459), .Q(n13206) );
  AND2X1 U14644 ( .IN1(n13209), .IN2(n6956), .Q(n13208) );
  AND2X1 U14645 ( .IN1(n13211), .IN2(n6955), .Q(n13210) );
  AND2X1 U14646 ( .IN1(P1_N3273), .IN2(n6910), .Q(n13212) );
  AND2X1 U14647 ( .IN1(P1_N4019), .IN2(n6887), .Q(n13213) );
  AND2X1 U14648 ( .IN1(P1_N3646), .IN2(n6904), .Q(n13214) );
  AND2X1 U14649 ( .IN1(P1_N4392), .IN2(n6887), .Q(n13215) );
  AND2X1 U14650 ( .IN1(n13217), .IN2(n6854), .Q(n13216) );
  AND2X1 U14651 ( .IN1(n13219), .IN2(n7459), .Q(n13218) );
  AND2X1 U14652 ( .IN1(P1_N4642), .IN2(n6955), .Q(n13220) );
  AND2X1 U14653 ( .IN1(n13222), .IN2(n6956), .Q(n13221) );
  AND2X1 U14654 ( .IN1(n13223), .IN2(n6976), .Q(n11407) );
  AND2X1 U14655 ( .IN1(n13224), .IN2(n6975), .Q(n11408) );
  AND2X1 U14656 ( .IN1(P1_N802), .IN2(n6910), .Q(n13225) );
  AND2X1 U14657 ( .IN1(P1_N1120), .IN2(n6887), .Q(n13226) );
  AND2X1 U14658 ( .IN1(P1_N382), .IN2(n6904), .Q(n13227) );
  AND2X1 U14659 ( .IN1(P1_N1375), .IN2(n6887), .Q(n13228) );
  AND2X1 U14660 ( .IN1(n13230), .IN2(n6854), .Q(n13229) );
  AND2X1 U14661 ( .IN1(n13232), .IN2(n7459), .Q(n13231) );
  AND2X1 U14662 ( .IN1(P1_N1782), .IN2(n6904), .Q(n13233) );
  AND2X1 U14663 ( .IN1(P1_N2528), .IN2(n6887), .Q(n13234) );
  AND2X1 U14664 ( .IN1(P1_N2155), .IN2(n6904), .Q(n13235) );
  AND2X1 U14665 ( .IN1(P1_N2901), .IN2(n6887), .Q(n13236) );
  AND2X1 U14666 ( .IN1(n13238), .IN2(n6854), .Q(n13237) );
  AND2X1 U14667 ( .IN1(n13240), .IN2(n7459), .Q(n13239) );
  AND2X1 U14668 ( .IN1(n13242), .IN2(n6956), .Q(n13241) );
  AND2X1 U14669 ( .IN1(n13244), .IN2(n6955), .Q(n13243) );
  AND2X1 U14670 ( .IN1(P1_N3274), .IN2(n6904), .Q(n13245) );
  AND2X1 U14671 ( .IN1(P1_N4020), .IN2(n6887), .Q(n13246) );
  AND2X1 U14672 ( .IN1(P1_N3647), .IN2(n6910), .Q(n13247) );
  AND2X1 U14673 ( .IN1(P1_N4393), .IN2(n6887), .Q(n13248) );
  AND2X1 U14674 ( .IN1(n13250), .IN2(n6854), .Q(n13249) );
  AND2X1 U14675 ( .IN1(n13252), .IN2(n7459), .Q(n13251) );
  AND2X1 U14676 ( .IN1(P1_N4643), .IN2(n6955), .Q(n13253) );
  AND2X1 U14677 ( .IN1(n13255), .IN2(n6956), .Q(n13254) );
  AND2X1 U14678 ( .IN1(n13256), .IN2(n6976), .Q(n11409) );
  AND2X1 U14679 ( .IN1(n13257), .IN2(n6975), .Q(n11410) );
  AND2X1 U14680 ( .IN1(P1_N803), .IN2(n6894), .Q(n13258) );
  AND2X1 U14681 ( .IN1(P1_N1121), .IN2(n6893), .Q(n13259) );
  AND2X1 U14682 ( .IN1(P1_N383), .IN2(n6894), .Q(n13260) );
  AND2X1 U14683 ( .IN1(P1_N1376), .IN2(n6893), .Q(n13261) );
  AND2X1 U14684 ( .IN1(n13263), .IN2(n6870), .Q(n13262) );
  AND2X1 U14685 ( .IN1(n13265), .IN2(n6869), .Q(n13264) );
  AND2X1 U14686 ( .IN1(P1_N1783), .IN2(n6894), .Q(n13266) );
  AND2X1 U14687 ( .IN1(P1_N2529), .IN2(n6893), .Q(n13267) );
  AND2X1 U14688 ( .IN1(P1_N2156), .IN2(n6894), .Q(n13268) );
  AND2X1 U14689 ( .IN1(P1_N2902), .IN2(n6893), .Q(n13269) );
  AND2X1 U14690 ( .IN1(n13271), .IN2(n6870), .Q(n13270) );
  AND2X1 U14691 ( .IN1(n13273), .IN2(n6869), .Q(n13272) );
  AND2X1 U14692 ( .IN1(n13275), .IN2(n6956), .Q(n13274) );
  AND2X1 U14693 ( .IN1(n13277), .IN2(n6949), .Q(n13276) );
  AND2X1 U14694 ( .IN1(P1_N3275), .IN2(n6894), .Q(n13278) );
  AND2X1 U14695 ( .IN1(P1_N4021), .IN2(n6893), .Q(n13279) );
  AND2X1 U14696 ( .IN1(P1_N3648), .IN2(n6894), .Q(n13280) );
  AND2X1 U14697 ( .IN1(P1_N4394), .IN2(n6893), .Q(n13281) );
  AND2X1 U14698 ( .IN1(n13283), .IN2(n6870), .Q(n13282) );
  AND2X1 U14699 ( .IN1(n13285), .IN2(n6869), .Q(n13284) );
  AND2X1 U14700 ( .IN1(P1_N4644), .IN2(n6949), .Q(n13286) );
  AND2X1 U14701 ( .IN1(n13288), .IN2(n6958), .Q(n13287) );
  AND2X1 U14702 ( .IN1(n13289), .IN2(n6980), .Q(n11411) );
  AND2X1 U14703 ( .IN1(n13290), .IN2(n6979), .Q(n11412) );
  AND2X1 U14704 ( .IN1(P1_N804), .IN2(n6894), .Q(n13291) );
  AND2X1 U14705 ( .IN1(P1_N1122), .IN2(n6895), .Q(n13292) );
  AND2X1 U14706 ( .IN1(P1_N384), .IN2(n6896), .Q(n13293) );
  AND2X1 U14707 ( .IN1(P1_N1377), .IN2(n6895), .Q(n13294) );
  AND2X1 U14708 ( .IN1(n13296), .IN2(n6870), .Q(n13295) );
  AND2X1 U14709 ( .IN1(n13298), .IN2(n6869), .Q(n13297) );
  AND2X1 U14710 ( .IN1(P1_N1784), .IN2(n6894), .Q(n13299) );
  AND2X1 U14711 ( .IN1(P1_N2530), .IN2(n6893), .Q(n13300) );
  AND2X1 U14712 ( .IN1(P1_N2157), .IN2(n6896), .Q(n13301) );
  AND2X1 U14713 ( .IN1(P1_N2903), .IN2(n6895), .Q(n13302) );
  AND2X1 U14714 ( .IN1(n13304), .IN2(n6870), .Q(n13303) );
  AND2X1 U14715 ( .IN1(n13306), .IN2(n6869), .Q(n13305) );
  AND2X1 U14716 ( .IN1(n13308), .IN2(n6962), .Q(n13307) );
  AND2X1 U14717 ( .IN1(n13310), .IN2(n6949), .Q(n13309) );
  AND2X1 U14718 ( .IN1(P1_N3276), .IN2(n6896), .Q(n13311) );
  AND2X1 U14719 ( .IN1(P1_N4022), .IN2(n6895), .Q(n13312) );
  AND2X1 U14720 ( .IN1(P1_N3649), .IN2(n6896), .Q(n13313) );
  AND2X1 U14721 ( .IN1(P1_N4395), .IN2(n6895), .Q(n13314) );
  AND2X1 U14722 ( .IN1(n13316), .IN2(n6870), .Q(n13315) );
  AND2X1 U14723 ( .IN1(n13318), .IN2(n6857), .Q(n13317) );
  AND2X1 U14538 ( .IN1(P1_N377), .IN2(n6890), .Q(n13062) );
  AND2X1 U14539 ( .IN1(P1_N1370), .IN2(n6901), .Q(n13063) );
  AND2X1 U14540 ( .IN1(n13065), .IN2(n6866), .Q(n13064) );
  AND2X1 U14541 ( .IN1(n13067), .IN2(n6865), .Q(n13066) );
  AND2X1 U14542 ( .IN1(P1_N1777), .IN2(n6926), .Q(n13068) );
  AND2X1 U14543 ( .IN1(P1_N2523), .IN2(n6901), .Q(n13069) );
  AND2X1 U14544 ( .IN1(P1_N2150), .IN2(n6926), .Q(n13070) );
  AND2X1 U14545 ( .IN1(P1_N2896), .IN2(n6901), .Q(n13071) );
  AND2X1 U14546 ( .IN1(n13073), .IN2(n6872), .Q(n13072) );
  AND2X1 U14547 ( .IN1(n13075), .IN2(n6871), .Q(n13074) );
  AND2X1 U14548 ( .IN1(n13077), .IN2(n6958), .Q(n13076) );
  AND2X1 U14549 ( .IN1(n13079), .IN2(n6957), .Q(n13078) );
  AND2X1 U14550 ( .IN1(P1_N3269), .IN2(n6926), .Q(n13080) );
  AND2X1 U14551 ( .IN1(P1_N4015), .IN2(n6901), .Q(n13081) );
  AND2X1 U14552 ( .IN1(P1_N3642), .IN2(n6926), .Q(n13082) );
  AND2X1 U14553 ( .IN1(P1_N4388), .IN2(n6901), .Q(n13083) );
  AND2X1 U14554 ( .IN1(n13085), .IN2(n6866), .Q(n13084) );
  AND2X1 U14555 ( .IN1(n13087), .IN2(n6865), .Q(n13086) );
  AND2X1 U14556 ( .IN1(P1_N4638), .IN2(n6957), .Q(n13088) );
  AND2X1 U14557 ( .IN1(n13090), .IN2(n6958), .Q(n13089) );
  AND2X1 U14558 ( .IN1(n13091), .IN2(n6976), .Q(n11399) );
  AND2X1 U14559 ( .IN1(n13092), .IN2(n6975), .Q(n11400) );
  AND2X1 U14560 ( .IN1(P1_N798), .IN2(n6920), .Q(n13093) );
  AND2X1 U14561 ( .IN1(P1_N1116), .IN2(n6919), .Q(n13094) );
  AND2X1 U14562 ( .IN1(P1_N378), .IN2(n6890), .Q(n13095) );
  AND2X1 U14563 ( .IN1(P1_N1371), .IN2(n6901), .Q(n13096) );
  AND2X1 U14564 ( .IN1(n13098), .IN2(n6866), .Q(n13097) );
  AND2X1 U14565 ( .IN1(n13100), .IN2(n6865), .Q(n13099) );
  AND2X1 U14566 ( .IN1(P1_N1778), .IN2(n6926), .Q(n13101) );
  AND2X1 U14567 ( .IN1(P1_N2524), .IN2(n6919), .Q(n13102) );
  AND2X1 U14568 ( .IN1(P1_N2151), .IN2(n6926), .Q(n13103) );
  AND2X1 U14569 ( .IN1(P1_N2897), .IN2(n6901), .Q(n13104) );
  AND2X1 U14570 ( .IN1(n13106), .IN2(n6866), .Q(n13105) );
  AND2X1 U14571 ( .IN1(n13108), .IN2(n6865), .Q(n13107) );
  AND2X1 U14572 ( .IN1(n13110), .IN2(n6956), .Q(n13109) );
  AND2X1 U14573 ( .IN1(n13112), .IN2(n6955), .Q(n13111) );
  AND2X1 U14574 ( .IN1(P1_N3270), .IN2(n6926), .Q(n13113) );
  AND2X1 U14575 ( .IN1(P1_N4016), .IN2(n6919), .Q(n13114) );
  AND2X1 U14576 ( .IN1(P1_N3643), .IN2(n6926), .Q(n13115) );
  AND2X1 U14577 ( .IN1(P1_N4389), .IN2(n6919), .Q(n13116) );
  AND2X1 U14578 ( .IN1(n13118), .IN2(n6866), .Q(n13117) );
  AND2X1 U14579 ( .IN1(n13120), .IN2(n6865), .Q(n13119) );
  AND2X1 U14580 ( .IN1(P1_N4639), .IN2(n6955), .Q(n13121) );
  AND2X1 U14581 ( .IN1(n13123), .IN2(n6956), .Q(n13122) );
  AND2X1 U14582 ( .IN1(n13124), .IN2(n6976), .Q(n11401) );
  AND2X1 U14583 ( .IN1(n13125), .IN2(n6975), .Q(n11402) );
  AND2X1 U14584 ( .IN1(P1_N799), .IN2(n6920), .Q(n13126) );
  AND2X1 U14585 ( .IN1(P1_N1117), .IN2(n6919), .Q(n13127) );
  AND2X1 U14586 ( .IN1(P1_N379), .IN2(n6920), .Q(n13128) );
  AND2X1 U14587 ( .IN1(P1_N1372), .IN2(n6919), .Q(n13129) );
  AND2X1 U14588 ( .IN1(n13131), .IN2(n6866), .Q(n13130) );
  AND2X1 U14589 ( .IN1(n13133), .IN2(n6865), .Q(n13132) );
  AND2X1 U14590 ( .IN1(P1_N1779), .IN2(n6926), .Q(n13134) );
  AND2X1 U14591 ( .IN1(P1_N2525), .IN2(n6919), .Q(n13135) );
  AND2X1 U14592 ( .IN1(P1_N2152), .IN2(n6926), .Q(n13136) );
  AND2X1 U14593 ( .IN1(P1_N2898), .IN2(n6901), .Q(n13137) );
  AND2X1 U14594 ( .IN1(n13139), .IN2(n6866), .Q(n13138) );
  AND2X1 U14595 ( .IN1(n13141), .IN2(n6865), .Q(n13140) );
  AND2X1 U14596 ( .IN1(n13143), .IN2(n6956), .Q(n13142) );
  AND2X1 U14597 ( .IN1(n13145), .IN2(n6955), .Q(n13144) );
  AND2X1 U14598 ( .IN1(P1_N3271), .IN2(n6926), .Q(n13146) );
  AND2X1 U14599 ( .IN1(P1_N4017), .IN2(n6901), .Q(n13147) );
  AND2X1 U14600 ( .IN1(P1_N3644), .IN2(n6926), .Q(n13148) );
  AND2X1 U14601 ( .IN1(P1_N4390), .IN2(n6901), .Q(n13149) );
  AND2X1 U14602 ( .IN1(n13151), .IN2(n6866), .Q(n13150) );
  AND2X1 U14603 ( .IN1(n13153), .IN2(n6865), .Q(n13152) );
  AND2X1 U14604 ( .IN1(P1_N4640), .IN2(n6955), .Q(n13154) );
  AND2X1 U14605 ( .IN1(n13156), .IN2(n6956), .Q(n13155) );
  AND2X1 U14606 ( .IN1(n13157), .IN2(n6976), .Q(n11403) );
  AND2X1 U14607 ( .IN1(n13158), .IN2(n6975), .Q(n11404) );
  AND2X1 U14608 ( .IN1(P1_N800), .IN2(n6890), .Q(n13159) );
  AND2X1 U14609 ( .IN1(P1_N1118), .IN2(n6901), .Q(n13160) );
  AND2X1 U14610 ( .IN1(P1_N380), .IN2(n6892), .Q(n13161) );
  AND2X1 U14611 ( .IN1(P1_N1373), .IN2(n6919), .Q(n13162) );
  AND2X1 U14612 ( .IN1(n13164), .IN2(n6854), .Q(n13163) );
  AND2X1 U14613 ( .IN1(n13166), .IN2(n7459), .Q(n13165) );
  AND2X1 U14614 ( .IN1(P1_N1780), .IN2(n6890), .Q(n13167) );
  AND2X1 U14615 ( .IN1(P1_N2526), .IN2(n6919), .Q(n13168) );
  AND2X1 U14616 ( .IN1(P1_N2153), .IN2(n6926), .Q(n13169) );
  AND2X1 U14617 ( .IN1(P1_N2899), .IN2(n6919), .Q(n13170) );
  AND2X1 U14618 ( .IN1(n13172), .IN2(n6854), .Q(n13171) );
  AND2X1 U14619 ( .IN1(n13174), .IN2(n7459), .Q(n13173) );
  AND2X1 U14620 ( .IN1(n13176), .IN2(n6956), .Q(n13175) );
  AND2X1 U14621 ( .IN1(n13178), .IN2(n6955), .Q(n13177) );
  AND2X1 U14622 ( .IN1(P1_N3272), .IN2(n6892), .Q(n13179) );
  AND2X1 U14623 ( .IN1(P1_N4018), .IN2(n6901), .Q(n13180) );
  AND2X1 U14624 ( .IN1(P1_N3645), .IN2(n6926), .Q(n13181) );
  AND2X1 U14625 ( .IN1(P1_N4391), .IN2(n6901), .Q(n13182) );
  AND2X1 U14626 ( .IN1(n13184), .IN2(n6866), .Q(n13183) );
  AND2X1 U14627 ( .IN1(n13186), .IN2(n7459), .Q(n13185) );
  AND2X1 U14628 ( .IN1(P1_N4641), .IN2(n6955), .Q(n13187) );
  AND2X1 U14629 ( .IN1(n13189), .IN2(n6956), .Q(n13188) );
  AND2X1 U14630 ( .IN1(n13190), .IN2(n6976), .Q(n11405) );
  AND2X1 U14445 ( .IN1(n12935), .IN2(n6857), .Q(n12934) );
  AND2X1 U14446 ( .IN1(P1_N1773), .IN2(n6890), .Q(n12936) );
  AND2X1 U14447 ( .IN1(P1_N2519), .IN2(P1_N292), .Q(n12937) );
  AND2X1 U14448 ( .IN1(P1_N2146), .IN2(n6890), .Q(n12938) );
  AND2X1 U14449 ( .IN1(P1_N2892), .IN2(P1_N292), .Q(n12939) );
  AND2X1 U14450 ( .IN1(n12941), .IN2(n6864), .Q(n12940) );
  AND2X1 U14451 ( .IN1(n12943), .IN2(n6867), .Q(n12942) );
  AND2X1 U14452 ( .IN1(n12945), .IN2(n6958), .Q(n12944) );
  AND2X1 U14453 ( .IN1(n12947), .IN2(n6957), .Q(n12946) );
  AND2X1 U14454 ( .IN1(P1_N3265), .IN2(n6890), .Q(n12948) );
  AND2X1 U14455 ( .IN1(P1_N4011), .IN2(P1_N292), .Q(n12949) );
  AND2X1 U14456 ( .IN1(P1_N3638), .IN2(n6890), .Q(n12950) );
  AND2X1 U14457 ( .IN1(P1_N4384), .IN2(P1_N292), .Q(n12951) );
  AND2X1 U14458 ( .IN1(n12953), .IN2(n6864), .Q(n12952) );
  AND2X1 U14459 ( .IN1(n12955), .IN2(n6867), .Q(n12954) );
  AND2X1 U14460 ( .IN1(P1_N4634), .IN2(n6961), .Q(n12956) );
  AND2X1 U14461 ( .IN1(n12958), .IN2(n6958), .Q(n12957) );
  AND2X1 U14462 ( .IN1(n12959), .IN2(n6982), .Q(n11391) );
  AND2X1 U14463 ( .IN1(n12960), .IN2(n6981), .Q(n11392) );
  AND2X1 U14464 ( .IN1(P1_N794), .IN2(n6892), .Q(n12961) );
  AND2X1 U14465 ( .IN1(P1_N1112), .IN2(n6891), .Q(n12962) );
  AND2X1 U14466 ( .IN1(P1_N374), .IN2(n6892), .Q(n12963) );
  AND2X1 U14467 ( .IN1(P1_N1367), .IN2(n6891), .Q(n12964) );
  AND2X1 U14468 ( .IN1(n12966), .IN2(n6872), .Q(n12965) );
  AND2X1 U14469 ( .IN1(n12968), .IN2(n6871), .Q(n12967) );
  AND2X1 U14470 ( .IN1(P1_N1774), .IN2(n6920), .Q(n12969) );
  AND2X1 U14471 ( .IN1(P1_N2520), .IN2(n6891), .Q(n12970) );
  AND2X1 U14472 ( .IN1(P1_N2147), .IN2(n6920), .Q(n12971) );
  AND2X1 U14473 ( .IN1(P1_N2893), .IN2(n6919), .Q(n12972) );
  AND2X1 U14474 ( .IN1(n12974), .IN2(n6872), .Q(n12973) );
  AND2X1 U14475 ( .IN1(n12976), .IN2(n6871), .Q(n12975) );
  AND2X1 U14476 ( .IN1(n12978), .IN2(n6958), .Q(n12977) );
  AND2X1 U14477 ( .IN1(n12980), .IN2(n6957), .Q(n12979) );
  AND2X1 U14478 ( .IN1(P1_N3266), .IN2(n6920), .Q(n12981) );
  AND2X1 U14479 ( .IN1(P1_N4012), .IN2(n6919), .Q(n12982) );
  AND2X1 U14480 ( .IN1(P1_N3639), .IN2(n6920), .Q(n12983) );
  AND2X1 U14481 ( .IN1(P1_N4385), .IN2(n6919), .Q(n12984) );
  AND2X1 U14482 ( .IN1(n12986), .IN2(n6872), .Q(n12985) );
  AND2X1 U14483 ( .IN1(n12988), .IN2(n6871), .Q(n12987) );
  AND2X1 U14484 ( .IN1(P1_N4635), .IN2(n6957), .Q(n12989) );
  AND2X1 U14485 ( .IN1(n12991), .IN2(n6958), .Q(n12990) );
  AND2X1 U14486 ( .IN1(n12992), .IN2(n6976), .Q(n11393) );
  AND2X1 U14487 ( .IN1(n12993), .IN2(n6975), .Q(n11394) );
  AND2X1 U14488 ( .IN1(P1_N795), .IN2(n6892), .Q(n12994) );
  AND2X1 U14489 ( .IN1(P1_N1113), .IN2(n6891), .Q(n12995) );
  AND2X1 U14490 ( .IN1(P1_N375), .IN2(n6890), .Q(n12996) );
  AND2X1 U14491 ( .IN1(P1_N1368), .IN2(n6901), .Q(n12997) );
  AND2X1 U14492 ( .IN1(n12999), .IN2(n6872), .Q(n12998) );
  AND2X1 U14493 ( .IN1(n13001), .IN2(n6871), .Q(n13000) );
  AND2X1 U14494 ( .IN1(P1_N1775), .IN2(n6920), .Q(n13002) );
  AND2X1 U14495 ( .IN1(P1_N2521), .IN2(n6919), .Q(n13003) );
  AND2X1 U14496 ( .IN1(P1_N2148), .IN2(n6920), .Q(n13004) );
  AND2X1 U14497 ( .IN1(P1_N2894), .IN2(n6919), .Q(n13005) );
  AND2X1 U14498 ( .IN1(n13007), .IN2(n6872), .Q(n13006) );
  AND2X1 U14499 ( .IN1(n13009), .IN2(n6871), .Q(n13008) );
  AND2X1 U14500 ( .IN1(n13011), .IN2(n6958), .Q(n13010) );
  AND2X1 U14501 ( .IN1(n13013), .IN2(n6957), .Q(n13012) );
  AND2X1 U14502 ( .IN1(P1_N3267), .IN2(n6920), .Q(n13014) );
  AND2X1 U14503 ( .IN1(P1_N4013), .IN2(n6919), .Q(n13015) );
  AND2X1 U14504 ( .IN1(P1_N3640), .IN2(n6920), .Q(n13016) );
  AND2X1 U14505 ( .IN1(P1_N4386), .IN2(n6919), .Q(n13017) );
  AND2X1 U14506 ( .IN1(n13019), .IN2(n6872), .Q(n13018) );
  AND2X1 U14507 ( .IN1(n13021), .IN2(n6871), .Q(n13020) );
  AND2X1 U14508 ( .IN1(P1_N4636), .IN2(n6957), .Q(n13022) );
  AND2X1 U14509 ( .IN1(n13024), .IN2(n6958), .Q(n13023) );
  AND2X1 U14510 ( .IN1(n13025), .IN2(n6976), .Q(n11395) );
  AND2X1 U14511 ( .IN1(n13026), .IN2(n6975), .Q(n11396) );
  AND2X1 U14512 ( .IN1(P1_N796), .IN2(n6890), .Q(n13027) );
  AND2X1 U14513 ( .IN1(P1_N1114), .IN2(n6901), .Q(n13028) );
  AND2X1 U14514 ( .IN1(P1_N376), .IN2(n6892), .Q(n13029) );
  AND2X1 U14515 ( .IN1(P1_N1369), .IN2(n6901), .Q(n13030) );
  AND2X1 U14516 ( .IN1(n13032), .IN2(n6872), .Q(n13031) );
  AND2X1 U14517 ( .IN1(n13034), .IN2(n6865), .Q(n13033) );
  AND2X1 U14518 ( .IN1(P1_N1776), .IN2(n6920), .Q(n13035) );
  AND2X1 U14519 ( .IN1(P1_N2522), .IN2(n6919), .Q(n13036) );
  AND2X1 U14520 ( .IN1(P1_N2149), .IN2(n6920), .Q(n13037) );
  AND2X1 U14521 ( .IN1(P1_N2895), .IN2(n6919), .Q(n13038) );
  AND2X1 U14522 ( .IN1(n13040), .IN2(n6872), .Q(n13039) );
  AND2X1 U14523 ( .IN1(n13042), .IN2(n6871), .Q(n13041) );
  AND2X1 U14524 ( .IN1(n13044), .IN2(n6958), .Q(n13043) );
  AND2X1 U14525 ( .IN1(n13046), .IN2(n6957), .Q(n13045) );
  AND2X1 U14526 ( .IN1(P1_N3268), .IN2(n6920), .Q(n13047) );
  AND2X1 U14527 ( .IN1(P1_N4014), .IN2(n6919), .Q(n13048) );
  AND2X1 U14528 ( .IN1(P1_N3641), .IN2(n6920), .Q(n13049) );
  AND2X1 U14529 ( .IN1(P1_N4387), .IN2(n6919), .Q(n13050) );
  AND2X1 U14530 ( .IN1(n13052), .IN2(n6872), .Q(n13051) );
  AND2X1 U14531 ( .IN1(n13054), .IN2(n6871), .Q(n13053) );
  AND2X1 U14532 ( .IN1(P1_N4637), .IN2(n6957), .Q(n13055) );
  AND2X1 U14533 ( .IN1(n13057), .IN2(n6958), .Q(n13056) );
  AND2X1 U14534 ( .IN1(n13058), .IN2(n6976), .Q(n11397) );
  AND2X1 U14535 ( .IN1(n13059), .IN2(n6975), .Q(n11398) );
  AND2X1 U14536 ( .IN1(P1_N797), .IN2(n6920), .Q(n13060) );
  AND2X1 U14537 ( .IN1(P1_N1115), .IN2(n6901), .Q(n13061) );
  AND2X1 U14352 ( .IN1(P1_N2142), .IN2(n6888), .Q(n12806) );
  AND2X1 U14353 ( .IN1(P1_N2888), .IN2(n6887), .Q(n12807) );
  AND2X1 U14354 ( .IN1(n12809), .IN2(n6874), .Q(n12808) );
  AND2X1 U14355 ( .IN1(n12811), .IN2(n7458), .Q(n12810) );
  AND2X1 U14356 ( .IN1(n12813), .IN2(n6954), .Q(n12812) );
  AND2X1 U14357 ( .IN1(n12815), .IN2(n7461), .Q(n12814) );
  AND2X1 U14358 ( .IN1(P1_N3261), .IN2(n6888), .Q(n12816) );
  AND2X1 U14359 ( .IN1(P1_N4007), .IN2(n6887), .Q(n12817) );
  AND2X1 U14360 ( .IN1(P1_N3634), .IN2(n6888), .Q(n12818) );
  AND2X1 U14361 ( .IN1(P1_N4380), .IN2(n6887), .Q(n12819) );
  AND2X1 U14362 ( .IN1(n12821), .IN2(n6874), .Q(n12820) );
  AND2X1 U14363 ( .IN1(n12823), .IN2(n7458), .Q(n12822) );
  AND2X1 U14364 ( .IN1(P1_N4630), .IN2(n7461), .Q(n12824) );
  AND2X1 U14365 ( .IN1(n12826), .IN2(n6954), .Q(n12825) );
  AND2X1 U14366 ( .IN1(n12827), .IN2(n6984), .Q(n11383) );
  AND2X1 U14367 ( .IN1(n12828), .IN2(P1_N294), .Q(n11384) );
  AND2X1 U14368 ( .IN1(P1_N790), .IN2(n6904), .Q(n12829) );
  AND2X1 U14369 ( .IN1(P1_N1108), .IN2(n7483), .Q(n12830) );
  AND2X1 U14370 ( .IN1(P1_N370), .IN2(n6904), .Q(n12831) );
  AND2X1 U14371 ( .IN1(P1_N1363), .IN2(n7483), .Q(n12832) );
  AND2X1 U14372 ( .IN1(n12834), .IN2(n6864), .Q(n12833) );
  AND2X1 U14373 ( .IN1(n12836), .IN2(n6867), .Q(n12835) );
  AND2X1 U14374 ( .IN1(P1_N1770), .IN2(n6904), .Q(n12837) );
  AND2X1 U14375 ( .IN1(P1_N2516), .IN2(n7483), .Q(n12838) );
  AND2X1 U14376 ( .IN1(P1_N2143), .IN2(n6904), .Q(n12839) );
  AND2X1 U14377 ( .IN1(P1_N2889), .IN2(n7483), .Q(n12840) );
  AND2X1 U14378 ( .IN1(n12842), .IN2(n6864), .Q(n12841) );
  AND2X1 U14379 ( .IN1(n12844), .IN2(n6867), .Q(n12843) );
  AND2X1 U14380 ( .IN1(n12846), .IN2(n6962), .Q(n12845) );
  AND2X1 U14381 ( .IN1(n12848), .IN2(n6961), .Q(n12847) );
  AND2X1 U14382 ( .IN1(P1_N3262), .IN2(n6904), .Q(n12849) );
  AND2X1 U14383 ( .IN1(P1_N4008), .IN2(n7483), .Q(n12850) );
  AND2X1 U14384 ( .IN1(P1_N3635), .IN2(n6904), .Q(n12851) );
  AND2X1 U14385 ( .IN1(P1_N4381), .IN2(n7483), .Q(n12852) );
  AND2X1 U14386 ( .IN1(n12854), .IN2(n6864), .Q(n12853) );
  AND2X1 U14387 ( .IN1(n12856), .IN2(n6867), .Q(n12855) );
  AND2X1 U14388 ( .IN1(P1_N4631), .IN2(n6961), .Q(n12857) );
  AND2X1 U14389 ( .IN1(n12859), .IN2(n6962), .Q(n12858) );
  AND2X1 U14390 ( .IN1(n12860), .IN2(n6982), .Q(n11385) );
  AND2X1 U14391 ( .IN1(n12861), .IN2(n6981), .Q(n11386) );
  AND2X1 U14392 ( .IN1(P1_N791), .IN2(n6890), .Q(n12862) );
  AND2X1 U14393 ( .IN1(P1_N1109), .IN2(P1_N292), .Q(n12863) );
  AND2X1 U14394 ( .IN1(P1_N371), .IN2(n6904), .Q(n12864) );
  AND2X1 U14395 ( .IN1(P1_N1364), .IN2(n7483), .Q(n12865) );
  AND2X1 U14396 ( .IN1(n12867), .IN2(n6864), .Q(n12866) );
  AND2X1 U14397 ( .IN1(n12869), .IN2(n6867), .Q(n12868) );
  AND2X1 U14398 ( .IN1(P1_N1771), .IN2(n6904), .Q(n12870) );
  AND2X1 U14399 ( .IN1(P1_N2517), .IN2(n7483), .Q(n12871) );
  AND2X1 U14400 ( .IN1(P1_N2144), .IN2(n6904), .Q(n12872) );
  AND2X1 U14401 ( .IN1(P1_N2890), .IN2(n7483), .Q(n12873) );
  AND2X1 U14402 ( .IN1(n12875), .IN2(n6864), .Q(n12874) );
  AND2X1 U14403 ( .IN1(n12877), .IN2(n6867), .Q(n12876) );
  AND2X1 U14404 ( .IN1(n12879), .IN2(n6962), .Q(n12878) );
  AND2X1 U14405 ( .IN1(n12881), .IN2(n6961), .Q(n12880) );
  AND2X1 U14406 ( .IN1(P1_N3263), .IN2(n6904), .Q(n12882) );
  AND2X1 U14407 ( .IN1(P1_N4009), .IN2(n7483), .Q(n12883) );
  AND2X1 U14408 ( .IN1(P1_N3636), .IN2(n6890), .Q(n12884) );
  AND2X1 U14409 ( .IN1(P1_N4382), .IN2(P1_N292), .Q(n12885) );
  AND2X1 U14410 ( .IN1(n12887), .IN2(n6864), .Q(n12886) );
  AND2X1 U14411 ( .IN1(n12889), .IN2(n6867), .Q(n12888) );
  AND2X1 U14412 ( .IN1(P1_N4632), .IN2(n6961), .Q(n12890) );
  AND2X1 U14413 ( .IN1(n12892), .IN2(n6962), .Q(n12891) );
  AND2X1 U14414 ( .IN1(n12893), .IN2(n6982), .Q(n11387) );
  AND2X1 U14415 ( .IN1(n12894), .IN2(n6981), .Q(n11388) );
  AND2X1 U14416 ( .IN1(P1_N792), .IN2(n6890), .Q(n12895) );
  AND2X1 U14417 ( .IN1(P1_N1110), .IN2(P1_N292), .Q(n12896) );
  AND2X1 U14418 ( .IN1(P1_N372), .IN2(n6890), .Q(n12897) );
  AND2X1 U14419 ( .IN1(P1_N1365), .IN2(P1_N292), .Q(n12898) );
  AND2X1 U14420 ( .IN1(n12900), .IN2(n6864), .Q(n12899) );
  AND2X1 U14421 ( .IN1(n12902), .IN2(n6857), .Q(n12901) );
  AND2X1 U14422 ( .IN1(P1_N1772), .IN2(n6890), .Q(n12903) );
  AND2X1 U14423 ( .IN1(P1_N2518), .IN2(P1_N292), .Q(n12904) );
  AND2X1 U14424 ( .IN1(P1_N2145), .IN2(n6890), .Q(n12905) );
  AND2X1 U14425 ( .IN1(P1_N2891), .IN2(P1_N292), .Q(n12906) );
  AND2X1 U14426 ( .IN1(n12908), .IN2(n6864), .Q(n12907) );
  AND2X1 U14427 ( .IN1(n12910), .IN2(n6867), .Q(n12909) );
  AND2X1 U14428 ( .IN1(n12912), .IN2(n6962), .Q(n12911) );
  AND2X1 U14429 ( .IN1(n12914), .IN2(n6961), .Q(n12913) );
  AND2X1 U14430 ( .IN1(P1_N3264), .IN2(n6890), .Q(n12915) );
  AND2X1 U14431 ( .IN1(P1_N4010), .IN2(P1_N292), .Q(n12916) );
  AND2X1 U14432 ( .IN1(P1_N3637), .IN2(n6890), .Q(n12917) );
  AND2X1 U14433 ( .IN1(P1_N4383), .IN2(P1_N292), .Q(n12918) );
  AND2X1 U14434 ( .IN1(n12920), .IN2(n6864), .Q(n12919) );
  AND2X1 U14435 ( .IN1(n12922), .IN2(n6857), .Q(n12921) );
  AND2X1 U14436 ( .IN1(P1_N4633), .IN2(n6961), .Q(n12923) );
  AND2X1 U14437 ( .IN1(n12925), .IN2(n6962), .Q(n12924) );
  AND2X1 U14438 ( .IN1(n12926), .IN2(n6982), .Q(n11389) );
  AND2X1 U14439 ( .IN1(n12927), .IN2(n6981), .Q(n11390) );
  AND2X1 U14440 ( .IN1(P1_N793), .IN2(n6890), .Q(n12928) );
  AND2X1 U14441 ( .IN1(P1_N1111), .IN2(P1_N292), .Q(n12929) );
  AND2X1 U14442 ( .IN1(P1_N373), .IN2(n6890), .Q(n12930) );
  AND2X1 U14443 ( .IN1(P1_N1366), .IN2(P1_N292), .Q(n12931) );
  AND2X1 U14444 ( .IN1(n12933), .IN2(n6864), .Q(n12932) );
  AND2X1 U14259 ( .IN1(n12679), .IN2(n6865), .Q(n12678) );
  AND2X1 U14260 ( .IN1(n12681), .IN2(n6954), .Q(n12680) );
  AND2X1 U14261 ( .IN1(n12683), .IN2(n7461), .Q(n12682) );
  AND2X1 U14262 ( .IN1(P1_N3257), .IN2(n6922), .Q(n12684) );
  AND2X1 U14263 ( .IN1(P1_N4003), .IN2(n6921), .Q(n12685) );
  AND2X1 U14264 ( .IN1(P1_N3630), .IN2(n6922), .Q(n12686) );
  AND2X1 U14265 ( .IN1(P1_N4376), .IN2(n6921), .Q(n12687) );
  AND2X1 U14266 ( .IN1(n12689), .IN2(n6860), .Q(n12688) );
  AND2X1 U14267 ( .IN1(n12691), .IN2(n6865), .Q(n12690) );
  AND2X1 U14268 ( .IN1(P1_N4626), .IN2(n7461), .Q(n12692) );
  AND2X1 U14269 ( .IN1(n12694), .IN2(n6954), .Q(n12693) );
  AND2X1 U14270 ( .IN1(n12695), .IN2(n6984), .Q(n11375) );
  AND2X1 U14271 ( .IN1(n12696), .IN2(P1_N294), .Q(n11376) );
  AND2X1 U14272 ( .IN1(P1_N786), .IN2(n6886), .Q(n12697) );
  AND2X1 U14273 ( .IN1(P1_N1104), .IN2(n6921), .Q(n12698) );
  AND2X1 U14274 ( .IN1(n6623), .IN2(n6886), .Q(n12699) );
  AND2X1 U14275 ( .IN1(P1_N1359), .IN2(n6921), .Q(n12700) );
  AND2X1 U14276 ( .IN1(n12702), .IN2(n6872), .Q(n12701) );
  AND2X1 U14277 ( .IN1(n12704), .IN2(n7458), .Q(n12703) );
  AND2X1 U14278 ( .IN1(P1_N1766), .IN2(n6922), .Q(n12705) );
  AND2X1 U14279 ( .IN1(P1_N2512), .IN2(n6921), .Q(n12706) );
  AND2X1 U14280 ( .IN1(P1_N2139), .IN2(n6922), .Q(n12707) );
  AND2X1 U14281 ( .IN1(P1_N2885), .IN2(n6921), .Q(n12708) );
  AND2X1 U14282 ( .IN1(n12710), .IN2(n6860), .Q(n12709) );
  AND2X1 U14283 ( .IN1(n12712), .IN2(n6865), .Q(n12711) );
  AND2X1 U14284 ( .IN1(n12714), .IN2(n6954), .Q(n12713) );
  AND2X1 U14285 ( .IN1(n12716), .IN2(n7461), .Q(n12715) );
  AND2X1 U14286 ( .IN1(P1_N3258), .IN2(n6922), .Q(n12717) );
  AND2X1 U14287 ( .IN1(P1_N4004), .IN2(n6921), .Q(n12718) );
  AND2X1 U14288 ( .IN1(P1_N3631), .IN2(n6922), .Q(n12719) );
  AND2X1 U14289 ( .IN1(P1_N4377), .IN2(n6921), .Q(n12720) );
  AND2X1 U14290 ( .IN1(n12722), .IN2(n6860), .Q(n12721) );
  AND2X1 U14291 ( .IN1(n12724), .IN2(n6865), .Q(n12723) );
  AND2X1 U14292 ( .IN1(P1_N4627), .IN2(n7461), .Q(n12725) );
  AND2X1 U14293 ( .IN1(n12727), .IN2(n6954), .Q(n12726) );
  AND2X1 U14294 ( .IN1(n12728), .IN2(n6984), .Q(n11377) );
  AND2X1 U14295 ( .IN1(n12729), .IN2(P1_N294), .Q(n11378) );
  AND2X1 U14296 ( .IN1(P1_N787), .IN2(n6886), .Q(n12730) );
  AND2X1 U14297 ( .IN1(P1_N1105), .IN2(n6921), .Q(n12731) );
  AND2X1 U14298 ( .IN1(n18451), .IN2(n6886), .Q(n12732) );
  AND2X1 U14299 ( .IN1(P1_N1360), .IN2(n6921), .Q(n12733) );
  AND2X1 U14300 ( .IN1(n12735), .IN2(n6872), .Q(n12734) );
  AND2X1 U14301 ( .IN1(n12737), .IN2(n7458), .Q(n12736) );
  AND2X1 U14302 ( .IN1(P1_N1767), .IN2(n6922), .Q(n12738) );
  AND2X1 U14303 ( .IN1(P1_N2513), .IN2(n6921), .Q(n12739) );
  AND2X1 U14304 ( .IN1(P1_N2140), .IN2(n6922), .Q(n12740) );
  AND2X1 U14305 ( .IN1(P1_N2886), .IN2(n6921), .Q(n12741) );
  AND2X1 U14306 ( .IN1(n12743), .IN2(n6860), .Q(n12742) );
  AND2X1 U14307 ( .IN1(n12745), .IN2(n6865), .Q(n12744) );
  AND2X1 U14308 ( .IN1(n12747), .IN2(n6954), .Q(n12746) );
  AND2X1 U14309 ( .IN1(n12749), .IN2(n7461), .Q(n12748) );
  AND2X1 U14310 ( .IN1(P1_N3259), .IN2(n6922), .Q(n12750) );
  AND2X1 U14311 ( .IN1(P1_N4005), .IN2(n6921), .Q(n12751) );
  AND2X1 U14312 ( .IN1(P1_N3632), .IN2(n6922), .Q(n12752) );
  AND2X1 U14313 ( .IN1(P1_N4378), .IN2(n6921), .Q(n12753) );
  AND2X1 U14314 ( .IN1(n12755), .IN2(n6860), .Q(n12754) );
  AND2X1 U14315 ( .IN1(n12757), .IN2(n6865), .Q(n12756) );
  AND2X1 U14316 ( .IN1(P1_N4628), .IN2(n7461), .Q(n12758) );
  AND2X1 U14317 ( .IN1(n12760), .IN2(n6954), .Q(n12759) );
  AND2X1 U14318 ( .IN1(n12761), .IN2(n6984), .Q(n11379) );
  AND2X1 U14319 ( .IN1(n12762), .IN2(P1_N294), .Q(n11380) );
  AND2X1 U14320 ( .IN1(P1_N788), .IN2(n6888), .Q(n12763) );
  AND2X1 U14321 ( .IN1(P1_N1106), .IN2(n6887), .Q(n12764) );
  AND2X1 U14322 ( .IN1(P1_N368), .IN2(n6886), .Q(n12765) );
  AND2X1 U14323 ( .IN1(P1_N1361), .IN2(n6887), .Q(n12766) );
  AND2X1 U14324 ( .IN1(n12768), .IN2(n6874), .Q(n12767) );
  AND2X1 U14325 ( .IN1(n12770), .IN2(n7458), .Q(n12769) );
  AND2X1 U14326 ( .IN1(P1_N1768), .IN2(n6888), .Q(n12771) );
  AND2X1 U14327 ( .IN1(P1_N2514), .IN2(n6887), .Q(n12772) );
  AND2X1 U14328 ( .IN1(P1_N2141), .IN2(n6888), .Q(n12773) );
  AND2X1 U14329 ( .IN1(P1_N2887), .IN2(n6887), .Q(n12774) );
  AND2X1 U14330 ( .IN1(n12776), .IN2(n6874), .Q(n12775) );
  AND2X1 U14331 ( .IN1(n12778), .IN2(n7458), .Q(n12777) );
  AND2X1 U14332 ( .IN1(n12780), .IN2(n6954), .Q(n12779) );
  AND2X1 U14333 ( .IN1(n12782), .IN2(n7461), .Q(n12781) );
  AND2X1 U14334 ( .IN1(P1_N3260), .IN2(n6888), .Q(n12783) );
  AND2X1 U14335 ( .IN1(P1_N4006), .IN2(n6887), .Q(n12784) );
  AND2X1 U14336 ( .IN1(P1_N3633), .IN2(n6888), .Q(n12785) );
  AND2X1 U14337 ( .IN1(P1_N4379), .IN2(n6887), .Q(n12786) );
  AND2X1 U14338 ( .IN1(n12788), .IN2(n6874), .Q(n12787) );
  AND2X1 U14339 ( .IN1(n12790), .IN2(n7458), .Q(n12789) );
  AND2X1 U14340 ( .IN1(P1_N4629), .IN2(n7461), .Q(n12791) );
  AND2X1 U14341 ( .IN1(n12793), .IN2(n6954), .Q(n12792) );
  AND2X1 U14342 ( .IN1(n12794), .IN2(n6984), .Q(n11381) );
  AND2X1 U14343 ( .IN1(n12795), .IN2(P1_N294), .Q(n11382) );
  AND2X1 U14344 ( .IN1(P1_N789), .IN2(n6888), .Q(n12796) );
  AND2X1 U14345 ( .IN1(P1_N1107), .IN2(n6887), .Q(n12797) );
  AND2X1 U14346 ( .IN1(P1_N369), .IN2(n6888), .Q(n12798) );
  AND2X1 U14347 ( .IN1(P1_N1362), .IN2(n6887), .Q(n12799) );
  AND2X1 U14348 ( .IN1(n12801), .IN2(n6874), .Q(n12800) );
  AND2X1 U14349 ( .IN1(n12803), .IN2(n7458), .Q(n12802) );
  AND2X1 U14350 ( .IN1(P1_N1769), .IN2(n6888), .Q(n12804) );
  AND2X1 U14351 ( .IN1(P1_N2515), .IN2(n6887), .Q(n12805) );
  AND2X1 U14166 ( .IN1(P1_N390), .IN2(n11309), .Q(n12551) );
  AND2X1 U14167 ( .IN1(P1_N4813), .IN2(n6992), .Q(n12552) );
  AND2X1 U14168 ( .IN1(n12554), .IN2(n6952), .Q(n12553) );
  AND2X1 U14169 ( .IN1(n12556), .IN2(n6955), .Q(n12555) );
  AND2X1 U14170 ( .IN1(n12557), .IN2(n6980), .Q(n11367) );
  AND2X1 U14171 ( .IN1(n12558), .IN2(n6977), .Q(n11368) );
  AND2X1 U14172 ( .IN1(P1_N966), .IN2(n6922), .Q(n12559) );
  AND2X1 U14173 ( .IN1(P1_N1312), .IN2(n6923), .Q(n12560) );
  AND2X1 U14174 ( .IN1(P1_N1038), .IN2(n6886), .Q(n12561) );
  AND2X1 U14175 ( .IN1(P1_N1567), .IN2(n6923), .Q(n12562) );
  AND2X1 U14176 ( .IN1(n12564), .IN2(n6856), .Q(n12563) );
  AND2X1 U14177 ( .IN1(n12566), .IN2(n6855), .Q(n12565) );
  AND2X1 U14178 ( .IN1(P1_N1940), .IN2(n6882), .Q(n12567) );
  AND2X1 U14179 ( .IN1(P1_N2686), .IN2(n6881), .Q(n12568) );
  AND2X1 U14180 ( .IN1(P1_N2313), .IN2(n6882), .Q(n12569) );
  AND2X1 U14181 ( .IN1(P1_N3059), .IN2(n6881), .Q(n12570) );
  AND2X1 U14182 ( .IN1(n12572), .IN2(n6856), .Q(n12571) );
  AND2X1 U14183 ( .IN1(n12574), .IN2(n6855), .Q(n12573) );
  AND2X1 U14184 ( .IN1(n12576), .IN2(n6952), .Q(n12575) );
  AND2X1 U14185 ( .IN1(n12578), .IN2(n6957), .Q(n12577) );
  AND2X1 U14186 ( .IN1(P1_N3432), .IN2(n6882), .Q(n12579) );
  AND2X1 U14187 ( .IN1(P1_N4178), .IN2(n6923), .Q(n12580) );
  AND2X1 U14188 ( .IN1(P1_N3805), .IN2(n6882), .Q(n12581) );
  AND2X1 U14189 ( .IN1(P1_N4551), .IN2(n6881), .Q(n12582) );
  AND2X1 U14190 ( .IN1(n12584), .IN2(n6856), .Q(n12583) );
  AND2X1 U14191 ( .IN1(n12586), .IN2(n6855), .Q(n12585) );
  AND2X1 U14192 ( .IN1(P1_N391), .IN2(n11309), .Q(n12587) );
  AND2X1 U14193 ( .IN1(P1_N4814), .IN2(n6992), .Q(n12588) );
  AND2X1 U14194 ( .IN1(n12590), .IN2(n6952), .Q(n12589) );
  AND2X1 U14195 ( .IN1(n12592), .IN2(n6959), .Q(n12591) );
  AND2X1 U14196 ( .IN1(n12593), .IN2(n6980), .Q(n11369) );
  AND2X1 U14197 ( .IN1(n12594), .IN2(n6977), .Q(n11370) );
  AND2X1 U14198 ( .IN1(P1_N967), .IN2(n6922), .Q(n12595) );
  AND2X1 U14199 ( .IN1(P1_N1313), .IN2(n6923), .Q(n12596) );
  AND2X1 U14200 ( .IN1(P1_N1039), .IN2(n6922), .Q(n12597) );
  AND2X1 U14201 ( .IN1(P1_N1568), .IN2(n6923), .Q(n12598) );
  AND2X1 U14202 ( .IN1(n12600), .IN2(n6856), .Q(n12599) );
  AND2X1 U14203 ( .IN1(n12602), .IN2(n6855), .Q(n12601) );
  AND2X1 U14204 ( .IN1(P1_N1941), .IN2(n6882), .Q(n12603) );
  AND2X1 U14205 ( .IN1(P1_N2687), .IN2(n6923), .Q(n12604) );
  AND2X1 U14206 ( .IN1(P1_N2314), .IN2(n6922), .Q(n12605) );
  AND2X1 U14207 ( .IN1(P1_N3060), .IN2(n6923), .Q(n12606) );
  AND2X1 U14208 ( .IN1(n12608), .IN2(n6856), .Q(n12607) );
  AND2X1 U14209 ( .IN1(n12610), .IN2(n6855), .Q(n12609) );
  AND2X1 U14210 ( .IN1(n12612), .IN2(n6952), .Q(n12611) );
  AND2X1 U14211 ( .IN1(n12614), .IN2(n6959), .Q(n12613) );
  AND2X1 U14212 ( .IN1(P1_N3433), .IN2(n6882), .Q(n12615) );
  AND2X1 U14213 ( .IN1(P1_N4179), .IN2(n6923), .Q(n12616) );
  AND2X1 U14214 ( .IN1(P1_N3806), .IN2(n6922), .Q(n12617) );
  AND2X1 U14215 ( .IN1(P1_N4552), .IN2(n6923), .Q(n12618) );
  AND2X1 U14216 ( .IN1(n12620), .IN2(n6856), .Q(n12619) );
  AND2X1 U14217 ( .IN1(n12622), .IN2(n6855), .Q(n12621) );
  AND2X1 U14218 ( .IN1(P1_N392), .IN2(n11309), .Q(n12623) );
  AND2X1 U14219 ( .IN1(P1_N4815), .IN2(n6992), .Q(n12624) );
  AND2X1 U14220 ( .IN1(n12626), .IN2(n6952), .Q(n12625) );
  AND2X1 U14221 ( .IN1(n12628), .IN2(n6959), .Q(n12627) );
  AND2X1 U14222 ( .IN1(n12629), .IN2(n6976), .Q(n11371) );
  AND2X1 U14223 ( .IN1(n12630), .IN2(n6977), .Q(n11372) );
  AND2X1 U14224 ( .IN1(P1_N630), .IN2(n6886), .Q(n12631) );
  AND2X1 U14225 ( .IN1(P1_N1102), .IN2(n6921), .Q(n12632) );
  AND2X1 U14226 ( .IN1(n6621), .IN2(n6886), .Q(n12633) );
  AND2X1 U14227 ( .IN1(P1_N1357), .IN2(n6881), .Q(n12634) );
  AND2X1 U14228 ( .IN1(n12636), .IN2(n6866), .Q(n12635) );
  AND2X1 U14229 ( .IN1(n12638), .IN2(n7458), .Q(n12637) );
  AND2X1 U14230 ( .IN1(P1_N1764), .IN2(n6906), .Q(n12639) );
  AND2X1 U14231 ( .IN1(P1_N2510), .IN2(n6921), .Q(n12640) );
  AND2X1 U14232 ( .IN1(P1_N2137), .IN2(n6906), .Q(n12641) );
  AND2X1 U14233 ( .IN1(P1_N2883), .IN2(n7481), .Q(n12642) );
  AND2X1 U14234 ( .IN1(n12644), .IN2(n6860), .Q(n12643) );
  AND2X1 U14235 ( .IN1(n12646), .IN2(n6865), .Q(n12645) );
  AND2X1 U14236 ( .IN1(n12648), .IN2(n6954), .Q(n12647) );
  AND2X1 U14237 ( .IN1(n12650), .IN2(n7461), .Q(n12649) );
  AND2X1 U14238 ( .IN1(P1_N3256), .IN2(n6922), .Q(n12651) );
  AND2X1 U14239 ( .IN1(P1_N4002), .IN2(n6921), .Q(n12652) );
  AND2X1 U14240 ( .IN1(P1_N3629), .IN2(n6922), .Q(n12653) );
  AND2X1 U14241 ( .IN1(P1_N4375), .IN2(n6921), .Q(n12654) );
  AND2X1 U14242 ( .IN1(n12656), .IN2(n6860), .Q(n12655) );
  AND2X1 U14243 ( .IN1(n12658), .IN2(n6865), .Q(n12657) );
  AND2X1 U14244 ( .IN1(P1_N4625), .IN2(n7461), .Q(n12659) );
  AND2X1 U14245 ( .IN1(n12661), .IN2(n6954), .Q(n12660) );
  AND2X1 U14246 ( .IN1(n12662), .IN2(n6984), .Q(n11373) );
  AND2X1 U14247 ( .IN1(n12663), .IN2(P1_N294), .Q(n11374) );
  AND2X1 U14248 ( .IN1(P1_N785), .IN2(n6886), .Q(n12664) );
  AND2X1 U14249 ( .IN1(P1_N1103), .IN2(n6921), .Q(n12665) );
  AND2X1 U14250 ( .IN1(n6622), .IN2(n6886), .Q(n12666) );
  AND2X1 U14251 ( .IN1(P1_N1358), .IN2(n6881), .Q(n12667) );
  AND2X1 U14252 ( .IN1(n12669), .IN2(n6866), .Q(n12668) );
  AND2X1 U14253 ( .IN1(n12671), .IN2(n7458), .Q(n12670) );
  AND2X1 U14254 ( .IN1(P1_N1765), .IN2(n6922), .Q(n12672) );
  AND2X1 U14255 ( .IN1(P1_N2511), .IN2(n7481), .Q(n12673) );
  AND2X1 U14256 ( .IN1(P1_N2138), .IN2(n6886), .Q(n12674) );
  AND2X1 U14257 ( .IN1(P1_N2884), .IN2(n7481), .Q(n12675) );
  AND2X1 U14258 ( .IN1(n12677), .IN2(n6860), .Q(n12676) );
  AND2X1 U14073 ( .IN1(n12422), .IN2(P1_N291), .Q(n12421) );
  AND2X1 U14074 ( .IN1(P1_N1936), .IN2(n6888), .Q(n12423) );
  AND2X1 U14075 ( .IN1(P1_N2682), .IN2(n6907), .Q(n12424) );
  AND2X1 U14076 ( .IN1(P1_N2309), .IN2(n6888), .Q(n12425) );
  AND2X1 U14077 ( .IN1(P1_N3055), .IN2(n6907), .Q(n12426) );
  AND2X1 U14078 ( .IN1(n12428), .IN2(n6878), .Q(n12427) );
  AND2X1 U14079 ( .IN1(n12430), .IN2(P1_N291), .Q(n12429) );
  AND2X1 U14080 ( .IN1(n12432), .IN2(n6962), .Q(n12431) );
  AND2X1 U14081 ( .IN1(n12434), .IN2(n6959), .Q(n12433) );
  AND2X1 U14082 ( .IN1(P1_N3428), .IN2(n6888), .Q(n12435) );
  AND2X1 U14083 ( .IN1(P1_N4174), .IN2(n6907), .Q(n12436) );
  AND2X1 U14084 ( .IN1(P1_N3801), .IN2(n6888), .Q(n12437) );
  AND2X1 U14085 ( .IN1(P1_N4547), .IN2(n6907), .Q(n12438) );
  AND2X1 U14086 ( .IN1(n12440), .IN2(n6878), .Q(n12439) );
  AND2X1 U14087 ( .IN1(n12442), .IN2(P1_N291), .Q(n12441) );
  AND2X1 U14088 ( .IN1(P1_N387), .IN2(n11309), .Q(n12443) );
  AND2X1 U14089 ( .IN1(P1_N4810), .IN2(n6992), .Q(n12444) );
  AND2X1 U14090 ( .IN1(n12446), .IN2(n6962), .Q(n12445) );
  AND2X1 U14091 ( .IN1(n12448), .IN2(n6959), .Q(n12447) );
  AND2X1 U14092 ( .IN1(n12449), .IN2(n6980), .Q(n11361) );
  AND2X1 U14093 ( .IN1(n12450), .IN2(n6977), .Q(n11362) );
  AND2X1 U14094 ( .IN1(P1_N963), .IN2(n6904), .Q(n12451) );
  AND2X1 U14095 ( .IN1(P1_N1309), .IN2(n6907), .Q(n12452) );
  AND2X1 U14096 ( .IN1(P1_N1035), .IN2(n6888), .Q(n12453) );
  AND2X1 U14097 ( .IN1(P1_N1564), .IN2(n6907), .Q(n12454) );
  AND2X1 U14098 ( .IN1(n12456), .IN2(n6878), .Q(n12455) );
  AND2X1 U14099 ( .IN1(n12458), .IN2(P1_N291), .Q(n12457) );
  AND2X1 U14100 ( .IN1(P1_N1937), .IN2(n6882), .Q(n12459) );
  AND2X1 U14101 ( .IN1(P1_N2683), .IN2(n6881), .Q(n12460) );
  AND2X1 U14102 ( .IN1(P1_N2310), .IN2(n6882), .Q(n12461) );
  AND2X1 U14103 ( .IN1(P1_N3056), .IN2(n6881), .Q(n12462) );
  AND2X1 U14104 ( .IN1(n12464), .IN2(n6856), .Q(n12463) );
  AND2X1 U14105 ( .IN1(n12466), .IN2(n6855), .Q(n12465) );
  AND2X1 U14106 ( .IN1(n12468), .IN2(n6962), .Q(n12467) );
  AND2X1 U14107 ( .IN1(n12470), .IN2(n6957), .Q(n12469) );
  AND2X1 U14108 ( .IN1(P1_N3429), .IN2(n6882), .Q(n12471) );
  AND2X1 U14109 ( .IN1(P1_N4175), .IN2(n6881), .Q(n12472) );
  AND2X1 U14110 ( .IN1(P1_N3802), .IN2(n6882), .Q(n12473) );
  AND2X1 U14111 ( .IN1(P1_N4548), .IN2(n6881), .Q(n12474) );
  AND2X1 U14112 ( .IN1(n12476), .IN2(n6856), .Q(n12475) );
  AND2X1 U14113 ( .IN1(n12478), .IN2(n6855), .Q(n12477) );
  AND2X1 U14114 ( .IN1(P1_N388), .IN2(n11309), .Q(n12479) );
  AND2X1 U14115 ( .IN1(P1_N4811), .IN2(n6992), .Q(n12480) );
  AND2X1 U14116 ( .IN1(n12482), .IN2(n6952), .Q(n12481) );
  AND2X1 U14117 ( .IN1(n12484), .IN2(n6959), .Q(n12483) );
  AND2X1 U14118 ( .IN1(n12485), .IN2(n6976), .Q(n11363) );
  AND2X1 U14119 ( .IN1(n12486), .IN2(n6977), .Q(n11364) );
  AND2X1 U14120 ( .IN1(P1_N964), .IN2(n6882), .Q(n12487) );
  AND2X1 U14121 ( .IN1(P1_N1310), .IN2(n6881), .Q(n12488) );
  AND2X1 U14122 ( .IN1(P1_N1036), .IN2(n6882), .Q(n12489) );
  AND2X1 U14123 ( .IN1(P1_N1565), .IN2(n6881), .Q(n12490) );
  AND2X1 U14124 ( .IN1(n12492), .IN2(n6856), .Q(n12491) );
  AND2X1 U14125 ( .IN1(n12494), .IN2(n6855), .Q(n12493) );
  AND2X1 U14126 ( .IN1(P1_N1938), .IN2(n6882), .Q(n12495) );
  AND2X1 U14127 ( .IN1(P1_N2684), .IN2(n6881), .Q(n12496) );
  AND2X1 U14128 ( .IN1(P1_N2311), .IN2(n6882), .Q(n12497) );
  AND2X1 U14129 ( .IN1(P1_N3057), .IN2(n6881), .Q(n12498) );
  AND2X1 U14130 ( .IN1(n12500), .IN2(n6856), .Q(n12499) );
  AND2X1 U14131 ( .IN1(n12502), .IN2(n6855), .Q(n12501) );
  AND2X1 U14132 ( .IN1(n12504), .IN2(n6952), .Q(n12503) );
  AND2X1 U14133 ( .IN1(n12506), .IN2(n6957), .Q(n12505) );
  AND2X1 U14134 ( .IN1(P1_N3430), .IN2(n6882), .Q(n12507) );
  AND2X1 U14135 ( .IN1(P1_N4176), .IN2(n6881), .Q(n12508) );
  AND2X1 U14136 ( .IN1(P1_N3803), .IN2(n6882), .Q(n12509) );
  AND2X1 U14137 ( .IN1(P1_N4549), .IN2(n6881), .Q(n12510) );
  AND2X1 U14138 ( .IN1(n12512), .IN2(n6856), .Q(n12511) );
  AND2X1 U14139 ( .IN1(n12514), .IN2(n6855), .Q(n12513) );
  AND2X1 U14140 ( .IN1(P1_N389), .IN2(n11309), .Q(n12515) );
  AND2X1 U14141 ( .IN1(P1_N4812), .IN2(n6992), .Q(n12516) );
  AND2X1 U14142 ( .IN1(n12518), .IN2(n6952), .Q(n12517) );
  AND2X1 U14143 ( .IN1(n12520), .IN2(n6959), .Q(n12519) );
  AND2X1 U14144 ( .IN1(n12521), .IN2(n6976), .Q(n11365) );
  AND2X1 U14145 ( .IN1(n12522), .IN2(n6977), .Q(n11366) );
  AND2X1 U14146 ( .IN1(P1_N965), .IN2(n6882), .Q(n12523) );
  AND2X1 U14147 ( .IN1(P1_N1311), .IN2(n6881), .Q(n12524) );
  AND2X1 U14148 ( .IN1(P1_N1037), .IN2(n6882), .Q(n12525) );
  AND2X1 U14149 ( .IN1(P1_N1566), .IN2(n6881), .Q(n12526) );
  AND2X1 U14150 ( .IN1(n12528), .IN2(n6856), .Q(n12527) );
  AND2X1 U14151 ( .IN1(n12530), .IN2(n6855), .Q(n12529) );
  AND2X1 U14152 ( .IN1(P1_N1939), .IN2(n6882), .Q(n12531) );
  AND2X1 U14153 ( .IN1(P1_N2685), .IN2(n6881), .Q(n12532) );
  AND2X1 U14154 ( .IN1(P1_N2312), .IN2(n6882), .Q(n12533) );
  AND2X1 U14155 ( .IN1(P1_N3058), .IN2(n6881), .Q(n12534) );
  AND2X1 U14156 ( .IN1(n12536), .IN2(n6856), .Q(n12535) );
  AND2X1 U14157 ( .IN1(n12538), .IN2(n6855), .Q(n12537) );
  AND2X1 U14158 ( .IN1(n12540), .IN2(n6952), .Q(n12539) );
  AND2X1 U14159 ( .IN1(n12542), .IN2(n6959), .Q(n12541) );
  AND2X1 U14160 ( .IN1(P1_N3431), .IN2(n6882), .Q(n12543) );
  AND2X1 U14161 ( .IN1(P1_N4177), .IN2(n6881), .Q(n12544) );
  AND2X1 U14162 ( .IN1(P1_N3804), .IN2(n6882), .Q(n12545) );
  AND2X1 U14163 ( .IN1(P1_N4550), .IN2(n6881), .Q(n12546) );
  AND2X1 U14164 ( .IN1(n12548), .IN2(n6856), .Q(n12547) );
  AND2X1 U14165 ( .IN1(n12550), .IN2(n6855), .Q(n12549) );
  AND2X1 U13980 ( .IN1(P1_N3797), .IN2(n6894), .Q(n12293) );
  AND2X1 U13981 ( .IN1(P1_N4543), .IN2(n6893), .Q(n12294) );
  AND2X1 U13982 ( .IN1(n12296), .IN2(n6870), .Q(n12295) );
  AND2X1 U13983 ( .IN1(n12298), .IN2(n6869), .Q(n12297) );
  AND2X1 U13984 ( .IN1(P1_N383), .IN2(n11309), .Q(n12299) );
  AND2X1 U13985 ( .IN1(P1_N4806), .IN2(n6992), .Q(n12300) );
  AND2X1 U13986 ( .IN1(n12302), .IN2(n6958), .Q(n12301) );
  AND2X1 U13987 ( .IN1(n12304), .IN2(n6949), .Q(n12303) );
  AND2X1 U13988 ( .IN1(n12305), .IN2(n6980), .Q(n11353) );
  AND2X1 U13989 ( .IN1(n12306), .IN2(n6979), .Q(n11354) );
  AND2X1 U13990 ( .IN1(P1_N959), .IN2(n6896), .Q(n12307) );
  AND2X1 U13991 ( .IN1(P1_N1305), .IN2(n6895), .Q(n12308) );
  AND2X1 U13992 ( .IN1(P1_N1031), .IN2(n6896), .Q(n12309) );
  AND2X1 U13993 ( .IN1(P1_N1560), .IN2(n6895), .Q(n12310) );
  AND2X1 U13994 ( .IN1(n12312), .IN2(n6870), .Q(n12311) );
  AND2X1 U13995 ( .IN1(n12314), .IN2(n6869), .Q(n12313) );
  AND2X1 U13996 ( .IN1(P1_N1933), .IN2(n6894), .Q(n12315) );
  AND2X1 U13997 ( .IN1(P1_N2679), .IN2(n6893), .Q(n12316) );
  AND2X1 U13998 ( .IN1(P1_N2306), .IN2(n6896), .Q(n12317) );
  AND2X1 U13999 ( .IN1(P1_N3052), .IN2(n6895), .Q(n12318) );
  AND2X1 U14000 ( .IN1(n12320), .IN2(n6870), .Q(n12319) );
  AND2X1 U14001 ( .IN1(n12322), .IN2(n6869), .Q(n12321) );
  AND2X1 U14002 ( .IN1(n12324), .IN2(n6958), .Q(n12323) );
  AND2X1 U14003 ( .IN1(n12326), .IN2(n6949), .Q(n12325) );
  AND2X1 U14004 ( .IN1(P1_N3425), .IN2(n6896), .Q(n12327) );
  AND2X1 U14005 ( .IN1(P1_N4171), .IN2(n6895), .Q(n12328) );
  AND2X1 U14006 ( .IN1(P1_N3798), .IN2(n6896), .Q(n12329) );
  AND2X1 U14007 ( .IN1(P1_N4544), .IN2(n6895), .Q(n12330) );
  AND2X1 U14008 ( .IN1(n12332), .IN2(n6856), .Q(n12331) );
  AND2X1 U14009 ( .IN1(n12334), .IN2(n6857), .Q(n12333) );
  AND2X1 U14010 ( .IN1(P1_N384), .IN2(n11309), .Q(n12335) );
  AND2X1 U14011 ( .IN1(P1_N4807), .IN2(n6992), .Q(n12336) );
  AND2X1 U14012 ( .IN1(n12338), .IN2(n6956), .Q(n12337) );
  AND2X1 U14013 ( .IN1(n12340), .IN2(n6949), .Q(n12339) );
  AND2X1 U14014 ( .IN1(n12341), .IN2(n6980), .Q(n11355) );
  AND2X1 U14015 ( .IN1(n12342), .IN2(n6979), .Q(n11356) );
  AND2X1 U14016 ( .IN1(P1_N960), .IN2(n6884), .Q(n12343) );
  AND2X1 U14017 ( .IN1(P1_N1306), .IN2(n6883), .Q(n12344) );
  AND2X1 U14018 ( .IN1(P1_N1032), .IN2(n6884), .Q(n12345) );
  AND2X1 U14019 ( .IN1(P1_N1561), .IN2(n6883), .Q(n12346) );
  AND2X1 U14020 ( .IN1(n12348), .IN2(n6856), .Q(n12347) );
  AND2X1 U14021 ( .IN1(n12350), .IN2(n6857), .Q(n12349) );
  AND2X1 U14022 ( .IN1(P1_N1934), .IN2(n6884), .Q(n12351) );
  AND2X1 U14023 ( .IN1(P1_N2680), .IN2(n6883), .Q(n12352) );
  AND2X1 U14024 ( .IN1(P1_N2307), .IN2(n6884), .Q(n12353) );
  AND2X1 U14025 ( .IN1(P1_N3053), .IN2(n6883), .Q(n12354) );
  AND2X1 U14026 ( .IN1(n12356), .IN2(n6856), .Q(n12355) );
  AND2X1 U14027 ( .IN1(n12358), .IN2(n6857), .Q(n12357) );
  AND2X1 U14028 ( .IN1(n12360), .IN2(n6956), .Q(n12359) );
  AND2X1 U14029 ( .IN1(n12362), .IN2(n6949), .Q(n12361) );
  AND2X1 U14030 ( .IN1(P1_N3426), .IN2(n6884), .Q(n12363) );
  AND2X1 U14031 ( .IN1(P1_N4172), .IN2(n6883), .Q(n12364) );
  AND2X1 U14032 ( .IN1(P1_N3799), .IN2(n6884), .Q(n12365) );
  AND2X1 U14033 ( .IN1(P1_N4545), .IN2(n6883), .Q(n12366) );
  AND2X1 U14034 ( .IN1(n12368), .IN2(n6864), .Q(n12367) );
  AND2X1 U14035 ( .IN1(n12370), .IN2(n6857), .Q(n12369) );
  AND2X1 U14036 ( .IN1(P1_N385), .IN2(n11309), .Q(n12371) );
  AND2X1 U14037 ( .IN1(P1_N4808), .IN2(n6992), .Q(n12372) );
  AND2X1 U14038 ( .IN1(n12374), .IN2(n6962), .Q(n12373) );
  AND2X1 U14039 ( .IN1(n12376), .IN2(n6949), .Q(n12375) );
  AND2X1 U14040 ( .IN1(n12377), .IN2(n6980), .Q(n11357) );
  AND2X1 U14041 ( .IN1(n12378), .IN2(n6979), .Q(n11358) );
  AND2X1 U14042 ( .IN1(P1_N961), .IN2(n6884), .Q(n12379) );
  AND2X1 U14043 ( .IN1(P1_N1307), .IN2(n6883), .Q(n12380) );
  AND2X1 U14044 ( .IN1(P1_N1033), .IN2(n6884), .Q(n12381) );
  AND2X1 U14045 ( .IN1(P1_N1562), .IN2(n6883), .Q(n12382) );
  AND2X1 U14046 ( .IN1(n12384), .IN2(n6864), .Q(n12383) );
  AND2X1 U14047 ( .IN1(n12386), .IN2(n6857), .Q(n12385) );
  AND2X1 U14048 ( .IN1(P1_N1935), .IN2(n6884), .Q(n12387) );
  AND2X1 U14049 ( .IN1(P1_N2681), .IN2(n6883), .Q(n12388) );
  AND2X1 U14050 ( .IN1(P1_N2308), .IN2(n6888), .Q(n12389) );
  AND2X1 U14051 ( .IN1(P1_N3054), .IN2(n6907), .Q(n12390) );
  AND2X1 U14052 ( .IN1(n12392), .IN2(n6864), .Q(n12391) );
  AND2X1 U14053 ( .IN1(n12394), .IN2(P1_N291), .Q(n12393) );
  AND2X1 U14054 ( .IN1(n12396), .IN2(n6962), .Q(n12395) );
  AND2X1 U14055 ( .IN1(n12398), .IN2(n6959), .Q(n12397) );
  AND2X1 U14056 ( .IN1(P1_N3427), .IN2(n6884), .Q(n12399) );
  AND2X1 U14057 ( .IN1(P1_N4173), .IN2(n6883), .Q(n12400) );
  AND2X1 U14058 ( .IN1(P1_N3800), .IN2(n6888), .Q(n12401) );
  AND2X1 U14059 ( .IN1(P1_N4546), .IN2(n6907), .Q(n12402) );
  AND2X1 U14060 ( .IN1(n12404), .IN2(n6878), .Q(n12403) );
  AND2X1 U14061 ( .IN1(n12406), .IN2(P1_N291), .Q(n12405) );
  AND2X1 U14062 ( .IN1(P1_N386), .IN2(n11309), .Q(n12407) );
  AND2X1 U14063 ( .IN1(P1_N4809), .IN2(n6992), .Q(n12408) );
  AND2X1 U14064 ( .IN1(n12410), .IN2(n6962), .Q(n12409) );
  AND2X1 U14065 ( .IN1(n12412), .IN2(n6959), .Q(n12411) );
  AND2X1 U14066 ( .IN1(n12413), .IN2(n6980), .Q(n11359) );
  AND2X1 U14067 ( .IN1(n12414), .IN2(n6979), .Q(n11360) );
  AND2X1 U14068 ( .IN1(P1_N962), .IN2(n6888), .Q(n12415) );
  AND2X1 U14069 ( .IN1(P1_N1308), .IN2(n6907), .Q(n12416) );
  AND2X1 U14070 ( .IN1(P1_N1034), .IN2(n6888), .Q(n12417) );
  AND2X1 U14071 ( .IN1(P1_N1563), .IN2(n6907), .Q(n12418) );
  AND2X1 U14072 ( .IN1(n12420), .IN2(n6878), .Q(n12419) );
  AND2X1 U13887 ( .IN1(P1_N1301), .IN2(n6919), .Q(n12164) );
  AND2X1 U13888 ( .IN1(P1_N1027), .IN2(n6890), .Q(n12165) );
  AND2X1 U13889 ( .IN1(P1_N1556), .IN2(n6919), .Q(n12166) );
  AND2X1 U13890 ( .IN1(n12168), .IN2(n6854), .Q(n12167) );
  AND2X1 U13891 ( .IN1(n12170), .IN2(n7459), .Q(n12169) );
  AND2X1 U13892 ( .IN1(P1_N1929), .IN2(n6890), .Q(n12171) );
  AND2X1 U13893 ( .IN1(P1_N2675), .IN2(n6919), .Q(n12172) );
  AND2X1 U13894 ( .IN1(P1_N2302), .IN2(n6920), .Q(n12173) );
  AND2X1 U13895 ( .IN1(P1_N3048), .IN2(n6901), .Q(n12174) );
  AND2X1 U13896 ( .IN1(n12176), .IN2(n6866), .Q(n12175) );
  AND2X1 U13897 ( .IN1(n12178), .IN2(n6865), .Q(n12177) );
  AND2X1 U13898 ( .IN1(n12180), .IN2(n6956), .Q(n12179) );
  AND2X1 U13899 ( .IN1(n12182), .IN2(n6955), .Q(n12181) );
  AND2X1 U13900 ( .IN1(P1_N3421), .IN2(n6890), .Q(n12183) );
  AND2X1 U13901 ( .IN1(P1_N4167), .IN2(n6919), .Q(n12184) );
  AND2X1 U13902 ( .IN1(P1_N3794), .IN2(n6920), .Q(n12185) );
  AND2X1 U13903 ( .IN1(P1_N4540), .IN2(n6919), .Q(n12186) );
  AND2X1 U13904 ( .IN1(n12188), .IN2(n6866), .Q(n12187) );
  AND2X1 U13905 ( .IN1(n12190), .IN2(n6865), .Q(n12189) );
  AND2X1 U13906 ( .IN1(P1_N380), .IN2(n11309), .Q(n12191) );
  AND2X1 U13907 ( .IN1(P1_N4803), .IN2(n6992), .Q(n12192) );
  AND2X1 U13908 ( .IN1(n12194), .IN2(n6956), .Q(n12193) );
  AND2X1 U13909 ( .IN1(n12196), .IN2(n6955), .Q(n12195) );
  AND2X1 U13910 ( .IN1(n12197), .IN2(n6976), .Q(n11347) );
  AND2X1 U13911 ( .IN1(n12198), .IN2(n6975), .Q(n11348) );
  AND2X1 U13912 ( .IN1(P1_N956), .IN2(n6904), .Q(n12199) );
  AND2X1 U13913 ( .IN1(P1_N1302), .IN2(n6919), .Q(n12200) );
  AND2X1 U13914 ( .IN1(P1_N1028), .IN2(n6904), .Q(n12201) );
  AND2X1 U13915 ( .IN1(P1_N1557), .IN2(n6919), .Q(n12202) );
  AND2X1 U13916 ( .IN1(n12204), .IN2(n6854), .Q(n12203) );
  AND2X1 U13917 ( .IN1(n12206), .IN2(n7459), .Q(n12205) );
  AND2X1 U13918 ( .IN1(P1_N1930), .IN2(n6920), .Q(n12207) );
  AND2X1 U13919 ( .IN1(P1_N2676), .IN2(n6919), .Q(n12208) );
  AND2X1 U13920 ( .IN1(P1_N2303), .IN2(n6920), .Q(n12209) );
  AND2X1 U13921 ( .IN1(P1_N3049), .IN2(n6919), .Q(n12210) );
  AND2X1 U13922 ( .IN1(n12212), .IN2(n6866), .Q(n12211) );
  AND2X1 U13923 ( .IN1(n12214), .IN2(n6865), .Q(n12213) );
  AND2X1 U13924 ( .IN1(n12216), .IN2(n6956), .Q(n12215) );
  AND2X1 U13925 ( .IN1(n12218), .IN2(n6955), .Q(n12217) );
  AND2X1 U13926 ( .IN1(P1_N3422), .IN2(n6910), .Q(n12219) );
  AND2X1 U13927 ( .IN1(P1_N4168), .IN2(n6887), .Q(n12220) );
  AND2X1 U13928 ( .IN1(P1_N3795), .IN2(n6904), .Q(n12221) );
  AND2X1 U13929 ( .IN1(P1_N4541), .IN2(n6887), .Q(n12222) );
  AND2X1 U13930 ( .IN1(n12224), .IN2(n6854), .Q(n12223) );
  AND2X1 U13931 ( .IN1(n12226), .IN2(n7459), .Q(n12225) );
  AND2X1 U13932 ( .IN1(P1_N381), .IN2(n11309), .Q(n12227) );
  AND2X1 U13933 ( .IN1(P1_N4804), .IN2(n6992), .Q(n12228) );
  AND2X1 U13934 ( .IN1(n12230), .IN2(n6956), .Q(n12229) );
  AND2X1 U13935 ( .IN1(n12232), .IN2(n6955), .Q(n12231) );
  AND2X1 U13936 ( .IN1(n12233), .IN2(n6976), .Q(n11349) );
  AND2X1 U13937 ( .IN1(n12234), .IN2(n6975), .Q(n11350) );
  AND2X1 U13938 ( .IN1(P1_N957), .IN2(n6904), .Q(n12235) );
  AND2X1 U13939 ( .IN1(P1_N1303), .IN2(n6887), .Q(n12236) );
  AND2X1 U13940 ( .IN1(P1_N1029), .IN2(n6910), .Q(n12237) );
  AND2X1 U13941 ( .IN1(P1_N1558), .IN2(n6887), .Q(n12238) );
  AND2X1 U13942 ( .IN1(n12240), .IN2(n6854), .Q(n12239) );
  AND2X1 U13943 ( .IN1(n12242), .IN2(n7459), .Q(n12241) );
  AND2X1 U13944 ( .IN1(P1_N1931), .IN2(n6904), .Q(n12243) );
  AND2X1 U13945 ( .IN1(P1_N2677), .IN2(n6887), .Q(n12244) );
  AND2X1 U13946 ( .IN1(P1_N2304), .IN2(n6904), .Q(n12245) );
  AND2X1 U13947 ( .IN1(P1_N3050), .IN2(n6887), .Q(n12246) );
  AND2X1 U13948 ( .IN1(n12248), .IN2(n6854), .Q(n12247) );
  AND2X1 U13949 ( .IN1(n12250), .IN2(n7459), .Q(n12249) );
  AND2X1 U13950 ( .IN1(n12252), .IN2(n6956), .Q(n12251) );
  AND2X1 U13951 ( .IN1(n12254), .IN2(n6955), .Q(n12253) );
  AND2X1 U13952 ( .IN1(P1_N3423), .IN2(n6904), .Q(n12255) );
  AND2X1 U13953 ( .IN1(P1_N4169), .IN2(n6887), .Q(n12256) );
  AND2X1 U13954 ( .IN1(P1_N3796), .IN2(n6894), .Q(n12257) );
  AND2X1 U13955 ( .IN1(P1_N4542), .IN2(n6893), .Q(n12258) );
  AND2X1 U13956 ( .IN1(n12260), .IN2(n6870), .Q(n12259) );
  AND2X1 U13957 ( .IN1(n12262), .IN2(n6869), .Q(n12261) );
  AND2X1 U13958 ( .IN1(P1_N382), .IN2(n11309), .Q(n12263) );
  AND2X1 U13959 ( .IN1(P1_N4805), .IN2(n6992), .Q(n12264) );
  AND2X1 U13960 ( .IN1(n12266), .IN2(n6958), .Q(n12265) );
  AND2X1 U13961 ( .IN1(n12268), .IN2(n6949), .Q(n12267) );
  AND2X1 U13962 ( .IN1(n12269), .IN2(n6976), .Q(n11351) );
  AND2X1 U13963 ( .IN1(n12270), .IN2(n6979), .Q(n11352) );
  AND2X1 U13964 ( .IN1(P1_N958), .IN2(n6896), .Q(n12271) );
  AND2X1 U13965 ( .IN1(P1_N1304), .IN2(n6893), .Q(n12272) );
  AND2X1 U13966 ( .IN1(P1_N1030), .IN2(n6894), .Q(n12273) );
  AND2X1 U13967 ( .IN1(P1_N1559), .IN2(n6893), .Q(n12274) );
  AND2X1 U13968 ( .IN1(n12276), .IN2(n6870), .Q(n12275) );
  AND2X1 U13969 ( .IN1(n12278), .IN2(n6869), .Q(n12277) );
  AND2X1 U13970 ( .IN1(P1_N1932), .IN2(n6894), .Q(n12279) );
  AND2X1 U13971 ( .IN1(P1_N2678), .IN2(n6893), .Q(n12280) );
  AND2X1 U13972 ( .IN1(P1_N2305), .IN2(n6894), .Q(n12281) );
  AND2X1 U13973 ( .IN1(P1_N3051), .IN2(n6893), .Q(n12282) );
  AND2X1 U13974 ( .IN1(n12284), .IN2(n6870), .Q(n12283) );
  AND2X1 U13975 ( .IN1(n12286), .IN2(n6869), .Q(n12285) );
  AND2X1 U13976 ( .IN1(n12288), .IN2(n6956), .Q(n12287) );
  AND2X1 U13977 ( .IN1(n12290), .IN2(n6949), .Q(n12289) );
  AND2X1 U13978 ( .IN1(P1_N3424), .IN2(n6894), .Q(n12291) );
  AND2X1 U13979 ( .IN1(P1_N4170), .IN2(n6893), .Q(n12292) );
  AND2X1 U13794 ( .IN1(n12036), .IN2(n6958), .Q(n12035) );
  AND2X1 U13795 ( .IN1(n12038), .IN2(n6957), .Q(n12037) );
  AND2X1 U13796 ( .IN1(P1_N3417), .IN2(n6920), .Q(n12039) );
  AND2X1 U13797 ( .IN1(P1_N4163), .IN2(n6919), .Q(n12040) );
  AND2X1 U13798 ( .IN1(P1_N3790), .IN2(n6890), .Q(n12041) );
  AND2X1 U13799 ( .IN1(P1_N4536), .IN2(n6901), .Q(n12042) );
  AND2X1 U13800 ( .IN1(n12044), .IN2(n6872), .Q(n12043) );
  AND2X1 U13801 ( .IN1(n12046), .IN2(n6871), .Q(n12045) );
  AND2X1 U13802 ( .IN1(P1_N376), .IN2(n11309), .Q(n12047) );
  AND2X1 U13803 ( .IN1(P1_N4799), .IN2(n6992), .Q(n12048) );
  AND2X1 U13804 ( .IN1(n12050), .IN2(n6958), .Q(n12049) );
  AND2X1 U13805 ( .IN1(n12052), .IN2(n6957), .Q(n12051) );
  AND2X1 U13806 ( .IN1(n12053), .IN2(n6976), .Q(n11339) );
  AND2X1 U13807 ( .IN1(n12054), .IN2(n6975), .Q(n11340) );
  AND2X1 U13808 ( .IN1(P1_N952), .IN2(n6920), .Q(n12055) );
  AND2X1 U13809 ( .IN1(P1_N1298), .IN2(n6901), .Q(n12056) );
  AND2X1 U13810 ( .IN1(P1_N1024), .IN2(n6892), .Q(n12057) );
  AND2X1 U13811 ( .IN1(P1_N1553), .IN2(n6901), .Q(n12058) );
  AND2X1 U13812 ( .IN1(n12060), .IN2(n6866), .Q(n12059) );
  AND2X1 U13813 ( .IN1(n12062), .IN2(n6865), .Q(n12061) );
  AND2X1 U13814 ( .IN1(P1_N1926), .IN2(n6920), .Q(n12063) );
  AND2X1 U13815 ( .IN1(P1_N2672), .IN2(n6901), .Q(n12064) );
  AND2X1 U13816 ( .IN1(P1_N2299), .IN2(n6920), .Q(n12065) );
  AND2X1 U13817 ( .IN1(P1_N3045), .IN2(n6901), .Q(n12066) );
  AND2X1 U13818 ( .IN1(n12068), .IN2(n6866), .Q(n12067) );
  AND2X1 U13819 ( .IN1(n12070), .IN2(n6865), .Q(n12069) );
  AND2X1 U13820 ( .IN1(n12072), .IN2(n6958), .Q(n12071) );
  AND2X1 U13821 ( .IN1(n12074), .IN2(n6957), .Q(n12073) );
  AND2X1 U13822 ( .IN1(P1_N3418), .IN2(n6920), .Q(n12075) );
  AND2X1 U13823 ( .IN1(P1_N4164), .IN2(n6901), .Q(n12076) );
  AND2X1 U13824 ( .IN1(P1_N3791), .IN2(n6890), .Q(n12077) );
  AND2X1 U13825 ( .IN1(P1_N4537), .IN2(n6901), .Q(n12078) );
  AND2X1 U13826 ( .IN1(n12080), .IN2(n6866), .Q(n12079) );
  AND2X1 U13827 ( .IN1(n12082), .IN2(n6865), .Q(n12081) );
  AND2X1 U13828 ( .IN1(P1_N377), .IN2(n11309), .Q(n12083) );
  AND2X1 U13829 ( .IN1(P1_N4800), .IN2(n6992), .Q(n12084) );
  AND2X1 U13830 ( .IN1(n12086), .IN2(n6958), .Q(n12085) );
  AND2X1 U13831 ( .IN1(n12088), .IN2(n6957), .Q(n12087) );
  AND2X1 U13832 ( .IN1(n12089), .IN2(n6976), .Q(n11341) );
  AND2X1 U13833 ( .IN1(n12090), .IN2(n6975), .Q(n11342) );
  AND2X1 U13834 ( .IN1(P1_N953), .IN2(n6890), .Q(n12091) );
  AND2X1 U13835 ( .IN1(P1_N1299), .IN2(n6901), .Q(n12092) );
  AND2X1 U13836 ( .IN1(P1_N1025), .IN2(n6890), .Q(n12093) );
  AND2X1 U13837 ( .IN1(P1_N1554), .IN2(n6901), .Q(n12094) );
  AND2X1 U13838 ( .IN1(n12096), .IN2(n6866), .Q(n12095) );
  AND2X1 U13839 ( .IN1(n12098), .IN2(n6865), .Q(n12097) );
  AND2X1 U13840 ( .IN1(P1_N1927), .IN2(n6920), .Q(n12099) );
  AND2X1 U13841 ( .IN1(P1_N2673), .IN2(n6901), .Q(n12100) );
  AND2X1 U13842 ( .IN1(P1_N2300), .IN2(n6920), .Q(n12101) );
  AND2X1 U13843 ( .IN1(P1_N3046), .IN2(n6901), .Q(n12102) );
  AND2X1 U13844 ( .IN1(n12104), .IN2(n6866), .Q(n12103) );
  AND2X1 U13845 ( .IN1(n12106), .IN2(n6865), .Q(n12105) );
  AND2X1 U13846 ( .IN1(n12108), .IN2(n6958), .Q(n12107) );
  AND2X1 U13847 ( .IN1(n12110), .IN2(n6957), .Q(n12109) );
  AND2X1 U13848 ( .IN1(P1_N3419), .IN2(n6920), .Q(n12111) );
  AND2X1 U13849 ( .IN1(P1_N4165), .IN2(n6901), .Q(n12112) );
  AND2X1 U13850 ( .IN1(P1_N3792), .IN2(n6920), .Q(n12113) );
  AND2X1 U13851 ( .IN1(P1_N4538), .IN2(n6901), .Q(n12114) );
  AND2X1 U13852 ( .IN1(n12116), .IN2(n6866), .Q(n12115) );
  AND2X1 U13853 ( .IN1(n12118), .IN2(n6865), .Q(n12117) );
  AND2X1 U13854 ( .IN1(P1_N378), .IN2(n11309), .Q(n12119) );
  AND2X1 U13855 ( .IN1(P1_N4801), .IN2(n6992), .Q(n12120) );
  AND2X1 U13856 ( .IN1(n12122), .IN2(n6956), .Q(n12121) );
  AND2X1 U13857 ( .IN1(n12124), .IN2(n6955), .Q(n12123) );
  AND2X1 U13858 ( .IN1(n12125), .IN2(n6976), .Q(n11343) );
  AND2X1 U13859 ( .IN1(n12126), .IN2(n6975), .Q(n11344) );
  AND2X1 U13860 ( .IN1(P1_N954), .IN2(n6920), .Q(n12127) );
  AND2X1 U13861 ( .IN1(P1_N1300), .IN2(n6901), .Q(n12128) );
  AND2X1 U13862 ( .IN1(P1_N1026), .IN2(n6920), .Q(n12129) );
  AND2X1 U13863 ( .IN1(P1_N1555), .IN2(n6919), .Q(n12130) );
  AND2X1 U13864 ( .IN1(n12132), .IN2(n6866), .Q(n12131) );
  AND2X1 U13865 ( .IN1(n12134), .IN2(n6865), .Q(n12133) );
  AND2X1 U13866 ( .IN1(P1_N1928), .IN2(n6920), .Q(n12135) );
  AND2X1 U13867 ( .IN1(P1_N2674), .IN2(n6919), .Q(n12136) );
  AND2X1 U13868 ( .IN1(P1_N2301), .IN2(n6892), .Q(n12137) );
  AND2X1 U13869 ( .IN1(P1_N3047), .IN2(n6901), .Q(n12138) );
  AND2X1 U13870 ( .IN1(n12140), .IN2(n6866), .Q(n12139) );
  AND2X1 U13871 ( .IN1(n12142), .IN2(n6865), .Q(n12141) );
  AND2X1 U13872 ( .IN1(n12144), .IN2(n6956), .Q(n12143) );
  AND2X1 U13873 ( .IN1(n12146), .IN2(n6955), .Q(n12145) );
  AND2X1 U13874 ( .IN1(P1_N3420), .IN2(n6920), .Q(n12147) );
  AND2X1 U13875 ( .IN1(P1_N4166), .IN2(n6919), .Q(n12148) );
  AND2X1 U13876 ( .IN1(P1_N3793), .IN2(n6920), .Q(n12149) );
  AND2X1 U13877 ( .IN1(P1_N4539), .IN2(n6919), .Q(n12150) );
  AND2X1 U13878 ( .IN1(n12152), .IN2(n6866), .Q(n12151) );
  AND2X1 U13879 ( .IN1(n12154), .IN2(n6865), .Q(n12153) );
  AND2X1 U13880 ( .IN1(P1_N379), .IN2(n11309), .Q(n12155) );
  AND2X1 U13881 ( .IN1(P1_N4802), .IN2(n6992), .Q(n12156) );
  AND2X1 U13882 ( .IN1(n12158), .IN2(n6956), .Q(n12157) );
  AND2X1 U13883 ( .IN1(n12160), .IN2(n6955), .Q(n12159) );
  AND2X1 U13884 ( .IN1(n12161), .IN2(n6976), .Q(n11345) );
  AND2X1 U13885 ( .IN1(n12162), .IN2(n6975), .Q(n11346) );
  AND2X1 U13886 ( .IN1(P1_N955), .IN2(n6926), .Q(n12163) );
  AND2X1 U13701 ( .IN1(n11908), .IN2(n6961), .Q(n11907) );
  AND2X1 U13702 ( .IN1(n11909), .IN2(n6982), .Q(n11331) );
  AND2X1 U13703 ( .IN1(n11910), .IN2(n6981), .Q(n11332) );
  AND2X1 U13704 ( .IN1(P1_N948), .IN2(n6890), .Q(n11911) );
  AND2X1 U13705 ( .IN1(P1_N1294), .IN2(P1_N292), .Q(n11912) );
  AND2X1 U13706 ( .IN1(P1_N1020), .IN2(n6892), .Q(n11913) );
  AND2X1 U13707 ( .IN1(P1_N1549), .IN2(n6891), .Q(n11914) );
  AND2X1 U13708 ( .IN1(n11916), .IN2(n6872), .Q(n11915) );
  AND2X1 U13709 ( .IN1(n11918), .IN2(n6871), .Q(n11917) );
  AND2X1 U13710 ( .IN1(P1_N1922), .IN2(n6890), .Q(n11919) );
  AND2X1 U13711 ( .IN1(P1_N2668), .IN2(P1_N292), .Q(n11920) );
  AND2X1 U13712 ( .IN1(P1_N2295), .IN2(n6890), .Q(n11921) );
  AND2X1 U13713 ( .IN1(P1_N3041), .IN2(n6891), .Q(n11922) );
  AND2X1 U13714 ( .IN1(n11924), .IN2(n6872), .Q(n11923) );
  AND2X1 U13715 ( .IN1(n11926), .IN2(n6871), .Q(n11925) );
  AND2X1 U13716 ( .IN1(n11928), .IN2(n6958), .Q(n11927) );
  AND2X1 U13717 ( .IN1(n11930), .IN2(n6957), .Q(n11929) );
  AND2X1 U13718 ( .IN1(P1_N3414), .IN2(n6892), .Q(n11931) );
  AND2X1 U13719 ( .IN1(P1_N4160), .IN2(n6891), .Q(n11932) );
  AND2X1 U13720 ( .IN1(P1_N3787), .IN2(n6892), .Q(n11933) );
  AND2X1 U13721 ( .IN1(P1_N4533), .IN2(n6891), .Q(n11934) );
  AND2X1 U13722 ( .IN1(n11936), .IN2(n6872), .Q(n11935) );
  AND2X1 U13723 ( .IN1(n11938), .IN2(n6871), .Q(n11937) );
  AND2X1 U13724 ( .IN1(P1_N373), .IN2(n11309), .Q(n11939) );
  AND2X1 U13725 ( .IN1(P1_N4796), .IN2(n6992), .Q(n11940) );
  AND2X1 U13726 ( .IN1(n11942), .IN2(n6958), .Q(n11941) );
  AND2X1 U13727 ( .IN1(n11944), .IN2(n6957), .Q(n11943) );
  AND2X1 U13728 ( .IN1(n11945), .IN2(n6976), .Q(n11333) );
  AND2X1 U13729 ( .IN1(n11946), .IN2(n6975), .Q(n11334) );
  AND2X1 U13730 ( .IN1(P1_N949), .IN2(n6892), .Q(n11947) );
  AND2X1 U13731 ( .IN1(P1_N1295), .IN2(n6891), .Q(n11948) );
  AND2X1 U13732 ( .IN1(P1_N1021), .IN2(n6892), .Q(n11949) );
  AND2X1 U13733 ( .IN1(P1_N1550), .IN2(n6891), .Q(n11950) );
  AND2X1 U13734 ( .IN1(n11952), .IN2(n6872), .Q(n11951) );
  AND2X1 U13735 ( .IN1(n11954), .IN2(n6871), .Q(n11953) );
  AND2X1 U13736 ( .IN1(P1_N1923), .IN2(n6892), .Q(n11955) );
  AND2X1 U13737 ( .IN1(P1_N2669), .IN2(n6891), .Q(n11956) );
  AND2X1 U13738 ( .IN1(P1_N2296), .IN2(n6892), .Q(n11957) );
  AND2X1 U13739 ( .IN1(P1_N3042), .IN2(n6891), .Q(n11958) );
  AND2X1 U13740 ( .IN1(n11960), .IN2(n6872), .Q(n11959) );
  AND2X1 U13741 ( .IN1(n11962), .IN2(n6871), .Q(n11961) );
  AND2X1 U13742 ( .IN1(n11964), .IN2(n6958), .Q(n11963) );
  AND2X1 U13743 ( .IN1(n11966), .IN2(n6957), .Q(n11965) );
  AND2X1 U13744 ( .IN1(P1_N3415), .IN2(n6892), .Q(n11967) );
  AND2X1 U13745 ( .IN1(P1_N4161), .IN2(n6891), .Q(n11968) );
  AND2X1 U13746 ( .IN1(P1_N3788), .IN2(n6892), .Q(n11969) );
  AND2X1 U13747 ( .IN1(P1_N4534), .IN2(n6891), .Q(n11970) );
  AND2X1 U13748 ( .IN1(n11972), .IN2(n6872), .Q(n11971) );
  AND2X1 U13749 ( .IN1(n11974), .IN2(n6871), .Q(n11973) );
  AND2X1 U13750 ( .IN1(P1_N374), .IN2(n11309), .Q(n11975) );
  AND2X1 U13751 ( .IN1(P1_N4797), .IN2(n6992), .Q(n11976) );
  AND2X1 U13752 ( .IN1(n11978), .IN2(n6958), .Q(n11977) );
  AND2X1 U13753 ( .IN1(n11980), .IN2(n6957), .Q(n11979) );
  AND2X1 U13754 ( .IN1(n11981), .IN2(n6976), .Q(n11335) );
  AND2X1 U13755 ( .IN1(n11982), .IN2(n6975), .Q(n11336) );
  AND2X1 U13756 ( .IN1(P1_N950), .IN2(n6892), .Q(n11983) );
  AND2X1 U13757 ( .IN1(P1_N1296), .IN2(n6891), .Q(n11984) );
  AND2X1 U13758 ( .IN1(P1_N1022), .IN2(n6892), .Q(n11985) );
  AND2X1 U13759 ( .IN1(P1_N1551), .IN2(n6891), .Q(n11986) );
  AND2X1 U13760 ( .IN1(n11988), .IN2(n6872), .Q(n11987) );
  AND2X1 U13761 ( .IN1(n11990), .IN2(n6871), .Q(n11989) );
  AND2X1 U13762 ( .IN1(P1_N1924), .IN2(n6892), .Q(n11991) );
  AND2X1 U13763 ( .IN1(P1_N2670), .IN2(n6891), .Q(n11992) );
  AND2X1 U13764 ( .IN1(P1_N2297), .IN2(n6892), .Q(n11993) );
  AND2X1 U13765 ( .IN1(P1_N3043), .IN2(n6891), .Q(n11994) );
  AND2X1 U13766 ( .IN1(n11996), .IN2(n6872), .Q(n11995) );
  AND2X1 U13767 ( .IN1(n11998), .IN2(n6871), .Q(n11997) );
  AND2X1 U13768 ( .IN1(n12000), .IN2(n6958), .Q(n11999) );
  AND2X1 U13769 ( .IN1(n12002), .IN2(n6957), .Q(n12001) );
  AND2X1 U13770 ( .IN1(P1_N3416), .IN2(n6890), .Q(n12003) );
  AND2X1 U13771 ( .IN1(P1_N4162), .IN2(n6901), .Q(n12004) );
  AND2X1 U13772 ( .IN1(P1_N3789), .IN2(n6892), .Q(n12005) );
  AND2X1 U13773 ( .IN1(P1_N4535), .IN2(n6891), .Q(n12006) );
  AND2X1 U13774 ( .IN1(n12008), .IN2(n6872), .Q(n12007) );
  AND2X1 U13775 ( .IN1(n12010), .IN2(n6871), .Q(n12009) );
  AND2X1 U13776 ( .IN1(P1_N375), .IN2(n11309), .Q(n12011) );
  AND2X1 U13777 ( .IN1(P1_N4798), .IN2(n6992), .Q(n12012) );
  AND2X1 U13778 ( .IN1(n12014), .IN2(n6958), .Q(n12013) );
  AND2X1 U13779 ( .IN1(n12016), .IN2(n6957), .Q(n12015) );
  AND2X1 U13780 ( .IN1(n12017), .IN2(n6976), .Q(n11337) );
  AND2X1 U13781 ( .IN1(n12018), .IN2(n6975), .Q(n11338) );
  AND2X1 U13782 ( .IN1(P1_N951), .IN2(n6926), .Q(n12019) );
  AND2X1 U13783 ( .IN1(P1_N1297), .IN2(n6901), .Q(n12020) );
  AND2X1 U13784 ( .IN1(P1_N1023), .IN2(n6920), .Q(n12021) );
  AND2X1 U13785 ( .IN1(P1_N1552), .IN2(n6901), .Q(n12022) );
  AND2X1 U13786 ( .IN1(n12024), .IN2(n6872), .Q(n12023) );
  AND2X1 U13787 ( .IN1(n12026), .IN2(n6871), .Q(n12025) );
  AND2X1 U13788 ( .IN1(P1_N1925), .IN2(n6890), .Q(n12027) );
  AND2X1 U13789 ( .IN1(P1_N2671), .IN2(n6901), .Q(n12028) );
  AND2X1 U13790 ( .IN1(P1_N2298), .IN2(n6920), .Q(n12029) );
  AND2X1 U13791 ( .IN1(P1_N3044), .IN2(n6901), .Q(n12030) );
  AND2X1 U13792 ( .IN1(n12032), .IN2(n6872), .Q(n12031) );
  AND2X1 U13793 ( .IN1(n12034), .IN2(n6871), .Q(n12033) );
  AND2X1 U13608 ( .IN1(P1_N2291), .IN2(n6888), .Q(n11777) );
  AND2X1 U13609 ( .IN1(P1_N3037), .IN2(n6887), .Q(n11778) );
  AND2X1 U13610 ( .IN1(n11780), .IN2(n6874), .Q(n11779) );
  AND2X1 U13611 ( .IN1(n11782), .IN2(n7458), .Q(n11781) );
  AND2X1 U13612 ( .IN1(n11784), .IN2(n6954), .Q(n11783) );
  AND2X1 U13613 ( .IN1(n11786), .IN2(n7461), .Q(n11785) );
  AND2X1 U13614 ( .IN1(P1_N3410), .IN2(n6888), .Q(n11787) );
  AND2X1 U13615 ( .IN1(P1_N4156), .IN2(n6887), .Q(n11788) );
  AND2X1 U13616 ( .IN1(P1_N3783), .IN2(n6888), .Q(n11789) );
  AND2X1 U13617 ( .IN1(P1_N4529), .IN2(n6887), .Q(n11790) );
  AND2X1 U13618 ( .IN1(n11792), .IN2(n6874), .Q(n11791) );
  AND2X1 U13619 ( .IN1(n11794), .IN2(n7458), .Q(n11793) );
  AND2X1 U13620 ( .IN1(P1_N369), .IN2(n11309), .Q(n11795) );
  AND2X1 U13621 ( .IN1(P1_N4792), .IN2(n6992), .Q(n11796) );
  AND2X1 U13622 ( .IN1(n11798), .IN2(n6954), .Q(n11797) );
  AND2X1 U13623 ( .IN1(n11800), .IN2(n7461), .Q(n11799) );
  AND2X1 U13624 ( .IN1(n11801), .IN2(n6984), .Q(n11325) );
  AND2X1 U13625 ( .IN1(n11802), .IN2(P1_N294), .Q(n11326) );
  AND2X1 U13626 ( .IN1(P1_N945), .IN2(n6904), .Q(n11803) );
  AND2X1 U13627 ( .IN1(P1_N1291), .IN2(n7483), .Q(n11804) );
  AND2X1 U13628 ( .IN1(P1_N1017), .IN2(n6904), .Q(n11805) );
  AND2X1 U13629 ( .IN1(P1_N1546), .IN2(n7483), .Q(n11806) );
  AND2X1 U13630 ( .IN1(n11808), .IN2(n6862), .Q(n11807) );
  AND2X1 U13631 ( .IN1(n11810), .IN2(n6857), .Q(n11809) );
  AND2X1 U13632 ( .IN1(P1_N1919), .IN2(n6904), .Q(n11811) );
  AND2X1 U13633 ( .IN1(P1_N2665), .IN2(n7483), .Q(n11812) );
  AND2X1 U13634 ( .IN1(P1_N2292), .IN2(n6904), .Q(n11813) );
  AND2X1 U13635 ( .IN1(P1_N3038), .IN2(n7483), .Q(n11814) );
  AND2X1 U13636 ( .IN1(n11816), .IN2(n6864), .Q(n11815) );
  AND2X1 U13637 ( .IN1(n11818), .IN2(n6857), .Q(n11817) );
  AND2X1 U13638 ( .IN1(n11820), .IN2(n6962), .Q(n11819) );
  AND2X1 U13639 ( .IN1(n11822), .IN2(n6961), .Q(n11821) );
  AND2X1 U13640 ( .IN1(P1_N3411), .IN2(n6904), .Q(n11823) );
  AND2X1 U13641 ( .IN1(P1_N4157), .IN2(n7483), .Q(n11824) );
  AND2X1 U13642 ( .IN1(P1_N3784), .IN2(n6904), .Q(n11825) );
  AND2X1 U13643 ( .IN1(P1_N4530), .IN2(n7483), .Q(n11826) );
  AND2X1 U13644 ( .IN1(n11828), .IN2(n6864), .Q(n11827) );
  AND2X1 U13645 ( .IN1(n11830), .IN2(n6867), .Q(n11829) );
  AND2X1 U13646 ( .IN1(P1_N370), .IN2(n11309), .Q(n11831) );
  AND2X1 U13647 ( .IN1(P1_N4793), .IN2(n6992), .Q(n11832) );
  AND2X1 U13648 ( .IN1(n11834), .IN2(n6962), .Q(n11833) );
  AND2X1 U13649 ( .IN1(n11836), .IN2(n6961), .Q(n11835) );
  AND2X1 U13650 ( .IN1(n11837), .IN2(n6982), .Q(n11327) );
  AND2X1 U13651 ( .IN1(n11838), .IN2(n6981), .Q(n11328) );
  AND2X1 U13652 ( .IN1(P1_N946), .IN2(n6890), .Q(n11839) );
  AND2X1 U13653 ( .IN1(P1_N1292), .IN2(P1_N292), .Q(n11840) );
  AND2X1 U13654 ( .IN1(P1_N1018), .IN2(n6890), .Q(n11841) );
  AND2X1 U13655 ( .IN1(P1_N1547), .IN2(P1_N292), .Q(n11842) );
  AND2X1 U13656 ( .IN1(n11844), .IN2(n6864), .Q(n11843) );
  AND2X1 U13657 ( .IN1(n11846), .IN2(n6867), .Q(n11845) );
  AND2X1 U13658 ( .IN1(P1_N1920), .IN2(n6904), .Q(n11847) );
  AND2X1 U13659 ( .IN1(P1_N2666), .IN2(n7483), .Q(n11848) );
  AND2X1 U13660 ( .IN1(P1_N2293), .IN2(n6904), .Q(n11849) );
  AND2X1 U13661 ( .IN1(P1_N3039), .IN2(n7483), .Q(n11850) );
  AND2X1 U13662 ( .IN1(n11852), .IN2(n6864), .Q(n11851) );
  AND2X1 U13663 ( .IN1(n11854), .IN2(n6857), .Q(n11853) );
  AND2X1 U13664 ( .IN1(n11856), .IN2(n6962), .Q(n11855) );
  AND2X1 U13665 ( .IN1(n11858), .IN2(n6961), .Q(n11857) );
  AND2X1 U13666 ( .IN1(P1_N3412), .IN2(n6904), .Q(n11859) );
  AND2X1 U13667 ( .IN1(P1_N4158), .IN2(n7483), .Q(n11860) );
  AND2X1 U13668 ( .IN1(P1_N3785), .IN2(n6904), .Q(n11861) );
  AND2X1 U13669 ( .IN1(P1_N4531), .IN2(n7483), .Q(n11862) );
  AND2X1 U13670 ( .IN1(n11864), .IN2(n6864), .Q(n11863) );
  AND2X1 U13671 ( .IN1(n11866), .IN2(n6857), .Q(n11865) );
  AND2X1 U13672 ( .IN1(P1_N371), .IN2(n11309), .Q(n11867) );
  AND2X1 U13673 ( .IN1(P1_N4794), .IN2(n6992), .Q(n11868) );
  AND2X1 U13674 ( .IN1(n11870), .IN2(n6962), .Q(n11869) );
  AND2X1 U13675 ( .IN1(n11872), .IN2(n6961), .Q(n11871) );
  AND2X1 U13676 ( .IN1(n11873), .IN2(n6982), .Q(n11329) );
  AND2X1 U13677 ( .IN1(n11874), .IN2(n6981), .Q(n11330) );
  AND2X1 U13678 ( .IN1(P1_N947), .IN2(n6890), .Q(n11875) );
  AND2X1 U13679 ( .IN1(P1_N1293), .IN2(P1_N292), .Q(n11876) );
  AND2X1 U13680 ( .IN1(P1_N1019), .IN2(n6890), .Q(n11877) );
  AND2X1 U13681 ( .IN1(P1_N1548), .IN2(P1_N292), .Q(n11878) );
  AND2X1 U13682 ( .IN1(n11880), .IN2(n6864), .Q(n11879) );
  AND2X1 U13683 ( .IN1(n11882), .IN2(n6857), .Q(n11881) );
  AND2X1 U13684 ( .IN1(P1_N1921), .IN2(n6890), .Q(n11883) );
  AND2X1 U13685 ( .IN1(P1_N2667), .IN2(P1_N292), .Q(n11884) );
  AND2X1 U13686 ( .IN1(P1_N2294), .IN2(n6890), .Q(n11885) );
  AND2X1 U13687 ( .IN1(P1_N3040), .IN2(P1_N292), .Q(n11886) );
  AND2X1 U13688 ( .IN1(n11888), .IN2(n6864), .Q(n11887) );
  AND2X1 U13689 ( .IN1(n11890), .IN2(n6867), .Q(n11889) );
  AND2X1 U13690 ( .IN1(n11892), .IN2(n6962), .Q(n11891) );
  AND2X1 U13691 ( .IN1(n11894), .IN2(n6961), .Q(n11893) );
  AND2X1 U13692 ( .IN1(P1_N3413), .IN2(n6890), .Q(n11895) );
  AND2X1 U13693 ( .IN1(P1_N4159), .IN2(P1_N292), .Q(n11896) );
  AND2X1 U13694 ( .IN1(P1_N3786), .IN2(n6890), .Q(n11897) );
  AND2X1 U13695 ( .IN1(P1_N4532), .IN2(P1_N292), .Q(n11898) );
  AND2X1 U13696 ( .IN1(n11900), .IN2(n6864), .Q(n11899) );
  AND2X1 U13697 ( .IN1(n11902), .IN2(n6857), .Q(n11901) );
  AND2X1 U13698 ( .IN1(P1_N372), .IN2(n11309), .Q(n11903) );
  AND2X1 U13699 ( .IN1(P1_N4795), .IN2(n6992), .Q(n11904) );
  AND2X1 U13700 ( .IN1(n11906), .IN2(n6962), .Q(n11905) );
  AND2X1 U13515 ( .IN1(n11650), .IN2(n6871), .Q(n11649) );
  AND2X1 U13516 ( .IN1(n6622), .IN2(n11309), .Q(n11651) );
  AND2X1 U13517 ( .IN1(P1_N4788), .IN2(n6992), .Q(n11652) );
  AND2X1 U13518 ( .IN1(n11654), .IN2(n6954), .Q(n11653) );
  AND2X1 U13519 ( .IN1(n11656), .IN2(n7461), .Q(n11655) );
  AND2X1 U13520 ( .IN1(n11657), .IN2(n6984), .Q(n11317) );
  AND2X1 U13521 ( .IN1(n11658), .IN2(P1_N294), .Q(n11318) );
  AND2X1 U13522 ( .IN1(P1_N941), .IN2(n6886), .Q(n11659) );
  AND2X1 U13523 ( .IN1(P1_N1287), .IN2(n6921), .Q(n11660) );
  AND2X1 U13524 ( .IN1(P1_N1013), .IN2(n6886), .Q(n11661) );
  AND2X1 U13525 ( .IN1(P1_N1542), .IN2(n6881), .Q(n11662) );
  AND2X1 U13526 ( .IN1(n11664), .IN2(n6872), .Q(n11663) );
  AND2X1 U13527 ( .IN1(n11666), .IN2(n7458), .Q(n11665) );
  AND2X1 U13528 ( .IN1(P1_N1915), .IN2(n6922), .Q(n11667) );
  AND2X1 U13529 ( .IN1(P1_N2661), .IN2(n6881), .Q(n11668) );
  AND2X1 U13530 ( .IN1(P1_N2288), .IN2(n6922), .Q(n11669) );
  AND2X1 U13531 ( .IN1(P1_N3034), .IN2(n6921), .Q(n11670) );
  AND2X1 U13532 ( .IN1(n11672), .IN2(n6860), .Q(n11671) );
  AND2X1 U13533 ( .IN1(n11674), .IN2(n6865), .Q(n11673) );
  AND2X1 U13534 ( .IN1(n11676), .IN2(n6954), .Q(n11675) );
  AND2X1 U13535 ( .IN1(n11678), .IN2(n7461), .Q(n11677) );
  AND2X1 U13536 ( .IN1(P1_N3407), .IN2(n6886), .Q(n11679) );
  AND2X1 U13537 ( .IN1(P1_N4153), .IN2(n6881), .Q(n11680) );
  AND2X1 U13538 ( .IN1(P1_N3780), .IN2(n6886), .Q(n11681) );
  AND2X1 U13539 ( .IN1(P1_N4526), .IN2(n6921), .Q(n11682) );
  AND2X1 U13540 ( .IN1(n11684), .IN2(n6872), .Q(n11683) );
  AND2X1 U13541 ( .IN1(n11686), .IN2(n7458), .Q(n11685) );
  AND2X1 U13542 ( .IN1(n6623), .IN2(n11309), .Q(n11687) );
  AND2X1 U13543 ( .IN1(P1_N4789), .IN2(n6992), .Q(n11688) );
  AND2X1 U13544 ( .IN1(n11690), .IN2(n6954), .Q(n11689) );
  AND2X1 U13545 ( .IN1(n11692), .IN2(n7461), .Q(n11691) );
  AND2X1 U13546 ( .IN1(n11693), .IN2(n6984), .Q(n11319) );
  AND2X1 U13547 ( .IN1(n11694), .IN2(P1_N294), .Q(n11320) );
  AND2X1 U13548 ( .IN1(P1_N942), .IN2(n6886), .Q(n11695) );
  AND2X1 U13549 ( .IN1(P1_N1288), .IN2(n6881), .Q(n11696) );
  AND2X1 U13550 ( .IN1(P1_N1014), .IN2(n6886), .Q(n11697) );
  AND2X1 U13551 ( .IN1(P1_N1543), .IN2(n6881), .Q(n11698) );
  AND2X1 U13552 ( .IN1(n11700), .IN2(n6874), .Q(n11699) );
  AND2X1 U13553 ( .IN1(n11702), .IN2(n7458), .Q(n11701) );
  AND2X1 U13554 ( .IN1(P1_N1916), .IN2(n6886), .Q(n11703) );
  AND2X1 U13555 ( .IN1(P1_N2662), .IN2(n6921), .Q(n11704) );
  AND2X1 U13556 ( .IN1(P1_N2289), .IN2(n6922), .Q(n11705) );
  AND2X1 U13557 ( .IN1(P1_N3035), .IN2(n6921), .Q(n11706) );
  AND2X1 U13558 ( .IN1(n11708), .IN2(n6872), .Q(n11707) );
  AND2X1 U13559 ( .IN1(n11710), .IN2(n7458), .Q(n11709) );
  AND2X1 U13560 ( .IN1(n11712), .IN2(n6954), .Q(n11711) );
  AND2X1 U13561 ( .IN1(n11714), .IN2(n7461), .Q(n11713) );
  AND2X1 U13562 ( .IN1(P1_N3408), .IN2(n6886), .Q(n11715) );
  AND2X1 U13563 ( .IN1(P1_N4154), .IN2(n6881), .Q(n11716) );
  AND2X1 U13564 ( .IN1(P1_N3781), .IN2(n6886), .Q(n11717) );
  AND2X1 U13565 ( .IN1(P1_N4527), .IN2(n6921), .Q(n11718) );
  AND2X1 U13566 ( .IN1(n11720), .IN2(n6872), .Q(n11719) );
  AND2X1 U13567 ( .IN1(n11722), .IN2(n7458), .Q(n11721) );
  AND2X1 U13568 ( .IN1(n18451), .IN2(n11309), .Q(n11723) );
  AND2X1 U13569 ( .IN1(P1_N4790), .IN2(n6992), .Q(n11724) );
  AND2X1 U13570 ( .IN1(n11726), .IN2(n6954), .Q(n11725) );
  AND2X1 U13571 ( .IN1(n11728), .IN2(n7461), .Q(n11727) );
  AND2X1 U13572 ( .IN1(n11729), .IN2(n6984), .Q(n11321) );
  AND2X1 U13573 ( .IN1(n11730), .IN2(P1_N294), .Q(n11322) );
  AND2X1 U13574 ( .IN1(P1_N943), .IN2(n6888), .Q(n11731) );
  AND2X1 U13575 ( .IN1(P1_N1289), .IN2(n6887), .Q(n11732) );
  AND2X1 U13576 ( .IN1(P1_N1015), .IN2(n6888), .Q(n11733) );
  AND2X1 U13577 ( .IN1(P1_N1544), .IN2(n6887), .Q(n11734) );
  AND2X1 U13578 ( .IN1(n11736), .IN2(n6874), .Q(n11735) );
  AND2X1 U13579 ( .IN1(n11738), .IN2(n7458), .Q(n11737) );
  AND2X1 U13580 ( .IN1(P1_N1917), .IN2(n6888), .Q(n11739) );
  AND2X1 U13581 ( .IN1(P1_N2663), .IN2(n6887), .Q(n11740) );
  AND2X1 U13582 ( .IN1(P1_N2290), .IN2(n6888), .Q(n11741) );
  AND2X1 U13583 ( .IN1(P1_N3036), .IN2(n6921), .Q(n11742) );
  AND2X1 U13584 ( .IN1(n11744), .IN2(n6874), .Q(n11743) );
  AND2X1 U13585 ( .IN1(n11746), .IN2(n7458), .Q(n11745) );
  AND2X1 U13586 ( .IN1(n11748), .IN2(n6954), .Q(n11747) );
  AND2X1 U13587 ( .IN1(n11750), .IN2(n7461), .Q(n11749) );
  AND2X1 U13588 ( .IN1(P1_N3409), .IN2(n6888), .Q(n11751) );
  AND2X1 U13589 ( .IN1(P1_N4155), .IN2(n6887), .Q(n11752) );
  AND2X1 U13590 ( .IN1(P1_N3782), .IN2(n6888), .Q(n11753) );
  AND2X1 U13591 ( .IN1(P1_N4528), .IN2(n6921), .Q(n11754) );
  AND2X1 U13592 ( .IN1(n11756), .IN2(n6874), .Q(n11755) );
  AND2X1 U13593 ( .IN1(n11758), .IN2(n7458), .Q(n11757) );
  AND2X1 U13594 ( .IN1(P1_N368), .IN2(n11309), .Q(n11759) );
  AND2X1 U13595 ( .IN1(P1_N4791), .IN2(n6992), .Q(n11760) );
  AND2X1 U13596 ( .IN1(n11762), .IN2(n6954), .Q(n11761) );
  AND2X1 U13597 ( .IN1(n11764), .IN2(n7461), .Q(n11763) );
  AND2X1 U13598 ( .IN1(n11765), .IN2(n6984), .Q(n11323) );
  AND2X1 U13599 ( .IN1(n11766), .IN2(P1_N294), .Q(n11324) );
  AND2X1 U13600 ( .IN1(P1_N944), .IN2(n6888), .Q(n11767) );
  AND2X1 U13601 ( .IN1(P1_N1290), .IN2(n6887), .Q(n11768) );
  AND2X1 U13602 ( .IN1(P1_N1016), .IN2(n6888), .Q(n11769) );
  AND2X1 U13603 ( .IN1(P1_N1545), .IN2(n6887), .Q(n11770) );
  AND2X1 U13604 ( .IN1(n11772), .IN2(n6874), .Q(n11771) );
  AND2X1 U13605 ( .IN1(n11774), .IN2(n7458), .Q(n11773) );
  AND2X1 U13606 ( .IN1(P1_N1918), .IN2(n6888), .Q(n11775) );
  AND2X1 U13607 ( .IN1(P1_N2664), .IN2(n6887), .Q(n11776) );
  OR2X1 U13422 ( .IN2(n11512), .IN1(n11511), .Q(P1_N4822) );
  OR2X1 U13423 ( .IN2(n11514), .IN1(n11513), .Q(P1_N4823) );
  OR2X1 U13424 ( .IN2(n11516), .IN1(n11515), .Q(P1_N4824) );
  OR2X1 U13425 ( .IN2(n11518), .IN1(n11517), .Q(P1_N4825) );
  OR2X1 U13426 ( .IN2(n11520), .IN1(n11519), .Q(P1_N4826) );
  OR2X1 U13427 ( .IN2(n11522), .IN1(n11521), .Q(P1_N4827) );
  OR2X1 U13428 ( .IN2(n11524), .IN1(n11523), .Q(P1_N4828) );
  OR2X1 U13429 ( .IN2(n11526), .IN1(n11525), .Q(P1_N4829) );
  OR2X1 U13430 ( .IN2(n11528), .IN1(n11527), .Q(P1_N4830) );
  OR2X1 U13431 ( .IN2(n11530), .IN1(n11529), .Q(P1_N4831) );
  OR2X1 U13432 ( .IN2(n11532), .IN1(n11531), .Q(P1_N4832) );
  OR2X1 U13433 ( .IN2(n11534), .IN1(n11533), .Q(P1_N4833) );
  OR2X1 U13434 ( .IN2(n11536), .IN1(n11535), .Q(P1_N4834) );
  OR2X1 U13435 ( .IN2(n11538), .IN1(n11537), .Q(P1_N4835) );
  OR2X1 U13436 ( .IN2(n11540), .IN1(n11539), .Q(P1_N4836) );
  OR2X1 U13437 ( .IN2(n11542), .IN1(n11541), .Q(P1_N4837) );
  OR2X1 U13438 ( .IN2(n11544), .IN1(n11543), .Q(P1_N4838) );
  AND2X1 U13439 ( .IN1(n11546), .IN2(n6952), .Q(n11545) );
  OR2X1 U13440 ( .IN2(n11548), .IN1(n11547), .Q(P1_N4818) );
  AND2X1 U13441 ( .IN1(P1_N5137), .IN2(n6884), .Q(n11311) );
  AND2X1 U13442 ( .IN1(P1_N5140), .IN2(n6883), .Q(n11312) );
  AND2X1 U13443 ( .IN1(n6857), .IN2(n11550), .Q(n11549) );
  AND2X1 U13444 ( .IN1(n11310), .IN2(n6864), .Q(n11551) );
  AND2X1 U13445 ( .IN1(n14521), .IN2(n6884), .Q(n11552) );
  AND2X1 U13446 ( .IN1(P1_N5213), .IN2(n6883), .Q(n11553) );
  AND2X1 U13447 ( .IN1(P1_N5143), .IN2(n6884), .Q(n11554) );
  AND2X1 U13448 ( .IN1(P1_N5282), .IN2(n6883), .Q(n11555) );
  AND2X1 U13449 ( .IN1(n11557), .IN2(n6864), .Q(n11556) );
  AND2X1 U13450 ( .IN1(n11559), .IN2(n6857), .Q(n11558) );
  AND2X1 U13451 ( .IN1(n11561), .IN2(n6958), .Q(n11560) );
  AND2X1 U13452 ( .IN1(n6949), .IN2(n11563), .Q(n11562) );
  AND2X1 U13453 ( .IN1(P1_N5284), .IN2(n6884), .Q(n11564) );
  AND2X1 U13454 ( .IN1(P1_N5288), .IN2(n6883), .Q(n11565) );
  AND2X1 U13455 ( .IN1(P1_N5286), .IN2(n6884), .Q(n11566) );
  AND2X1 U13456 ( .IN1(P1_N5290), .IN2(n6883), .Q(n11567) );
  AND2X1 U13457 ( .IN1(n11569), .IN2(n6864), .Q(n11568) );
  AND2X1 U13458 ( .IN1(n11571), .IN2(n6857), .Q(n11570) );
  AND2X1 U13459 ( .IN1(P1_N5292), .IN2(n6884), .Q(n11572) );
  AND2X1 U13460 ( .IN1(P1_N5363), .IN2(n6883), .Q(n11573) );
  AND2X1 U13461 ( .IN1(P1_N5294), .IN2(n6884), .Q(n11574) );
  AND2X1 U13462 ( .IN1(P1_N5432), .IN2(n6883), .Q(n11575) );
  AND2X1 U13463 ( .IN1(n11577), .IN2(n6856), .Q(n11576) );
  AND2X1 U13464 ( .IN1(n11579), .IN2(n6857), .Q(n11578) );
  AND2X1 U13465 ( .IN1(n11581), .IN2(n6956), .Q(n11580) );
  AND2X1 U13466 ( .IN1(n11583), .IN2(n6949), .Q(n11582) );
  AND2X1 U13468 ( .IN1(n11585), .IN2(n6980), .Q(n11313) );
  AND2X1 U13469 ( .IN1(n6979), .IN2(n11586), .Q(n11314) );
  AND2X1 U13470 ( .IN1(P1_N939), .IN2(n6886), .Q(n11587) );
  AND2X1 U13471 ( .IN1(P1_N1285), .IN2(n6881), .Q(n11588) );
  AND2X1 U13472 ( .IN1(P1_N1011), .IN2(n6886), .Q(n11589) );
  AND2X1 U13473 ( .IN1(P1_N1540), .IN2(n6921), .Q(n11590) );
  AND2X1 U13474 ( .IN1(n11592), .IN2(n6872), .Q(n11591) );
  AND2X1 U13475 ( .IN1(n11594), .IN2(n7458), .Q(n11593) );
  AND2X1 U13476 ( .IN1(P1_N1913), .IN2(n6906), .Q(n11595) );
  AND2X1 U13477 ( .IN1(P1_N2659), .IN2(n7481), .Q(n11596) );
  AND2X1 U13478 ( .IN1(P1_N2286), .IN2(n6906), .Q(n11597) );
  AND2X1 U13479 ( .IN1(P1_N3032), .IN2(n7481), .Q(n11598) );
  AND2X1 U13480 ( .IN1(n11600), .IN2(n6860), .Q(n11599) );
  AND2X1 U13481 ( .IN1(n11602), .IN2(n6871), .Q(n11601) );
  AND2X1 U13482 ( .IN1(n11604), .IN2(n6954), .Q(n11603) );
  AND2X1 U13483 ( .IN1(n11606), .IN2(n7461), .Q(n11605) );
  AND2X1 U13484 ( .IN1(P1_N3405), .IN2(n6886), .Q(n11607) );
  AND2X1 U13485 ( .IN1(P1_N4151), .IN2(n6881), .Q(n11608) );
  AND2X1 U13486 ( .IN1(P1_N3778), .IN2(n6886), .Q(n11609) );
  AND2X1 U13487 ( .IN1(P1_N4524), .IN2(n6921), .Q(n11610) );
  AND2X1 U13488 ( .IN1(n11612), .IN2(n6860), .Q(n11611) );
  AND2X1 U13489 ( .IN1(n11614), .IN2(n7458), .Q(n11613) );
  AND2X1 U13490 ( .IN1(n6621), .IN2(n11309), .Q(n11615) );
  AND2X1 U13491 ( .IN1(P1_N4787), .IN2(n6992), .Q(n11616) );
  AND2X1 U13492 ( .IN1(n11618), .IN2(n6954), .Q(n11617) );
  AND2X1 U13493 ( .IN1(n11620), .IN2(n7461), .Q(n11619) );
  AND2X1 U13494 ( .IN1(n11621), .IN2(n6984), .Q(n11315) );
  AND2X1 U13495 ( .IN1(n11622), .IN2(P1_N294), .Q(n11316) );
  AND2X1 U13496 ( .IN1(P1_N940), .IN2(n6886), .Q(n11623) );
  AND2X1 U13497 ( .IN1(P1_N1286), .IN2(n6921), .Q(n11624) );
  AND2X1 U13498 ( .IN1(P1_N1012), .IN2(n6886), .Q(n11625) );
  AND2X1 U13499 ( .IN1(P1_N1541), .IN2(n6881), .Q(n11626) );
  AND2X1 U13500 ( .IN1(n11628), .IN2(n6872), .Q(n11627) );
  AND2X1 U13501 ( .IN1(n11630), .IN2(n7458), .Q(n11629) );
  AND2X1 U13502 ( .IN1(P1_N1914), .IN2(n6922), .Q(n11631) );
  AND2X1 U13503 ( .IN1(P1_N2660), .IN2(n6921), .Q(n11632) );
  AND2X1 U13504 ( .IN1(P1_N2287), .IN2(n6922), .Q(n11633) );
  AND2X1 U13505 ( .IN1(P1_N3033), .IN2(n6921), .Q(n11634) );
  AND2X1 U13506 ( .IN1(n11636), .IN2(n6860), .Q(n11635) );
  AND2X1 U13507 ( .IN1(n11638), .IN2(n6871), .Q(n11637) );
  AND2X1 U13508 ( .IN1(n11640), .IN2(n6954), .Q(n11639) );
  AND2X1 U13509 ( .IN1(n11642), .IN2(n7461), .Q(n11641) );
  AND2X1 U13510 ( .IN1(P1_N3406), .IN2(n6886), .Q(n11643) );
  AND2X1 U13511 ( .IN1(P1_N4152), .IN2(n6921), .Q(n11644) );
  AND2X1 U13512 ( .IN1(P1_N3779), .IN2(n6886), .Q(n11645) );
  AND2X1 U13513 ( .IN1(P1_N4525), .IN2(n6921), .Q(n11646) );
  AND2X1 U13514 ( .IN1(n11648), .IN2(n6860), .Q(n11647) );
  OR2X1 U13329 ( .IN2(n11330), .IN1(n11329), .Q(P1_N4945) );
  OR2X1 U13330 ( .IN2(n11332), .IN1(n11331), .Q(P1_N4946) );
  OR2X1 U13331 ( .IN2(n11334), .IN1(n11333), .Q(P1_N4947) );
  OR2X1 U13332 ( .IN2(n11336), .IN1(n11335), .Q(P1_N4948) );
  OR2X1 U13333 ( .IN2(n11338), .IN1(n11337), .Q(P1_N4949) );
  OR2X1 U13334 ( .IN2(n11340), .IN1(n11339), .Q(P1_N4950) );
  OR2X1 U13335 ( .IN2(n11342), .IN1(n11341), .Q(P1_N4951) );
  OR2X1 U13336 ( .IN2(n11344), .IN1(n11343), .Q(P1_N4952) );
  OR2X1 U13337 ( .IN2(n11346), .IN1(n11345), .Q(P1_N4953) );
  OR2X1 U13338 ( .IN2(n11348), .IN1(n11347), .Q(P1_N4954) );
  OR2X1 U13339 ( .IN2(n11350), .IN1(n11349), .Q(P1_N4955) );
  OR2X1 U13340 ( .IN2(n11352), .IN1(n11351), .Q(P1_N4956) );
  OR2X1 U13341 ( .IN2(n11354), .IN1(n11353), .Q(P1_N4957) );
  OR2X1 U13342 ( .IN2(n11356), .IN1(n11355), .Q(P1_N4958) );
  OR2X1 U13343 ( .IN2(n11358), .IN1(n11357), .Q(P1_N4959) );
  OR2X1 U13344 ( .IN2(n11360), .IN1(n11359), .Q(P1_N4960) );
  OR2X1 U13345 ( .IN2(n11362), .IN1(n11361), .Q(P1_N4961) );
  OR2X1 U13346 ( .IN2(n11364), .IN1(n11363), .Q(P1_N4962) );
  OR2X1 U13347 ( .IN2(n11366), .IN1(n11365), .Q(P1_N4963) );
  OR2X1 U13348 ( .IN2(n11368), .IN1(n11367), .Q(P1_N4964) );
  OR2X1 U13349 ( .IN2(n11370), .IN1(n11369), .Q(P1_N4965) );
  OR2X1 U13350 ( .IN2(n11372), .IN1(n11371), .Q(P1_N4966) );
  OR2X1 U13351 ( .IN2(n11374), .IN1(n11373), .Q(P1_N4906) );
  OR2X1 U13352 ( .IN2(n11376), .IN1(n11375), .Q(P1_N4907) );
  OR2X1 U13353 ( .IN2(n11378), .IN1(n11377), .Q(P1_N4908) );
  OR2X1 U13354 ( .IN2(n11380), .IN1(n11379), .Q(P1_N4909) );
  OR2X1 U13355 ( .IN2(n11382), .IN1(n11381), .Q(P1_N4910) );
  OR2X1 U13356 ( .IN2(n11384), .IN1(n11383), .Q(P1_N4911) );
  OR2X1 U13357 ( .IN2(n11386), .IN1(n11385), .Q(P1_N4912) );
  OR2X1 U13358 ( .IN2(n11388), .IN1(n11387), .Q(P1_N4913) );
  OR2X1 U13359 ( .IN2(n11390), .IN1(n11389), .Q(P1_N4914) );
  OR2X1 U13360 ( .IN2(n11392), .IN1(n11391), .Q(P1_N4915) );
  OR2X1 U13361 ( .IN2(n11394), .IN1(n11393), .Q(P1_N4916) );
  OR2X1 U13362 ( .IN2(n11396), .IN1(n11395), .Q(P1_N4917) );
  OR2X1 U13363 ( .IN2(n11398), .IN1(n11397), .Q(P1_N4918) );
  OR2X1 U13364 ( .IN2(n11400), .IN1(n11399), .Q(P1_N4919) );
  OR2X1 U13365 ( .IN2(n11402), .IN1(n11401), .Q(P1_N4920) );
  OR2X1 U13366 ( .IN2(n11404), .IN1(n11403), .Q(P1_N4921) );
  OR2X1 U13367 ( .IN2(n11406), .IN1(n11405), .Q(P1_N4922) );
  OR2X1 U13368 ( .IN2(n11408), .IN1(n11407), .Q(P1_N4923) );
  OR2X1 U13369 ( .IN2(n11410), .IN1(n11409), .Q(P1_N4924) );
  OR2X1 U13370 ( .IN2(n11412), .IN1(n11411), .Q(P1_N4925) );
  OR2X1 U13371 ( .IN2(n11414), .IN1(n11413), .Q(P1_N4926) );
  OR2X1 U13372 ( .IN2(n11416), .IN1(n11415), .Q(P1_N4927) );
  OR2X1 U13373 ( .IN2(n11418), .IN1(n11417), .Q(P1_N4928) );
  OR2X1 U13374 ( .IN2(n11420), .IN1(n11419), .Q(P1_N4929) );
  OR2X1 U13375 ( .IN2(n11422), .IN1(n11421), .Q(P1_N4930) );
  OR2X1 U13376 ( .IN2(n11424), .IN1(n11423), .Q(P1_N4931) );
  OR2X1 U13377 ( .IN2(n11426), .IN1(n11425), .Q(P1_N4932) );
  OR2X1 U13378 ( .IN2(n11428), .IN1(n11427), .Q(P1_N4933) );
  OR2X1 U13379 ( .IN2(n11430), .IN1(n11429), .Q(P1_N4934) );
  OR2X1 U13380 ( .IN2(n11432), .IN1(n11431), .Q(P1_N4935) );
  OR2X1 U13381 ( .IN2(n11434), .IN1(n11433), .Q(P1_N4873) );
  OR2X1 U13382 ( .IN2(n11436), .IN1(n11435), .Q(P1_N4874) );
  OR2X1 U13383 ( .IN2(n11438), .IN1(n11437), .Q(P1_N4875) );
  OR2X1 U13384 ( .IN2(n11440), .IN1(n11439), .Q(P1_N4876) );
  OR2X1 U13385 ( .IN2(n11442), .IN1(n11441), .Q(P1_N4877) );
  OR2X1 U13386 ( .IN2(n11444), .IN1(n11443), .Q(P1_N4878) );
  OR2X1 U13387 ( .IN2(n11446), .IN1(n11445), .Q(P1_N4879) );
  OR2X1 U13388 ( .IN2(n11448), .IN1(n11447), .Q(P1_N4880) );
  OR2X1 U13389 ( .IN2(n11450), .IN1(n11449), .Q(P1_N4881) );
  OR2X1 U13390 ( .IN2(n11452), .IN1(n11451), .Q(P1_N4882) );
  OR2X1 U13391 ( .IN2(n11454), .IN1(n11453), .Q(P1_N4883) );
  OR2X1 U13392 ( .IN2(n11456), .IN1(n11455), .Q(P1_N4884) );
  OR2X1 U13393 ( .IN2(n11458), .IN1(n11457), .Q(P1_N4885) );
  OR2X1 U13394 ( .IN2(n11460), .IN1(n11459), .Q(P1_N4886) );
  OR2X1 U13395 ( .IN2(n11462), .IN1(n11461), .Q(P1_N4887) );
  OR2X1 U13396 ( .IN2(n11464), .IN1(n11463), .Q(P1_N4888) );
  OR2X1 U13397 ( .IN2(n11466), .IN1(n11465), .Q(P1_N4889) );
  OR2X1 U13398 ( .IN2(n11468), .IN1(n11467), .Q(P1_N4890) );
  OR2X1 U13399 ( .IN2(n11470), .IN1(n11469), .Q(P1_N4891) );
  OR2X1 U13400 ( .IN2(n11472), .IN1(n11471), .Q(P1_N4892) );
  OR2X1 U13401 ( .IN2(n11474), .IN1(n11473), .Q(P1_N4893) );
  OR2X1 U13402 ( .IN2(n11476), .IN1(n11475), .Q(P1_N4894) );
  OR2X1 U13403 ( .IN2(n11478), .IN1(n11477), .Q(P1_N4895) );
  OR2X1 U13404 ( .IN2(n11480), .IN1(n11479), .Q(P1_N4896) );
  OR2X1 U13405 ( .IN2(n11482), .IN1(n11481), .Q(P1_N4897) );
  OR2X1 U13406 ( .IN2(n11484), .IN1(n11483), .Q(P1_N4898) );
  OR2X1 U13407 ( .IN2(n11486), .IN1(n11485), .Q(P1_N4899) );
  OR2X1 U13408 ( .IN2(n11488), .IN1(n11487), .Q(P1_N4900) );
  OR2X1 U13409 ( .IN2(n11490), .IN1(n11489), .Q(P1_N4901) );
  OR2X1 U13410 ( .IN2(n11492), .IN1(n11491), .Q(P1_N4902) );
  AND2X1 U13411 ( .IN1(P1_N4786), .IN2(n6992), .Q(n11493) );
  OR2X1 U13412 ( .IN2(n11496), .IN1(n11495), .Q(P1_N4905) );
  AND2X1 U13413 ( .IN1(P1_N4817), .IN2(n6992), .Q(n11497) );
  AND2X1 U13414 ( .IN1(P1_N1570), .IN2(n6907), .Q(n11498) );
  OR2X1 U13415 ( .IN2(n11500), .IN1(n11499), .Q(P1_N4872) );
  AND2X1 U13416 ( .IN1(P1_N4816), .IN2(n6992), .Q(n11501) );
  AND2X1 U13417 ( .IN1(P1_N1569), .IN2(n6923), .Q(n11502) );
  OR2X1 U13418 ( .IN2(n11504), .IN1(n11503), .Q(P1_N4839) );
  OR2X1 U13419 ( .IN2(n11506), .IN1(n11505), .Q(P1_N4819) );
  OR2X1 U13420 ( .IN2(n11508), .IN1(n11507), .Q(P1_N4820) );
  OR2X1 U13421 ( .IN2(n11510), .IN1(n11509), .Q(P1_N4821) );
  OR2X1 U13319 ( .IN2(n6893), .IN1(n6869), .Q(n11309) );
  OR2X1 U13320 ( .IN2(n11312), .IN1(n11311), .Q(n11310) );
  OR2X1 U13321 ( .IN2(n11314), .IN1(n11313), .Q(P1_N5433) );
  OR2X1 U13322 ( .IN2(n11316), .IN1(n11315), .Q(P1_N4938) );
  OR2X1 U13323 ( .IN2(n11318), .IN1(n11317), .Q(P1_N4939) );
  OR2X1 U13324 ( .IN2(n11320), .IN1(n11319), .Q(P1_N4940) );
  OR2X1 U13325 ( .IN2(n11322), .IN1(n11321), .Q(P1_N4941) );
  OR2X1 U13326 ( .IN2(n11324), .IN1(n11323), .Q(P1_N4942) );
  OR2X1 U13327 ( .IN2(n11326), .IN1(n11325), .Q(P1_N4943) );
  OR2X1 U13328 ( .IN2(n11328), .IN1(n11327), .Q(P1_N4944) );
  INVX0 U12434 ( .ZN(n10368), .INP(n18348) );
  INVX0 U12435 ( .ZN(n10369), .INP(n10368) );
  INVX0 U12437 ( .ZN(n10372), .INP(n18698) );
  INVX0 U12438 ( .ZN(n10373), .INP(n10372) );
  INVX0 U12440 ( .ZN(n10376), .INP(n18318) );
  INVX0 U12441 ( .ZN(n10377), .INP(n10376) );
  INVX0 U12443 ( .ZN(n10380), .INP(n18666) );
  INVX0 U12444 ( .ZN(n10381), .INP(n10380) );
  INVX0 U12339 ( .ZN(n10249), .INP(n18190) );
  INVX0 U12340 ( .ZN(n10250), .INP(n18190) );
  INVX0 U12165 ( .ZN(n10022), .INP(n18706) );
  INVX0 U12166 ( .ZN(n10023), .INP(n10022) );
  INVX0 U12168 ( .ZN(n10026), .INP(n18708) );
  INVX0 U12169 ( .ZN(n10027), .INP(n10026) );
  INVX0 U12171 ( .ZN(n10030), .INP(n18710) );
  INVX0 U12172 ( .ZN(n10031), .INP(n10030) );
  INVX0 U12174 ( .ZN(n10034), .INP(n18712) );
  INVX0 U12175 ( .ZN(n10035), .INP(n10034) );
  INVX0 U12177 ( .ZN(n10038), .INP(n18714) );
  INVX0 U12178 ( .ZN(n10039), .INP(n10038) );
  INVX0 U12180 ( .ZN(n10042), .INP(n18716) );
  INVX0 U12181 ( .ZN(n10043), .INP(n10042) );
  INVX0 U12183 ( .ZN(n10046), .INP(n18718) );
  INVX0 U12184 ( .ZN(n10047), .INP(n10046) );
  INVX0 U12186 ( .ZN(n10050), .INP(n18720) );
  INVX0 U12187 ( .ZN(n10051), .INP(n10050) );
  INVX0 U12189 ( .ZN(n10054), .INP(n18722) );
  INVX0 U12190 ( .ZN(n10055), .INP(n10054) );
  INVX0 U12192 ( .ZN(n10058), .INP(n18724) );
  INVX0 U12193 ( .ZN(n10059), .INP(n10058) );
  INVX0 U12195 ( .ZN(n10062), .INP(n18726) );
  INVX0 U12196 ( .ZN(n10063), .INP(n10062) );
  INVX0 U12198 ( .ZN(n10066), .INP(n18728) );
  INVX0 U12199 ( .ZN(n10067), .INP(n10066) );
  INVX0 U12201 ( .ZN(n10070), .INP(n18730) );
  INVX0 U12202 ( .ZN(n10071), .INP(n10070) );
  INVX0 U12204 ( .ZN(n10074), .INP(n18732) );
  INVX0 U12205 ( .ZN(n10075), .INP(n10074) );
  INVX0 U12207 ( .ZN(n10078), .INP(n18734) );
  INVX0 U12208 ( .ZN(n10079), .INP(n10078) );
  INVX0 U12210 ( .ZN(n10082), .INP(n18736) );
  INVX0 U12211 ( .ZN(n10083), .INP(n10082) );
  INVX0 U12213 ( .ZN(n10086), .INP(n18738) );
  INVX0 U12214 ( .ZN(n10087), .INP(n10086) );
  INVX0 U12216 ( .ZN(n10090), .INP(n18740) );
  INVX0 U12217 ( .ZN(n10091), .INP(n10090) );
  INVX0 U12219 ( .ZN(n10094), .INP(n19006) );
  INVX0 U12220 ( .ZN(n10095), .INP(n10094) );
  INVX0 U12222 ( .ZN(n10098), .INP(n19018) );
  INVX0 U12223 ( .ZN(n10099), .INP(n10098) );
  INVX0 U12226 ( .ZN(n10103), .INP(n18192) );
  INVX0 U12229 ( .ZN(n10107), .INP(n18193) );
  INVX0 U12231 ( .ZN(n10110), .INP(n18904) );
  INVX0 U12232 ( .ZN(n10111), .INP(n10110) );
  INVX0 U12233 ( .ZN(n10112), .INP(n10110) );
  INVX0 U12236 ( .ZN(n10116), .INP(n18191) );
  INVX0 U12237 ( .ZN(n10117), .INP(n18191) );
  INVX0 U12242 ( .ZN(n10124), .INP(n18696) );
  INVX0 U12243 ( .ZN(n10125), .INP(n10124) );
  INVX0 U12245 ( .ZN(n10128), .INP(n18700) );
  INVX0 U12246 ( .ZN(n10129), .INP(n10128) );
  INVX0 U12248 ( .ZN(n10132), .INP(n19004) );
  INVX0 U12249 ( .ZN(n10133), .INP(n10132) );
  INVX0 U12251 ( .ZN(n10136), .INP(n19020) );
  INVX0 U12252 ( .ZN(n10137), .INP(n10136) );
  INVX0 U12254 ( .ZN(n10140), .INP(n18350) );
  INVX0 U12255 ( .ZN(n10141), .INP(n10140) );
  INVX0 U12257 ( .ZN(n10144), .INP(n18702) );
  INVX0 U12258 ( .ZN(n10145), .INP(n10144) );
  INVX0 U12286 ( .ZN(n10182), .INP(n18320) );
  INVX0 U12287 ( .ZN(n10183), .INP(n10182) );
  INVX0 U12289 ( .ZN(n10186), .INP(n18668) );
  INVX0 U12290 ( .ZN(n10187), .INP(n10186) );
  INVX0 U12292 ( .ZN(n10190), .INP(n18316) );
  INVX0 U12293 ( .ZN(n10191), .INP(n10190) );
  INVX0 U12295 ( .ZN(n10194), .INP(n18664) );
  INVX0 U12296 ( .ZN(n10195), .INP(n10194) );
  INVX0 U12026 ( .ZN(n9837), .INP(n9836) );
  INVX0 U12027 ( .ZN(n9838), .INP(n9836) );
  INVX0 U12029 ( .ZN(n9841), .INP(n18998) );
  INVX0 U12030 ( .ZN(n9842), .INP(n9841) );
  INVX0 U12031 ( .ZN(n9843), .INP(n9841) );
  INVX0 U12036 ( .ZN(n9850), .INP(n18390) );
  INVX0 U12037 ( .ZN(n9851), .INP(n9850) );
  INVX0 U12039 ( .ZN(n9854), .INP(n18398) );
  INVX0 U12040 ( .ZN(n9855), .INP(n9854) );
  INVX0 U12042 ( .ZN(n9858), .INP(n18406) );
  INVX0 U12043 ( .ZN(n9859), .INP(n9858) );
  INVX0 U12045 ( .ZN(n9862), .INP(n18414) );
  INVX0 U12046 ( .ZN(n9863), .INP(n9862) );
  INVX0 U12048 ( .ZN(n9866), .INP(n18422) );
  INVX0 U12049 ( .ZN(n9867), .INP(n9866) );
  INVX0 U12051 ( .ZN(n9870), .INP(n18428) );
  INVX0 U12052 ( .ZN(n9871), .INP(n9870) );
  INVX0 U12054 ( .ZN(n9874), .INP(n18432) );
  INVX0 U12055 ( .ZN(n9875), .INP(n9874) );
  INVX0 U12057 ( .ZN(n9878), .INP(n18436) );
  INVX0 U12058 ( .ZN(n9879), .INP(n9878) );
  INVX0 U12060 ( .ZN(n9882), .INP(n18440) );
  INVX0 U12061 ( .ZN(n9883), .INP(n9882) );
  INVX0 U12063 ( .ZN(n9886), .INP(n18444) );
  INVX0 U12064 ( .ZN(n9887), .INP(n9886) );
  INVX0 U12066 ( .ZN(n9890), .INP(n18448) );
  INVX0 U12067 ( .ZN(n9891), .INP(n9890) );
  INVX0 U12069 ( .ZN(n9894), .INP(n18452) );
  INVX0 U12070 ( .ZN(n9895), .INP(n9894) );
  INVX0 U12072 ( .ZN(n9898), .INP(n18456) );
  INVX0 U12073 ( .ZN(n9899), .INP(n9898) );
  INVX0 U12075 ( .ZN(n9902), .INP(n18742) );
  INVX0 U12076 ( .ZN(n9903), .INP(n9902) );
  INVX0 U12078 ( .ZN(n9906), .INP(n18744) );
  INVX0 U12079 ( .ZN(n9907), .INP(n9906) );
  INVX0 U12081 ( .ZN(n9910), .INP(n18746) );
  INVX0 U12082 ( .ZN(n9911), .INP(n9910) );
  INVX0 U12084 ( .ZN(n9914), .INP(n18748) );
  INVX0 U12085 ( .ZN(n9915), .INP(n9914) );
  INVX0 U12087 ( .ZN(n9918), .INP(n18750) );
  INVX0 U12088 ( .ZN(n9919), .INP(n9918) );
  INVX0 U12090 ( .ZN(n9922), .INP(n18752) );
  INVX0 U12091 ( .ZN(n9923), .INP(n9922) );
  INVX0 U12093 ( .ZN(n9926), .INP(n18754) );
  INVX0 U12094 ( .ZN(n9927), .INP(n9926) );
  INVX0 U12096 ( .ZN(n9930), .INP(n18756) );
  INVX0 U12097 ( .ZN(n9931), .INP(n9930) );
  INVX0 U12099 ( .ZN(n9934), .INP(n18352) );
  INVX0 U12100 ( .ZN(n9935), .INP(n9934) );
  INVX0 U12102 ( .ZN(n9938), .INP(n18356) );
  INVX0 U12103 ( .ZN(n9939), .INP(n9938) );
  INVX0 U12105 ( .ZN(n9942), .INP(n18360) );
  INVX0 U12106 ( .ZN(n9943), .INP(n9942) );
  INVX0 U12108 ( .ZN(n9946), .INP(n18364) );
  INVX0 U12109 ( .ZN(n9947), .INP(n9946) );
  INVX0 U12111 ( .ZN(n9950), .INP(n18368) );
  INVX0 U12112 ( .ZN(n9951), .INP(n9950) );
  INVX0 U12114 ( .ZN(n9954), .INP(n18372) );
  INVX0 U12115 ( .ZN(n9955), .INP(n9954) );
  INVX0 U12117 ( .ZN(n9958), .INP(n18376) );
  INVX0 U12118 ( .ZN(n9959), .INP(n9958) );
  INVX0 U12120 ( .ZN(n9962), .INP(n18380) );
  INVX0 U12121 ( .ZN(n9963), .INP(n9962) );
  INVX0 U12123 ( .ZN(n9966), .INP(n18384) );
  INVX0 U12124 ( .ZN(n9967), .INP(n9966) );
  INVX0 U12126 ( .ZN(n9970), .INP(n18388) );
  INVX0 U12127 ( .ZN(n9971), .INP(n9970) );
  INVX0 U12129 ( .ZN(n9974), .INP(n18392) );
  INVX0 U12130 ( .ZN(n9975), .INP(n9974) );
  INVX0 U12132 ( .ZN(n9978), .INP(n18396) );
  INVX0 U12133 ( .ZN(n9979), .INP(n9978) );
  INVX0 U12135 ( .ZN(n9982), .INP(n18400) );
  INVX0 U12136 ( .ZN(n9983), .INP(n9982) );
  INVX0 U12138 ( .ZN(n9986), .INP(n18404) );
  INVX0 U12139 ( .ZN(n9987), .INP(n9986) );
  INVX0 U12141 ( .ZN(n9990), .INP(n18408) );
  INVX0 U12142 ( .ZN(n9991), .INP(n9990) );
  INVX0 U12144 ( .ZN(n9994), .INP(n18412) );
  INVX0 U12145 ( .ZN(n9995), .INP(n9994) );
  INVX0 U12147 ( .ZN(n9998), .INP(n18416) );
  INVX0 U12148 ( .ZN(n9999), .INP(n9998) );
  INVX0 U12150 ( .ZN(n10002), .INP(n18420) );
  INVX0 U12151 ( .ZN(n10003), .INP(n10002) );
  INVX0 U12153 ( .ZN(n10006), .INP(n18424) );
  INVX0 U12154 ( .ZN(n10007), .INP(n10006) );
  INVX0 U12156 ( .ZN(n10010), .INP(n18430) );
  INVX0 U12157 ( .ZN(n10011), .INP(n10010) );
  INVX0 U12159 ( .ZN(n10014), .INP(n18438) );
  INVX0 U12160 ( .ZN(n10015), .INP(n10014) );
  INVX0 U12162 ( .ZN(n10018), .INP(n18704) );
  INVX0 U12163 ( .ZN(n10019), .INP(n10018) );
  INVX0 U11885 ( .ZN(n9649), .INP(n9648) );
  INVX0 U11890 ( .ZN(n9656), .INP(n18446) );
  INVX0 U11891 ( .ZN(n9657), .INP(n9656) );
  INVX0 U11893 ( .ZN(n9660), .INP(n18386) );
  INVX0 U11894 ( .ZN(n9661), .INP(n9660) );
  INVX0 U11896 ( .ZN(n9664), .INP(n18394) );
  INVX0 U11897 ( .ZN(n9665), .INP(n9664) );
  INVX0 U11899 ( .ZN(n9668), .INP(n18402) );
  INVX0 U11900 ( .ZN(n9669), .INP(n9668) );
  INVX0 U11902 ( .ZN(n9672), .INP(n18410) );
  INVX0 U11903 ( .ZN(n9673), .INP(n9672) );
  INVX0 U11905 ( .ZN(n9676), .INP(n18418) );
  INVX0 U11906 ( .ZN(n9677), .INP(n9676) );
  INVX0 U11908 ( .ZN(n9680), .INP(n18426) );
  INVX0 U11909 ( .ZN(n9681), .INP(n9680) );
  INVX0 U11911 ( .ZN(n9684), .INP(n18434) );
  INVX0 U11912 ( .ZN(n9685), .INP(n9684) );
  INVX0 U11914 ( .ZN(n9688), .INP(n18442) );
  INVX0 U11915 ( .ZN(n9689), .INP(n9688) );
  INVX0 U11917 ( .ZN(n9692), .INP(n18552) );
  INVX0 U11918 ( .ZN(n9693), .INP(n9692) );
  INVX0 U11920 ( .ZN(n9696), .INP(n18554) );
  INVX0 U11921 ( .ZN(n9697), .INP(n9696) );
  INVX0 U11923 ( .ZN(n9700), .INP(n18556) );
  INVX0 U11924 ( .ZN(n9701), .INP(n9700) );
  INVX0 U11926 ( .ZN(n9704), .INP(n18558) );
  INVX0 U11927 ( .ZN(n9705), .INP(n9704) );
  INVX0 U11929 ( .ZN(n9708), .INP(n18560) );
  INVX0 U11930 ( .ZN(n9709), .INP(n9708) );
  INVX0 U11932 ( .ZN(n9712), .INP(n18562) );
  INVX0 U11933 ( .ZN(n9713), .INP(n9712) );
  INVX0 U11935 ( .ZN(n9716), .INP(n18564) );
  INVX0 U11936 ( .ZN(n9717), .INP(n9716) );
  INVX0 U11938 ( .ZN(n9720), .INP(n18566) );
  INVX0 U11939 ( .ZN(n9721), .INP(n9720) );
  INVX0 U11941 ( .ZN(n9724), .INP(n18568) );
  INVX0 U11942 ( .ZN(n9725), .INP(n9724) );
  INVX0 U11944 ( .ZN(n9728), .INP(n18570) );
  INVX0 U11945 ( .ZN(n9729), .INP(n9728) );
  INVX0 U11948 ( .ZN(n9733), .INP(n18187) );
  INVX0 U11950 ( .ZN(n9736), .INP(n18572) );
  INVX0 U11951 ( .ZN(n9737), .INP(n9736) );
  INVX0 U11953 ( .ZN(n9740), .INP(n18574) );
  INVX0 U11954 ( .ZN(n9741), .INP(n9740) );
  INVX0 U11956 ( .ZN(n9744), .INP(n18576) );
  INVX0 U11957 ( .ZN(n9745), .INP(n9744) );
  INVX0 U11959 ( .ZN(n9748), .INP(n18578) );
  INVX0 U11960 ( .ZN(n9749), .INP(n9748) );
  INVX0 U11962 ( .ZN(n9752), .INP(n18580) );
  INVX0 U11963 ( .ZN(n9753), .INP(n9752) );
  INVX0 U11965 ( .ZN(n9756), .INP(n18582) );
  INVX0 U11966 ( .ZN(n9757), .INP(n9756) );
  INVX0 U11968 ( .ZN(n9760), .INP(n18584) );
  INVX0 U11969 ( .ZN(n9761), .INP(n9760) );
  INVX0 U11971 ( .ZN(n9764), .INP(n18606) );
  INVX0 U11972 ( .ZN(n9765), .INP(n9764) );
  INVX0 U11974 ( .ZN(n9768), .INP(n18608) );
  INVX0 U11975 ( .ZN(n9769), .INP(n9768) );
  INVX0 U11977 ( .ZN(n9772), .INP(n18610) );
  INVX0 U11978 ( .ZN(n9773), .INP(n9772) );
  INVX0 U11980 ( .ZN(n9776), .INP(n18612) );
  INVX0 U11981 ( .ZN(n9777), .INP(n9776) );
  INVX0 U11983 ( .ZN(n9780), .INP(n18614) );
  INVX0 U11984 ( .ZN(n9781), .INP(n9780) );
  INVX0 U11986 ( .ZN(n9784), .INP(n18616) );
  INVX0 U11987 ( .ZN(n9785), .INP(n9784) );
  INVX0 U11989 ( .ZN(n9788), .INP(n18618) );
  INVX0 U11990 ( .ZN(n9789), .INP(n9788) );
  INVX0 U11992 ( .ZN(n9792), .INP(n18620) );
  INVX0 U11993 ( .ZN(n9793), .INP(n9792) );
  INVX0 U11995 ( .ZN(n9796), .INP(n18622) );
  INVX0 U11996 ( .ZN(n9797), .INP(n9796) );
  INVX0 U11998 ( .ZN(n9800), .INP(n18624) );
  INVX0 U11999 ( .ZN(n9801), .INP(n9800) );
  INVX0 U12001 ( .ZN(n9804), .INP(n18626) );
  INVX0 U12002 ( .ZN(n9805), .INP(n9804) );
  INVX0 U12004 ( .ZN(n9808), .INP(n18628) );
  INVX0 U12005 ( .ZN(n9809), .INP(n9808) );
  INVX0 U12007 ( .ZN(n9812), .INP(n18630) );
  INVX0 U12008 ( .ZN(n9813), .INP(n9812) );
  INVX0 U12010 ( .ZN(n9816), .INP(n18632) );
  INVX0 U12011 ( .ZN(n9817), .INP(n9816) );
  INVX0 U12013 ( .ZN(n9820), .INP(n18634) );
  INVX0 U12014 ( .ZN(n9821), .INP(n9820) );
  INVX0 U12016 ( .ZN(n9824), .INP(n18636) );
  INVX0 U12017 ( .ZN(n9825), .INP(n9824) );
  INVX0 U12019 ( .ZN(n9828), .INP(n18638) );
  INVX0 U12020 ( .ZN(n9829), .INP(n9828) );
  INVX0 U12022 ( .ZN(n9832), .INP(n18640) );
  INVX0 U12023 ( .ZN(n9833), .INP(n9832) );
  INVX0 U12025 ( .ZN(n9836), .INP(n18940) );
  INVX0 U11745 ( .ZN(n9464), .INP(n18233) );
  INVX0 U11746 ( .ZN(n9465), .INP(n9464) );
  INVX0 U11748 ( .ZN(n9468), .INP(n18235) );
  INVX0 U11749 ( .ZN(n9469), .INP(n9468) );
  INVX0 U11751 ( .ZN(n9472), .INP(n18237) );
  INVX0 U11752 ( .ZN(n9473), .INP(n9472) );
  INVX0 U11754 ( .ZN(n9476), .INP(n18239) );
  INVX0 U11755 ( .ZN(n9477), .INP(n9476) );
  INVX0 U11757 ( .ZN(n9480), .INP(n18241) );
  INVX0 U11758 ( .ZN(n9481), .INP(n9480) );
  INVX0 U11760 ( .ZN(n9484), .INP(n18243) );
  INVX0 U11761 ( .ZN(n9485), .INP(n9484) );
  INVX0 U11763 ( .ZN(n9488), .INP(n19002) );
  INVX0 U11764 ( .ZN(n9489), .INP(n9488) );
  INVX0 U11766 ( .ZN(n9492), .INP(n18550) );
  INVX0 U11767 ( .ZN(n9493), .INP(n9492) );
  INVX0 U11770 ( .ZN(n9497), .INP(n18188) );
  INVX0 U11772 ( .ZN(n9500), .INP(n18780) );
  INVX0 U11773 ( .ZN(n9501), .INP(n9500) );
  INVX0 U11775 ( .ZN(n9504), .INP(n18782) );
  INVX0 U11776 ( .ZN(n9505), .INP(n9504) );
  INVX0 U11778 ( .ZN(n9508), .INP(n18784) );
  INVX0 U11779 ( .ZN(n9509), .INP(n9508) );
  INVX0 U11781 ( .ZN(n9512), .INP(n18786) );
  INVX0 U11782 ( .ZN(n9513), .INP(n9512) );
  INVX0 U11784 ( .ZN(n9516), .INP(n18788) );
  INVX0 U11785 ( .ZN(n9517), .INP(n9516) );
  INVX0 U11787 ( .ZN(n9520), .INP(n18790) );
  INVX0 U11788 ( .ZN(n9521), .INP(n9520) );
  INVX0 U11790 ( .ZN(n9524), .INP(n18792) );
  INVX0 U11791 ( .ZN(n9525), .INP(n9524) );
  INVX0 U11793 ( .ZN(n9528), .INP(n18794) );
  INVX0 U11794 ( .ZN(n9529), .INP(n9528) );
  INVX0 U11796 ( .ZN(n9532), .INP(n18796) );
  INVX0 U11797 ( .ZN(n9533), .INP(n9532) );
  INVX0 U11799 ( .ZN(n9536), .INP(n18798) );
  INVX0 U11800 ( .ZN(n9537), .INP(n9536) );
  INVX0 U11802 ( .ZN(n9540), .INP(n18800) );
  INVX0 U11803 ( .ZN(n9541), .INP(n9540) );
  INVX0 U11805 ( .ZN(n9544), .INP(n18802) );
  INVX0 U11806 ( .ZN(n9545), .INP(n9544) );
  INVX0 U11808 ( .ZN(n9548), .INP(n18804) );
  INVX0 U11809 ( .ZN(n9549), .INP(n9548) );
  INVX0 U11811 ( .ZN(n9552), .INP(n18806) );
  INVX0 U11812 ( .ZN(n9553), .INP(n9552) );
  INVX0 U11814 ( .ZN(n9556), .INP(n18808) );
  INVX0 U11815 ( .ZN(n9557), .INP(n9556) );
  INVX0 U11821 ( .ZN(n9564), .INP(n18247) );
  INVX0 U11822 ( .ZN(n9565), .INP(n9564) );
  INVX0 U11824 ( .ZN(n9568), .INP(n18249) );
  INVX0 U11825 ( .ZN(n9569), .INP(n9568) );
  INVX0 U11827 ( .ZN(n9572), .INP(n18251) );
  INVX0 U11828 ( .ZN(n9573), .INP(n9572) );
  INVX0 U11830 ( .ZN(n9576), .INP(n18253) );
  INVX0 U11831 ( .ZN(n9577), .INP(n9576) );
  INVX0 U11833 ( .ZN(n9580), .INP(n18255) );
  INVX0 U11834 ( .ZN(n9581), .INP(n9580) );
  INVX0 U11836 ( .ZN(n9584), .INP(n18257) );
  INVX0 U11837 ( .ZN(n9585), .INP(n9584) );
  INVX0 U11839 ( .ZN(n9588), .INP(n18259) );
  INVX0 U11840 ( .ZN(n9589), .INP(n9588) );
  INVX0 U11842 ( .ZN(n9592), .INP(n18261) );
  INVX0 U11843 ( .ZN(n9593), .INP(n9592) );
  INVX0 U11845 ( .ZN(n9596), .INP(n18263) );
  INVX0 U11846 ( .ZN(n9597), .INP(n9596) );
  INVX0 U11849 ( .ZN(n9601), .INP(n18186) );
  INVX0 U11851 ( .ZN(n9604), .INP(n18265) );
  INVX0 U11852 ( .ZN(n9605), .INP(n9604) );
  INVX0 U11854 ( .ZN(n9608), .INP(n18267) );
  INVX0 U11855 ( .ZN(n9609), .INP(n9608) );
  INVX0 U11857 ( .ZN(n9612), .INP(n18269) );
  INVX0 U11858 ( .ZN(n9613), .INP(n9612) );
  INVX0 U11860 ( .ZN(n9616), .INP(n18271) );
  INVX0 U11861 ( .ZN(n9617), .INP(n9616) );
  INVX0 U11863 ( .ZN(n9620), .INP(n18273) );
  INVX0 U11864 ( .ZN(n9621), .INP(n9620) );
  INVX0 U11866 ( .ZN(n9624), .INP(n18275) );
  INVX0 U11867 ( .ZN(n9625), .INP(n9624) );
  INVX0 U11869 ( .ZN(n9628), .INP(n18277) );
  INVX0 U11870 ( .ZN(n9629), .INP(n9628) );
  INVX0 U11872 ( .ZN(n9632), .INP(n18293) );
  INVX0 U11873 ( .ZN(n9633), .INP(n9632) );
  INVX0 U11875 ( .ZN(n9636), .INP(n18358) );
  INVX0 U11876 ( .ZN(n9637), .INP(n9636) );
  INVX0 U11878 ( .ZN(n9640), .INP(n18366) );
  INVX0 U11879 ( .ZN(n9641), .INP(n9640) );
  INVX0 U11881 ( .ZN(n9644), .INP(n18374) );
  INVX0 U11882 ( .ZN(n9645), .INP(n9644) );
  INVX0 U11884 ( .ZN(n9648), .INP(n18382) );
  INVX0 U11604 ( .ZN(n9277), .INP(n18948) );
  INVX0 U11605 ( .ZN(n9278), .INP(n9277) );
  INVX0 U11607 ( .ZN(n9281), .INP(n18950) );
  INVX0 U11608 ( .ZN(n9282), .INP(n9281) );
  INVX0 U11610 ( .ZN(n9285), .INP(n18952) );
  INVX0 U11611 ( .ZN(n9286), .INP(n9285) );
  INVX0 U11613 ( .ZN(n9289), .INP(n18954) );
  INVX0 U11614 ( .ZN(n9290), .INP(n9289) );
  INVX0 U11616 ( .ZN(n9293), .INP(n18956) );
  INVX0 U11617 ( .ZN(n9294), .INP(n9293) );
  INVX0 U11619 ( .ZN(n9297), .INP(n18958) );
  INVX0 U11620 ( .ZN(n9298), .INP(n9297) );
  INVX0 U11622 ( .ZN(n9301), .INP(n18960) );
  INVX0 U11623 ( .ZN(n9302), .INP(n9301) );
  INVX0 U11625 ( .ZN(n9305), .INP(n19012) );
  INVX0 U11626 ( .ZN(n9306), .INP(n9305) );
  INVX0 U11628 ( .ZN(n9309), .INP(n19016) );
  INVX0 U11629 ( .ZN(n9310), .INP(n9309) );
  INVX0 U11631 ( .ZN(n9313), .INP(n19022) );
  INVX0 U11632 ( .ZN(n9314), .INP(n9313) );
  INVX0 U11634 ( .ZN(n9317), .INP(n18279) );
  INVX0 U11635 ( .ZN(n9318), .INP(n9317) );
  INVX0 U11637 ( .ZN(n9321), .INP(n18283) );
  INVX0 U11638 ( .ZN(n9322), .INP(n9321) );
  INVX0 U11641 ( .ZN(n9325), .INP(n18183) );
  INVX0 U11643 ( .ZN(n9328), .INP(n18281) );
  INVX0 U11644 ( .ZN(n9329), .INP(n9328) );
  INVX0 U11646 ( .ZN(n9332), .INP(n18460) );
  INVX0 U11647 ( .ZN(n9333), .INP(n9332) );
  INVX0 U11649 ( .ZN(n9336), .INP(n18758) );
  INVX0 U11650 ( .ZN(n9337), .INP(n9336) );
  INVX0 U11652 ( .ZN(n9340), .INP(n19010) );
  INVX0 U11653 ( .ZN(n9341), .INP(n9340) );
  INVX0 U11655 ( .ZN(n9344), .INP(n19014) );
  INVX0 U11656 ( .ZN(n9345), .INP(n9344) );
  INVX0 U11658 ( .ZN(n9348), .INP(n18762) );
  INVX0 U11659 ( .ZN(n9349), .INP(n9348) );
  INVX0 U11661 ( .ZN(n9352), .INP(n18764) );
  INVX0 U11662 ( .ZN(n9353), .INP(n9352) );
  INVX0 U11664 ( .ZN(n9356), .INP(n18766) );
  INVX0 U11665 ( .ZN(n9357), .INP(n9356) );
  INVX0 U11667 ( .ZN(n9360), .INP(n18768) );
  INVX0 U11668 ( .ZN(n9361), .INP(n9360) );
  INVX0 U11670 ( .ZN(n9364), .INP(n18770) );
  INVX0 U11671 ( .ZN(n9365), .INP(n9364) );
  INVX0 U11673 ( .ZN(n9368), .INP(n18772) );
  INVX0 U11674 ( .ZN(n9369), .INP(n9368) );
  INVX0 U11676 ( .ZN(n9372), .INP(n18774) );
  INVX0 U11677 ( .ZN(n9373), .INP(n9372) );
  INVX0 U11679 ( .ZN(n9376), .INP(n18776) );
  INVX0 U11680 ( .ZN(n9377), .INP(n9376) );
  INVX0 U11682 ( .ZN(n9380), .INP(n18778) );
  INVX0 U11683 ( .ZN(n9381), .INP(n9380) );
  INVX0 U11685 ( .ZN(n9384), .INP(n18462) );
  INVX0 U11686 ( .ZN(n9385), .INP(n9384) );
  INVX0 U11688 ( .ZN(n9388), .INP(n18760) );
  INVX0 U11689 ( .ZN(n9389), .INP(n9388) );
  INVX0 U11694 ( .ZN(n9396), .INP(n18810) );
  INVX0 U11695 ( .ZN(n9397), .INP(n9396) );
  INVX0 U11697 ( .ZN(n9400), .INP(n18354) );
  INVX0 U11698 ( .ZN(n9401), .INP(n9400) );
  INVX0 U11700 ( .ZN(n9404), .INP(n18362) );
  INVX0 U11701 ( .ZN(n9405), .INP(n9404) );
  INVX0 U11703 ( .ZN(n9408), .INP(n18370) );
  INVX0 U11704 ( .ZN(n9409), .INP(n9408) );
  INVX0 U11706 ( .ZN(n9412), .INP(n18378) );
  INVX0 U11707 ( .ZN(n9413), .INP(n9412) );
  INVX0 U11709 ( .ZN(n9416), .INP(n18211) );
  INVX0 U11710 ( .ZN(n9417), .INP(n9416) );
  INVX0 U11712 ( .ZN(n9420), .INP(n18213) );
  INVX0 U11713 ( .ZN(n9421), .INP(n9420) );
  INVX0 U11715 ( .ZN(n9424), .INP(n18215) );
  INVX0 U11716 ( .ZN(n9425), .INP(n9424) );
  INVX0 U11718 ( .ZN(n9428), .INP(n18217) );
  INVX0 U11719 ( .ZN(n9429), .INP(n9428) );
  INVX0 U11721 ( .ZN(n9432), .INP(n18219) );
  INVX0 U11722 ( .ZN(n9433), .INP(n9432) );
  INVX0 U11724 ( .ZN(n9436), .INP(n18221) );
  INVX0 U11725 ( .ZN(n9437), .INP(n9436) );
  INVX0 U11727 ( .ZN(n9440), .INP(n18223) );
  INVX0 U11728 ( .ZN(n9441), .INP(n9440) );
  INVX0 U11730 ( .ZN(n9444), .INP(n18225) );
  INVX0 U11731 ( .ZN(n9445), .INP(n9444) );
  INVX0 U11733 ( .ZN(n9448), .INP(n18227) );
  INVX0 U11734 ( .ZN(n9449), .INP(n9448) );
  INVX0 U11737 ( .ZN(n9453), .INP(n18185) );
  INVX0 U11739 ( .ZN(n9456), .INP(n18229) );
  INVX0 U11740 ( .ZN(n9457), .INP(n9456) );
  INVX0 U11742 ( .ZN(n9460), .INP(n18231) );
  INVX0 U11743 ( .ZN(n9461), .INP(n9460) );
  INVX0 U11464 ( .ZN(n9090), .INP(n9089) );
  INVX0 U11466 ( .ZN(n9093), .INP(n18604) );
  INVX0 U11467 ( .ZN(n9094), .INP(n9093) );
  INVX0 U11469 ( .ZN(n9097), .INP(n18820) );
  INVX0 U11470 ( .ZN(n9098), .INP(n9097) );
  INVX0 U11472 ( .ZN(n9101), .INP(n18822) );
  INVX0 U11473 ( .ZN(n9102), .INP(n9101) );
  INVX0 U11475 ( .ZN(n9105), .INP(n18824) );
  INVX0 U11476 ( .ZN(n9106), .INP(n9105) );
  INVX0 U11478 ( .ZN(n9109), .INP(n18826) );
  INVX0 U11479 ( .ZN(n9110), .INP(n9109) );
  INVX0 U11481 ( .ZN(n9113), .INP(n18828) );
  INVX0 U11482 ( .ZN(n9114), .INP(n9113) );
  INVX0 U11484 ( .ZN(n9117), .INP(n18830) );
  INVX0 U11485 ( .ZN(n9118), .INP(n9117) );
  INVX0 U11487 ( .ZN(n9121), .INP(n18832) );
  INVX0 U11488 ( .ZN(n9122), .INP(n9121) );
  INVX0 U11490 ( .ZN(n9125), .INP(n18834) );
  INVX0 U11491 ( .ZN(n9126), .INP(n9125) );
  INVX0 U11493 ( .ZN(n9129), .INP(n18836) );
  INVX0 U11494 ( .ZN(n9130), .INP(n9129) );
  INVX0 U11496 ( .ZN(n9133), .INP(n18838) );
  INVX0 U11497 ( .ZN(n9134), .INP(n9133) );
  INVX0 U11499 ( .ZN(n9137), .INP(n18840) );
  INVX0 U11500 ( .ZN(n9138), .INP(n9137) );
  INVX0 U11502 ( .ZN(n9141), .INP(n18842) );
  INVX0 U11503 ( .ZN(n9142), .INP(n9141) );
  INVX0 U11505 ( .ZN(n9145), .INP(n18844) );
  INVX0 U11506 ( .ZN(n9146), .INP(n9145) );
  INVX0 U11508 ( .ZN(n9149), .INP(n18846) );
  INVX0 U11509 ( .ZN(n9150), .INP(n9149) );
  INVX0 U11511 ( .ZN(n9153), .INP(n18848) );
  INVX0 U11512 ( .ZN(n9154), .INP(n9153) );
  INVX0 U11514 ( .ZN(n9157), .INP(n18850) );
  INVX0 U11515 ( .ZN(n9158), .INP(n9157) );
  INVX0 U11517 ( .ZN(n9161), .INP(n18852) );
  INVX0 U11518 ( .ZN(n9162), .INP(n9161) );
  INVX0 U11520 ( .ZN(n9165), .INP(n18854) );
  INVX0 U11521 ( .ZN(n9166), .INP(n9165) );
  INVX0 U11523 ( .ZN(n9169), .INP(n18856) );
  INVX0 U11524 ( .ZN(n9170), .INP(n9169) );
  INVX0 U11526 ( .ZN(n9173), .INP(n18858) );
  INVX0 U11527 ( .ZN(n9174), .INP(n9173) );
  INVX0 U11529 ( .ZN(n9177), .INP(n18860) );
  INVX0 U11530 ( .ZN(n9178), .INP(n9177) );
  INVX0 U11532 ( .ZN(n9181), .INP(n18862) );
  INVX0 U11533 ( .ZN(n9182), .INP(n9181) );
  INVX0 U11535 ( .ZN(n9185), .INP(n18864) );
  INVX0 U11536 ( .ZN(n9186), .INP(n9185) );
  INVX0 U11538 ( .ZN(n9189), .INP(n18866) );
  INVX0 U11539 ( .ZN(n9190), .INP(n9189) );
  INVX0 U11541 ( .ZN(n9193), .INP(n18868) );
  INVX0 U11542 ( .ZN(n9194), .INP(n9193) );
  INVX0 U11544 ( .ZN(n9197), .INP(n18870) );
  INVX0 U11545 ( .ZN(n9198), .INP(n9197) );
  INVX0 U11547 ( .ZN(n9201), .INP(n18872) );
  INVX0 U11548 ( .ZN(n9202), .INP(n9201) );
  INVX0 U11550 ( .ZN(n9205), .INP(n18874) );
  INVX0 U11551 ( .ZN(n9206), .INP(n9205) );
  INVX0 U11553 ( .ZN(n9209), .INP(n18876) );
  INVX0 U11554 ( .ZN(n9210), .INP(n9209) );
  INVX0 U11556 ( .ZN(n9213), .INP(n18878) );
  INVX0 U11557 ( .ZN(n9214), .INP(n9213) );
  INVX0 U11559 ( .ZN(n9217), .INP(n18880) );
  INVX0 U11560 ( .ZN(n9218), .INP(n9217) );
  INVX0 U11562 ( .ZN(n9221), .INP(n18882) );
  INVX0 U11563 ( .ZN(n9222), .INP(n9221) );
  INVX0 U11565 ( .ZN(n9225), .INP(n18884) );
  INVX0 U11566 ( .ZN(n9226), .INP(n9225) );
  INVX0 U11568 ( .ZN(n9229), .INP(n18886) );
  INVX0 U11569 ( .ZN(n9230), .INP(n9229) );
  INVX0 U11571 ( .ZN(n9233), .INP(n18888) );
  INVX0 U11572 ( .ZN(n9234), .INP(n9233) );
  INVX0 U11574 ( .ZN(n9237), .INP(n18890) );
  INVX0 U11575 ( .ZN(n9238), .INP(n9237) );
  INVX0 U11577 ( .ZN(n9241), .INP(n18892) );
  INVX0 U11578 ( .ZN(n9242), .INP(n9241) );
  INVX0 U11580 ( .ZN(n9245), .INP(n18894) );
  INVX0 U11581 ( .ZN(n9246), .INP(n9245) );
  INVX0 U11583 ( .ZN(n9249), .INP(n18896) );
  INVX0 U11584 ( .ZN(n9250), .INP(n9249) );
  INVX0 U11586 ( .ZN(n9253), .INP(n18898) );
  INVX0 U11587 ( .ZN(n9254), .INP(n9253) );
  INVX0 U11589 ( .ZN(n9257), .INP(n18900) );
  INVX0 U11590 ( .ZN(n9258), .INP(n9257) );
  INVX0 U11592 ( .ZN(n9261), .INP(n18902) );
  INVX0 U11593 ( .ZN(n9262), .INP(n9261) );
  INVX0 U11595 ( .ZN(n9265), .INP(n18942) );
  INVX0 U11596 ( .ZN(n9266), .INP(n9265) );
  INVX0 U11598 ( .ZN(n9269), .INP(n18944) );
  INVX0 U11599 ( .ZN(n9270), .INP(n9269) );
  INVX0 U11601 ( .ZN(n9273), .INP(n18946) );
  INVX0 U11602 ( .ZN(n9274), .INP(n9273) );
  INVX0 U11325 ( .ZN(n8905), .INP(n18474) );
  INVX0 U11326 ( .ZN(n8906), .INP(n8905) );
  INVX0 U11328 ( .ZN(n8909), .INP(n18476) );
  INVX0 U11329 ( .ZN(n8910), .INP(n8909) );
  INVX0 U11331 ( .ZN(n8913), .INP(n18478) );
  INVX0 U11332 ( .ZN(n8914), .INP(n8913) );
  INVX0 U11334 ( .ZN(n8917), .INP(n18480) );
  INVX0 U11335 ( .ZN(n8918), .INP(n8917) );
  INVX0 U11337 ( .ZN(n8921), .INP(n18482) );
  INVX0 U11338 ( .ZN(n8922), .INP(n8921) );
  INVX0 U11340 ( .ZN(n8925), .INP(n18484) );
  INVX0 U11341 ( .ZN(n8926), .INP(n8925) );
  INVX0 U11343 ( .ZN(n8929), .INP(n18486) );
  INVX0 U11344 ( .ZN(n8930), .INP(n8929) );
  INVX0 U11346 ( .ZN(n8933), .INP(n18488) );
  INVX0 U11347 ( .ZN(n8934), .INP(n8933) );
  INVX0 U11349 ( .ZN(n8937), .INP(n18490) );
  INVX0 U11350 ( .ZN(n8938), .INP(n8937) );
  INVX0 U11352 ( .ZN(n8941), .INP(n18492) );
  INVX0 U11353 ( .ZN(n8942), .INP(n8941) );
  INVX0 U11355 ( .ZN(n8945), .INP(n18494) );
  INVX0 U11356 ( .ZN(n8946), .INP(n8945) );
  INVX0 U11358 ( .ZN(n8949), .INP(n18496) );
  INVX0 U11359 ( .ZN(n8950), .INP(n8949) );
  INVX0 U11361 ( .ZN(n8953), .INP(n18498) );
  INVX0 U11362 ( .ZN(n8954), .INP(n8953) );
  INVX0 U11364 ( .ZN(n8957), .INP(n18500) );
  INVX0 U11365 ( .ZN(n8958), .INP(n8957) );
  INVX0 U11367 ( .ZN(n8961), .INP(n18502) );
  INVX0 U11368 ( .ZN(n8962), .INP(n8961) );
  INVX0 U11370 ( .ZN(n8965), .INP(n18504) );
  INVX0 U11371 ( .ZN(n8966), .INP(n8965) );
  INVX0 U11373 ( .ZN(n8969), .INP(n18506) );
  INVX0 U11374 ( .ZN(n8970), .INP(n8969) );
  INVX0 U11376 ( .ZN(n8973), .INP(n18508) );
  INVX0 U11377 ( .ZN(n8974), .INP(n8973) );
  INVX0 U11379 ( .ZN(n8977), .INP(n18510) );
  INVX0 U11380 ( .ZN(n8978), .INP(n8977) );
  INVX0 U11382 ( .ZN(n8981), .INP(n18512) );
  INVX0 U11383 ( .ZN(n8982), .INP(n8981) );
  INVX0 U11385 ( .ZN(n8985), .INP(n18514) );
  INVX0 U11386 ( .ZN(n8986), .INP(n8985) );
  INVX0 U11388 ( .ZN(n8989), .INP(n18516) );
  INVX0 U11389 ( .ZN(n8990), .INP(n8989) );
  INVX0 U11391 ( .ZN(n8993), .INP(n18518) );
  INVX0 U11392 ( .ZN(n8994), .INP(n8993) );
  INVX0 U11394 ( .ZN(n8997), .INP(n18520) );
  INVX0 U11395 ( .ZN(n8998), .INP(n8997) );
  INVX0 U11397 ( .ZN(n9001), .INP(n18522) );
  INVX0 U11398 ( .ZN(n9002), .INP(n9001) );
  INVX0 U11400 ( .ZN(n9005), .INP(n18524) );
  INVX0 U11401 ( .ZN(n9006), .INP(n9005) );
  INVX0 U11403 ( .ZN(n9009), .INP(n18526) );
  INVX0 U11404 ( .ZN(n9010), .INP(n9009) );
  INVX0 U11406 ( .ZN(n9013), .INP(n18528) );
  INVX0 U11407 ( .ZN(n9014), .INP(n9013) );
  INVX0 U11409 ( .ZN(n9017), .INP(n18530) );
  INVX0 U11410 ( .ZN(n9018), .INP(n9017) );
  INVX0 U11412 ( .ZN(n9021), .INP(n18532) );
  INVX0 U11413 ( .ZN(n9022), .INP(n9021) );
  INVX0 U11415 ( .ZN(n9025), .INP(n18534) );
  INVX0 U11416 ( .ZN(n9026), .INP(n9025) );
  INVX0 U11418 ( .ZN(n9029), .INP(n18536) );
  INVX0 U11419 ( .ZN(n9030), .INP(n9029) );
  INVX0 U11421 ( .ZN(n9033), .INP(n18538) );
  INVX0 U11422 ( .ZN(n9034), .INP(n9033) );
  INVX0 U11424 ( .ZN(n9037), .INP(n18540) );
  INVX0 U11425 ( .ZN(n9038), .INP(n9037) );
  INVX0 U11427 ( .ZN(n9041), .INP(n18542) );
  INVX0 U11428 ( .ZN(n9042), .INP(n9041) );
  INVX0 U11430 ( .ZN(n9045), .INP(n18544) );
  INVX0 U11431 ( .ZN(n9046), .INP(n9045) );
  INVX0 U11433 ( .ZN(n9049), .INP(n18546) );
  INVX0 U11434 ( .ZN(n9050), .INP(n9049) );
  INVX0 U11436 ( .ZN(n9053), .INP(n18548) );
  INVX0 U11437 ( .ZN(n9054), .INP(n9053) );
  INVX0 U11439 ( .ZN(n9057), .INP(n18586) );
  INVX0 U11440 ( .ZN(n9058), .INP(n9057) );
  INVX0 U11442 ( .ZN(n9061), .INP(n18588) );
  INVX0 U11443 ( .ZN(n9062), .INP(n9061) );
  INVX0 U11445 ( .ZN(n9065), .INP(n18590) );
  INVX0 U11446 ( .ZN(n9066), .INP(n9065) );
  INVX0 U11448 ( .ZN(n9069), .INP(n18592) );
  INVX0 U11449 ( .ZN(n9070), .INP(n9069) );
  INVX0 U11451 ( .ZN(n9073), .INP(n18594) );
  INVX0 U11452 ( .ZN(n9074), .INP(n9073) );
  INVX0 U11454 ( .ZN(n9077), .INP(n18596) );
  INVX0 U11455 ( .ZN(n9078), .INP(n9077) );
  INVX0 U11457 ( .ZN(n9081), .INP(n18598) );
  INVX0 U11458 ( .ZN(n9082), .INP(n9081) );
  INVX0 U11460 ( .ZN(n9085), .INP(n18600) );
  INVX0 U11461 ( .ZN(n9086), .INP(n9085) );
  INVX0 U11463 ( .ZN(n9089), .INP(n18602) );
  INVX0 U8781 ( .ZN(n6371), .INP(P2_N196) );
  NAND2X0 U8782 ( .IN1(P2_N244), .IN2(n6371), .QN(n6370) );
  INVX0 U8783 ( .ZN(n6376), .INP(P2_N244) );
  NAND2X0 U8784 ( .IN1(P2_N196), .IN2(n6376), .QN(n6369) );
  NAND2X0 U8785 ( .IN1(n6370), .IN2(n6369), .QN(P2_N245) );
  NOR2X0 U8786 ( .QN(n6372), .IN1(n6371), .IN2(n6376) );
  NAND2X0 U8788 ( .IN1(n6372), .IN2(n7350), .QN(n6374) );
  OR2X1 U8789 ( .IN2(n6372), .IN1(n7350), .Q(n6373) );
  NAND2X0 U8790 ( .IN1(n6374), .IN2(n6373), .QN(P2_N246) );
  NOR2X0 U8791 ( .QN(n6377), .IN1(n6376), .IN2(n7350) );
  NAND2X0 U8792 ( .IN1(n6377), .IN2(P2_N196), .QN(n6378) );
  OR2X1 U8793 ( .IN2(P2_N194), .IN1(n6378), .Q(n6380) );
  NAND2X0 U8794 ( .IN1(P2_N194), .IN2(n6378), .QN(n6379) );
  NAND2X0 U8795 ( .IN1(n6380), .IN2(n6379), .QN(P2_N247) );
  AND2X1 U8796 ( .IN1(P2_N247), .IN2(P2_N246), .Q(n6381) );
  INVX0 U8798 ( .ZN(n6392), .INP(P2_N252) );
  NAND2X0 U8799 ( .IN1(P2_N290), .IN2(n6392), .QN(n6383) );
  INVX0 U8800 ( .ZN(n6391), .INP(P2_N290) );
  NAND2X0 U8801 ( .IN1(P2_N252), .IN2(n6391), .QN(n6382) );
  NAND2X0 U8803 ( .IN1(P2_N290), .IN2(P2_N252), .QN(n6386) );
  OR2X1 U8804 ( .IN2(P2_N251), .IN1(n6386), .Q(n6385) );
  NAND2X0 U8805 ( .IN1(P2_N251), .IN2(n6386), .QN(n6384) );
  INVX0 U8807 ( .ZN(n6393), .INP(P2_N251) );
  NOR2X0 U8808 ( .QN(n6387), .IN1(n6386), .IN2(n6393) );
  NAND2X0 U8810 ( .IN1(n6387), .IN2(n7353), .QN(n6389) );
  OR2X1 U8811 ( .IN2(n6387), .IN1(n7353), .Q(n6388) );
  NOR2X0 U8813 ( .QN(n6395), .IN1(n6391), .IN2(n7353) );
  NOR2X0 U8814 ( .QN(n6394), .IN1(n6393), .IN2(n6392) );
  NAND2X0 U8815 ( .IN1(n6395), .IN2(n6394), .QN(n6396) );
  OR2X1 U8816 ( .IN2(P2_N249), .IN1(n6396), .Q(n6398) );
  NAND2X0 U8817 ( .IN1(P2_N249), .IN2(n6396), .QN(n6397) );
  INVX0 U8819 ( .ZN(n6399), .INP(P2_N190) );
  OR2X1 U8820 ( .IN2(P2_N136), .IN1(n6399), .Q(n6401) );
  NAND2X0 U8821 ( .IN1(P2_N136), .IN2(n6399), .QN(n6400) );
  NAND2X0 U8823 ( .IN1(P2_N136), .IN2(P2_N190), .QN(n6402) );
  OR2X1 U8824 ( .IN2(P2_N135), .IN1(n6402), .Q(n6404) );
  NAND2X0 U8825 ( .IN1(P2_N135), .IN2(n6402), .QN(n6403) );
  INVX0 U8827 ( .ZN(n6405), .INP(P2_N245) );
  NOR2X0 U8828 ( .QN(n6406), .IN1(P2_N246), .IN2(n6405) );
  AND2X1 U8829 ( .IN1(n6406), .IN2(P2_N247), .Q(P2_N504) );
  NOR2X0 U8830 ( .QN(n6407), .IN1(P2_N246), .IN2(P2_N245) );
  AND2X1 U8831 ( .IN1(n6407), .IN2(P2_N247), .Q(P2_N508) );
  NOR2X0 U8833 ( .QN(n6409), .IN1(P2_N247), .IN2(n6405) );
  AND2X1 U8834 ( .IN1(n6409), .IN2(P2_N246), .Q(P2_N511) );
  NOR2X0 U8835 ( .QN(n6410), .IN1(P2_N247), .IN2(P2_N245) );
  AND2X1 U8836 ( .IN1(n6410), .IN2(P2_N246), .Q(P2_N514) );
  NOR2X0 U8837 ( .QN(n6411), .IN1(P2_N247), .IN2(P2_N246) );
  AND2X1 U8838 ( .IN1(n6411), .IN2(P2_N245), .Q(P2_N517) );
  OR2X1 U8839 ( .IN2(P2_N246), .IN1(P2_N247), .Q(n6412) );
  NOR2X0 U8840 ( .QN(P2_N519), .IN1(P2_N245), .IN2(n6412) );
  INVX0 U8841 ( .ZN(n6413), .INP(P2_N455) );
  OR2X1 U8842 ( .IN2(P2_N397), .IN1(n6413), .Q(n6415) );
  NAND2X0 U8843 ( .IN1(P2_N397), .IN2(n6413), .QN(n6414) );
  NAND2X0 U8845 ( .IN1(P2_N397), .IN2(P2_N455), .QN(n6416) );
  OR2X1 U8846 ( .IN2(P2_N396), .IN1(n6416), .Q(n6418) );
  NAND2X0 U8847 ( .IN1(P2_N396), .IN2(n6416), .QN(n6417) );
  AND2X1 U8849 ( .IN1(P1_N247), .IN2(P1_N246), .Q(n6419) );
  AND2X1 U8850 ( .IN1(n6419), .IN2(P1_N245), .Q(P1_N4969) );
  AND2X1 U8851 ( .IN1(P2_N247), .IN2(P2_N246), .Q(n6420) );
  AND2X1 U8852 ( .IN1(n6420), .IN2(P2_N245), .Q(P2_N4841) );
  INVX0 U11298 ( .ZN(n8869), .INP(n18198) );
  INVX0 U11299 ( .ZN(n8870), .INP(n8869) );
  INVX0 U11301 ( .ZN(n8873), .INP(n18200) );
  INVX0 U11302 ( .ZN(n8874), .INP(n8873) );
  INVX0 U11304 ( .ZN(n8877), .INP(n18202) );
  INVX0 U11305 ( .ZN(n8878), .INP(n8877) );
  INVX0 U11307 ( .ZN(n8881), .INP(n18289) );
  INVX0 U11308 ( .ZN(n8882), .INP(n8881) );
  INVX0 U11310 ( .ZN(n8885), .INP(n18291) );
  INVX0 U11311 ( .ZN(n8886), .INP(n8885) );
  INVX0 U11313 ( .ZN(n8889), .INP(n18466) );
  INVX0 U11314 ( .ZN(n8890), .INP(n8889) );
  INVX0 U11316 ( .ZN(n8893), .INP(n18468) );
  INVX0 U11317 ( .ZN(n8894), .INP(n8893) );
  INVX0 U11319 ( .ZN(n8897), .INP(n18470) );
  INVX0 U11320 ( .ZN(n8898), .INP(n8897) );
  INVX0 U11322 ( .ZN(n8901), .INP(n18472) );
  INVX0 U11323 ( .ZN(n8902), .INP(n8901) );
  NAND2X0 U8688 ( .IN1(N10), .IN2(n6736), .QN(n5943) );
  NAND2X0 U8689 ( .IN1(n9927), .IN2(n6737), .QN(n5942) );
  NAND2X0 U8690 ( .IN1(P1_N583), .IN2(P1_N360), .QN(n4145) );
  NAND2X0 U8691 ( .IN1(n4148), .IN2(n5944), .QN(P1_N1013) );
  NAND2X0 U8692 ( .IN1(n7026), .IN2(n4150), .QN(n5944) );
  NAND2X0 U8694 ( .IN1(n9931), .IN2(n6737), .QN(n5946) );
  NAND2X0 U8695 ( .IN1(N9), .IN2(n6736), .QN(n5945) );
  NAND2X0 U8696 ( .IN1(P1_N583), .IN2(P1_N361), .QN(n4148) );
  NAND2X0 U8697 ( .IN1(n4151), .IN2(n5947), .QN(P1_N1012) );
  NAND2X0 U8698 ( .IN1(n7022), .IN2(n4153), .QN(n5947) );
  NAND2X0 U8700 ( .IN1(n9337), .IN2(n6739), .QN(n5949) );
  NAND2X0 U8701 ( .IN1(N8), .IN2(n6736), .QN(n5948) );
  NAND2X0 U8702 ( .IN1(P1_N583), .IN2(P1_N362), .QN(n4151) );
  NAND2X0 U8703 ( .IN1(n4154), .IN2(n5950), .QN(P1_N1011) );
  NAND2X0 U8704 ( .IN1(n7022), .IN2(n4156), .QN(n5950) );
  NAND2X0 U8706 ( .IN1(n9389), .IN2(n6739), .QN(n5952) );
  NAND2X0 U8708 ( .IN1(N7), .IN2(N5), .QN(n5951) );
  NAND2X0 U8709 ( .IN1(P1_N583), .IN2(P1_N363), .QN(n4154) );
  INVX0 U8711 ( .ZN(n4158), .INP(n7330) );
  INVX0 U8712 ( .ZN(n4157), .INP(n7331) );
  INVX0 U8713 ( .ZN(n6321), .INP(P1_N196) );
  NAND2X0 U8714 ( .IN1(P1_N244), .IN2(n6321), .QN(n6320) );
  INVX0 U8715 ( .ZN(n6326), .INP(P1_N244) );
  NAND2X0 U8716 ( .IN1(P1_N196), .IN2(n6326), .QN(n6319) );
  NAND2X0 U8717 ( .IN1(n6320), .IN2(n6319), .QN(P1_N245) );
  NOR2X0 U8718 ( .QN(n6322), .IN1(n6321), .IN2(n6326) );
  NAND2X0 U8720 ( .IN1(n6322), .IN2(n7351), .QN(n6324) );
  OR2X1 U8721 ( .IN2(n6322), .IN1(n7351), .Q(n6323) );
  NAND2X0 U8722 ( .IN1(n6324), .IN2(n6323), .QN(P1_N246) );
  NOR2X0 U8723 ( .QN(n6327), .IN1(n6326), .IN2(n7351) );
  NAND2X0 U8724 ( .IN1(n6327), .IN2(P1_N196), .QN(n6328) );
  OR2X1 U8725 ( .IN2(P1_N194), .IN1(n6328), .Q(n6330) );
  NAND2X0 U8726 ( .IN1(P1_N194), .IN2(n6328), .QN(n6329) );
  NAND2X0 U8727 ( .IN1(n6330), .IN2(n6329), .QN(P1_N247) );
  AND2X1 U8728 ( .IN1(P1_N247), .IN2(P1_N246), .Q(n6331) );
  INVX0 U8730 ( .ZN(n6342), .INP(P1_N252) );
  NAND2X0 U8731 ( .IN1(P1_N290), .IN2(n6342), .QN(n6333) );
  INVX0 U8732 ( .ZN(n6341), .INP(P1_N290) );
  NAND2X0 U8733 ( .IN1(P1_N252), .IN2(n6341), .QN(n6332) );
  NAND2X0 U8735 ( .IN1(P1_N290), .IN2(P1_N252), .QN(n6336) );
  OR2X1 U8736 ( .IN2(P1_N251), .IN1(n6336), .Q(n6335) );
  NAND2X0 U8737 ( .IN1(P1_N251), .IN2(n6336), .QN(n6334) );
  INVX0 U8739 ( .ZN(n6343), .INP(P1_N251) );
  NOR2X0 U8740 ( .QN(n6337), .IN1(n6336), .IN2(n6343) );
  NAND2X0 U8742 ( .IN1(n6337), .IN2(n7352), .QN(n6339) );
  OR2X1 U8743 ( .IN2(n6337), .IN1(n7352), .Q(n6338) );
  NOR2X0 U8745 ( .QN(n6345), .IN1(n6341), .IN2(n7352) );
  NOR2X0 U8746 ( .QN(n6344), .IN1(n6343), .IN2(n6342) );
  NAND2X0 U8747 ( .IN1(n6345), .IN2(n6344), .QN(n6346) );
  OR2X1 U8748 ( .IN2(P1_N249), .IN1(n6346), .Q(n6348) );
  NAND2X0 U8749 ( .IN1(P1_N249), .IN2(n6346), .QN(n6347) );
  INVX0 U8751 ( .ZN(n6349), .INP(P1_N190) );
  OR2X1 U8752 ( .IN2(P1_N136), .IN1(n6349), .Q(n6351) );
  NAND2X0 U8753 ( .IN1(P1_N136), .IN2(n6349), .QN(n6350) );
  NAND2X0 U8755 ( .IN1(P1_N136), .IN2(P1_N190), .QN(n6352) );
  OR2X1 U8756 ( .IN2(P1_N135), .IN1(n6352), .Q(n6354) );
  NAND2X0 U8757 ( .IN1(P1_N135), .IN2(n6352), .QN(n6353) );
  INVX0 U8759 ( .ZN(n6355), .INP(P1_N245) );
  NOR2X0 U8760 ( .QN(n6356), .IN1(P1_N246), .IN2(n6355) );
  AND2X1 U8761 ( .IN1(n6356), .IN2(P1_N247), .Q(P1_N504) );
  NOR2X0 U8762 ( .QN(n6357), .IN1(P1_N246), .IN2(P1_N245) );
  AND2X1 U8763 ( .IN1(n6357), .IN2(P1_N247), .Q(P1_N508) );
  NOR2X0 U8765 ( .QN(n6359), .IN1(P1_N247), .IN2(n6355) );
  AND2X1 U8766 ( .IN1(n6359), .IN2(P1_N246), .Q(P1_N511) );
  NOR2X0 U8767 ( .QN(n6360), .IN1(P1_N247), .IN2(P1_N245) );
  AND2X1 U8768 ( .IN1(n6360), .IN2(P1_N246), .Q(P1_N514) );
  NOR2X0 U8769 ( .QN(n6361), .IN1(P1_N247), .IN2(P1_N246) );
  AND2X1 U8770 ( .IN1(n6361), .IN2(P1_N245), .Q(P1_N517) );
  OR2X1 U8771 ( .IN2(P1_N246), .IN1(P1_N247), .Q(n6362) );
  NOR2X0 U8772 ( .QN(P1_N519), .IN1(P1_N245), .IN2(n6362) );
  INVX0 U8773 ( .ZN(n6363), .INP(P1_N455) );
  OR2X1 U8774 ( .IN2(P1_N397), .IN1(n6363), .Q(n6365) );
  NAND2X0 U8775 ( .IN1(P1_N397), .IN2(n6363), .QN(n6364) );
  NAND2X0 U8777 ( .IN1(P1_N397), .IN2(P1_N455), .QN(n6366) );
  OR2X1 U8778 ( .IN2(P1_N396), .IN1(n6366), .Q(n6368) );
  NAND2X0 U8779 ( .IN1(P1_N396), .IN2(n6366), .QN(n6367) );
  NAND2X0 U8594 ( .IN1(P1_N583), .IN2(P1_N344), .QN(n4097) );
  NAND2X0 U8595 ( .IN1(n4100), .IN2(n5896), .QN(P1_N1029) );
  NAND2X0 U8596 ( .IN1(n7028), .IN2(n4102), .QN(n5896) );
  NAND2X0 U8597 ( .IN1(n5897), .IN2(n5898), .QN(n4102) );
  NAND2X0 U8598 ( .IN1(N25), .IN2(n6736), .QN(n5898) );
  NAND2X0 U8599 ( .IN1(n10059), .IN2(n6737), .QN(n5897) );
  NAND2X0 U8600 ( .IN1(P1_N583), .IN2(P1_N345), .QN(n4100) );
  NAND2X0 U8601 ( .IN1(n4103), .IN2(n5899), .QN(P1_N1028) );
  NAND2X0 U8602 ( .IN1(n7028), .IN2(n4105), .QN(n5899) );
  NAND2X0 U8603 ( .IN1(n5900), .IN2(n5901), .QN(n4105) );
  NAND2X0 U8604 ( .IN1(N24), .IN2(n6736), .QN(n5901) );
  NAND2X0 U8605 ( .IN1(n10063), .IN2(n6737), .QN(n5900) );
  NAND2X0 U8606 ( .IN1(P1_N583), .IN2(P1_N346), .QN(n4103) );
  NAND2X0 U8607 ( .IN1(n4106), .IN2(n5902), .QN(P1_N1027) );
  NAND2X0 U8608 ( .IN1(n7028), .IN2(n4108), .QN(n5902) );
  NAND2X0 U8610 ( .IN1(N23), .IN2(n6736), .QN(n5904) );
  NAND2X0 U8611 ( .IN1(n10067), .IN2(n6737), .QN(n5903) );
  NAND2X0 U8612 ( .IN1(P1_N583), .IN2(P1_N347), .QN(n4106) );
  NAND2X0 U8613 ( .IN1(n4109), .IN2(n5905), .QN(P1_N1026) );
  NAND2X0 U8614 ( .IN1(n7028), .IN2(n4111), .QN(n5905) );
  NAND2X0 U8616 ( .IN1(N22), .IN2(n6736), .QN(n5907) );
  NAND2X0 U8617 ( .IN1(n10071), .IN2(n6737), .QN(n5906) );
  NAND2X0 U8618 ( .IN1(P1_N583), .IN2(P1_N348), .QN(n4109) );
  NAND2X0 U8619 ( .IN1(n4112), .IN2(n5908), .QN(P1_N1025) );
  NAND2X0 U8620 ( .IN1(n7028), .IN2(n4114), .QN(n5908) );
  NAND2X0 U8622 ( .IN1(N21), .IN2(n6736), .QN(n5910) );
  NAND2X0 U8623 ( .IN1(n10075), .IN2(n6737), .QN(n5909) );
  NAND2X0 U8625 ( .IN1(n4115), .IN2(n5911), .QN(P1_N1024) );
  NAND2X0 U8626 ( .IN1(n7024), .IN2(n4117), .QN(n5911) );
  NAND2X0 U8628 ( .IN1(N20), .IN2(n6736), .QN(n5913) );
  NAND2X0 U8629 ( .IN1(n10079), .IN2(n6737), .QN(n5912) );
  NAND2X0 U8631 ( .IN1(n4118), .IN2(n5914), .QN(P1_N1023) );
  NAND2X0 U8632 ( .IN1(n7024), .IN2(n4120), .QN(n5914) );
  NAND2X0 U8634 ( .IN1(N19), .IN2(n6736), .QN(n5916) );
  NAND2X0 U8635 ( .IN1(n10083), .IN2(n6737), .QN(n5915) );
  NAND2X0 U8637 ( .IN1(n4121), .IN2(n5917), .QN(P1_N1022) );
  NAND2X0 U8638 ( .IN1(n7024), .IN2(n4123), .QN(n5917) );
  NAND2X0 U8640 ( .IN1(N18), .IN2(n6736), .QN(n5919) );
  NAND2X0 U8641 ( .IN1(n10087), .IN2(n6737), .QN(n5918) );
  NAND2X0 U8643 ( .IN1(n4124), .IN2(n5920), .QN(P1_N1021) );
  NAND2X0 U8644 ( .IN1(n7024), .IN2(n4126), .QN(n5920) );
  NAND2X0 U8646 ( .IN1(N17), .IN2(n6736), .QN(n5922) );
  NAND2X0 U8647 ( .IN1(n10091), .IN2(n6737), .QN(n5921) );
  NAND2X0 U8649 ( .IN1(n4127), .IN2(n5923), .QN(P1_N1020) );
  NAND2X0 U8650 ( .IN1(n7463), .IN2(n4129), .QN(n5923) );
  NAND2X0 U8652 ( .IN1(N16), .IN2(n6736), .QN(n5925) );
  NAND2X0 U8653 ( .IN1(n9903), .IN2(n6737), .QN(n5924) );
  NAND2X0 U8655 ( .IN1(n4130), .IN2(n5926), .QN(P1_N1019) );
  NAND2X0 U8656 ( .IN1(n7463), .IN2(n4132), .QN(n5926) );
  NAND2X0 U8657 ( .IN1(n5927), .IN2(n5928), .QN(n4132) );
  NAND2X0 U8658 ( .IN1(N15), .IN2(n6736), .QN(n5928) );
  NAND2X0 U8659 ( .IN1(n9907), .IN2(n6737), .QN(n5927) );
  NAND2X0 U8660 ( .IN1(P1_N583), .IN2(P1_N355), .QN(n4130) );
  NAND2X0 U8661 ( .IN1(n4133), .IN2(n5929), .QN(P1_N1018) );
  NAND2X0 U8662 ( .IN1(n7463), .IN2(n4135), .QN(n5929) );
  NAND2X0 U8663 ( .IN1(n5930), .IN2(n5931), .QN(n4135) );
  NAND2X0 U8664 ( .IN1(N14), .IN2(n6736), .QN(n5931) );
  NAND2X0 U8665 ( .IN1(n9911), .IN2(n6737), .QN(n5930) );
  NAND2X0 U8666 ( .IN1(P1_N583), .IN2(P1_N356), .QN(n4133) );
  NAND2X0 U8667 ( .IN1(n4136), .IN2(n5932), .QN(P1_N1017) );
  NAND2X0 U8668 ( .IN1(n7463), .IN2(n4138), .QN(n5932) );
  NAND2X0 U8670 ( .IN1(N13), .IN2(n6736), .QN(n5934) );
  NAND2X0 U8671 ( .IN1(n9915), .IN2(n6737), .QN(n5933) );
  NAND2X0 U8673 ( .IN1(n4139), .IN2(n5935), .QN(P1_N1016) );
  NAND2X0 U8674 ( .IN1(n7026), .IN2(n4141), .QN(n5935) );
  NAND2X0 U8676 ( .IN1(N12), .IN2(n6736), .QN(n5937) );
  NAND2X0 U8677 ( .IN1(n9919), .IN2(n6737), .QN(n5936) );
  NAND2X0 U8678 ( .IN1(P1_N583), .IN2(P1_N358), .QN(n4139) );
  NAND2X0 U8679 ( .IN1(n4142), .IN2(n5938), .QN(P1_N1015) );
  NAND2X0 U8680 ( .IN1(n7026), .IN2(n4144), .QN(n5938) );
  NAND2X0 U8682 ( .IN1(N11), .IN2(n6736), .QN(n5940) );
  NAND2X0 U8683 ( .IN1(n9923), .IN2(n6737), .QN(n5939) );
  NAND2X0 U8684 ( .IN1(P1_N583), .IN2(P1_N359), .QN(n4142) );
  NAND2X0 U8685 ( .IN1(n4145), .IN2(n5941), .QN(P1_N1014) );
  NAND2X0 U8686 ( .IN1(n7026), .IN2(n4147), .QN(n5941) );
  AND2X1 U8500 ( .IN1(n5840), .IN2(n5841), .Q(n5838) );
  NAND2X0 U8501 ( .IN1(P1_N355), .IN2(n6996), .QN(n5841) );
  NAND2X0 U8502 ( .IN1(n203), .IN2(n7337), .QN(n5840) );
  NAND2X0 U8503 ( .IN1(n5842), .IN2(n5843), .QN(P1_N670) );
  NAND2X0 U8504 ( .IN1(n183), .IN2(n7340), .QN(n5843) );
  AND2X1 U8505 ( .IN1(n5844), .IN2(n5845), .Q(n5842) );
  NAND2X0 U8506 ( .IN1(P1_N356), .IN2(n6996), .QN(n5845) );
  NAND2X0 U8507 ( .IN1(n204), .IN2(n7337), .QN(n5844) );
  NAND2X0 U8508 ( .IN1(n5846), .IN2(n5847), .QN(P1_N669) );
  NAND2X0 U8509 ( .IN1(n184), .IN2(n7340), .QN(n5847) );
  AND2X1 U8510 ( .IN1(n5848), .IN2(n5849), .Q(n5846) );
  NAND2X0 U8511 ( .IN1(P1_N357), .IN2(n6996), .QN(n5849) );
  NAND2X0 U8512 ( .IN1(n205), .IN2(n7337), .QN(n5848) );
  NAND2X0 U8513 ( .IN1(n5850), .IN2(n5851), .QN(P1_N668) );
  NAND2X0 U8514 ( .IN1(n185), .IN2(n7340), .QN(n5851) );
  AND2X1 U8515 ( .IN1(n5852), .IN2(n5853), .Q(n5850) );
  NAND2X0 U8516 ( .IN1(P1_N358), .IN2(n6996), .QN(n5853) );
  NAND2X0 U8517 ( .IN1(n206), .IN2(n7337), .QN(n5852) );
  NAND2X0 U8518 ( .IN1(n5854), .IN2(n5855), .QN(P1_N667) );
  NAND2X0 U8519 ( .IN1(n186), .IN2(n7340), .QN(n5855) );
  AND2X1 U8520 ( .IN1(n5856), .IN2(n5857), .Q(n5854) );
  NAND2X0 U8521 ( .IN1(P1_N359), .IN2(n6996), .QN(n5857) );
  NAND2X0 U8522 ( .IN1(n207), .IN2(n7337), .QN(n5856) );
  NAND2X0 U8523 ( .IN1(n5858), .IN2(n5859), .QN(P1_N666) );
  NAND2X0 U8524 ( .IN1(n187), .IN2(n7340), .QN(n5859) );
  AND2X1 U8525 ( .IN1(n5860), .IN2(n5861), .Q(n5858) );
  NAND2X0 U8526 ( .IN1(P1_N360), .IN2(n6996), .QN(n5861) );
  NAND2X0 U8527 ( .IN1(n208), .IN2(n7337), .QN(n5860) );
  NAND2X0 U8528 ( .IN1(n5862), .IN2(n5863), .QN(P1_N665) );
  NAND2X0 U8529 ( .IN1(n188), .IN2(n7340), .QN(n5863) );
  AND2X1 U8530 ( .IN1(n5864), .IN2(n5865), .Q(n5862) );
  NAND2X0 U8531 ( .IN1(P1_N361), .IN2(n6996), .QN(n5865) );
  NAND2X0 U8532 ( .IN1(n209), .IN2(n7337), .QN(n5864) );
  NAND2X0 U8533 ( .IN1(n5866), .IN2(n5867), .QN(P1_N664) );
  NAND2X0 U8534 ( .IN1(n189), .IN2(n7340), .QN(n5867) );
  AND2X1 U8535 ( .IN1(n5868), .IN2(n5869), .Q(n5866) );
  NAND2X0 U8536 ( .IN1(P1_N362), .IN2(n6996), .QN(n5869) );
  NAND2X0 U8537 ( .IN1(n210), .IN2(n7337), .QN(n5868) );
  NAND2X0 U8538 ( .IN1(n5870), .IN2(n5871), .QN(P1_N663) );
  NAND2X0 U8539 ( .IN1(n190), .IN2(n7340), .QN(n5871) );
  AND2X1 U8540 ( .IN1(n5872), .IN2(n5873), .Q(n5870) );
  NAND2X0 U8541 ( .IN1(P1_N363), .IN2(n6996), .QN(n5873) );
  NAND2X0 U8542 ( .IN1(n211), .IN2(n7337), .QN(n5872) );
  NOR2X0 U8543 ( .QN(P1_N1039), .IN1(n7326), .IN2(n7029) );
  NAND2X0 U8545 ( .IN1(n5875), .IN2(n5876), .QN(n4184) );
  NAND2X0 U8546 ( .IN1(N35), .IN2(N5), .QN(n5876) );
  NAND2X0 U8547 ( .IN1(n10019), .IN2(n6739), .QN(n5875) );
  NOR2X0 U8548 ( .QN(P1_N1038), .IN1(n7324), .IN2(n7029) );
  NAND2X0 U8550 ( .IN1(n5877), .IN2(n5878), .QN(n4187) );
  NAND2X0 U8551 ( .IN1(N34), .IN2(N5), .QN(n5878) );
  NAND2X0 U8552 ( .IN1(n10023), .IN2(n6739), .QN(n5877) );
  NOR2X0 U8553 ( .QN(P1_N1037), .IN1(n7322), .IN2(n7029) );
  NAND2X0 U8555 ( .IN1(n5879), .IN2(n5880), .QN(n4190) );
  NAND2X0 U8556 ( .IN1(N33), .IN2(N5), .QN(n5880) );
  NAND2X0 U8557 ( .IN1(n10027), .IN2(n6739), .QN(n5879) );
  NOR2X0 U8558 ( .QN(P1_N1036), .IN1(n7320), .IN2(n7029) );
  NAND2X0 U8560 ( .IN1(n5881), .IN2(n5882), .QN(n4193) );
  NAND2X0 U8561 ( .IN1(N32), .IN2(N5), .QN(n5882) );
  NAND2X0 U8562 ( .IN1(n10031), .IN2(n6739), .QN(n5881) );
  NOR2X0 U8563 ( .QN(P1_N1035), .IN1(n7318), .IN2(n7029) );
  NAND2X0 U8565 ( .IN1(n5883), .IN2(n5884), .QN(n4196) );
  NAND2X0 U8566 ( .IN1(N31), .IN2(N5), .QN(n5884) );
  NAND2X0 U8567 ( .IN1(n10035), .IN2(n6739), .QN(n5883) );
  NOR2X0 U8568 ( .QN(P1_N1034), .IN1(n7316), .IN2(n7027) );
  NAND2X0 U8570 ( .IN1(n5885), .IN2(n5886), .QN(n4199) );
  NAND2X0 U8571 ( .IN1(N30), .IN2(N5), .QN(n5886) );
  NAND2X0 U8572 ( .IN1(n10039), .IN2(n6739), .QN(n5885) );
  NOR2X0 U8573 ( .QN(P1_N1033), .IN1(n7314), .IN2(n7027) );
  NAND2X0 U8575 ( .IN1(n5887), .IN2(n5888), .QN(n4202) );
  NAND2X0 U8576 ( .IN1(N29), .IN2(N5), .QN(n5888) );
  NAND2X0 U8577 ( .IN1(n10043), .IN2(n6739), .QN(n5887) );
  NOR2X0 U8578 ( .QN(P1_N1032), .IN1(n7312), .IN2(n7027) );
  NAND2X0 U8580 ( .IN1(n5889), .IN2(n5890), .QN(n4205) );
  NAND2X0 U8581 ( .IN1(N28), .IN2(N5), .QN(n5890) );
  NAND2X0 U8582 ( .IN1(n10047), .IN2(n6739), .QN(n5889) );
  NOR2X0 U8583 ( .QN(P1_N1031), .IN1(n7310), .IN2(n7023) );
  NAND2X0 U8586 ( .IN1(n5891), .IN2(n5892), .QN(n4208) );
  NAND2X0 U8587 ( .IN1(N27), .IN2(N5), .QN(n5892) );
  NAND2X0 U8588 ( .IN1(n10051), .IN2(n6739), .QN(n5891) );
  NAND2X0 U8589 ( .IN1(n4097), .IN2(n5893), .QN(P1_N1030) );
  NAND2X0 U8590 ( .IN1(n7019), .IN2(n4099), .QN(n5893) );
  NAND2X0 U8592 ( .IN1(N26), .IN2(n6736), .QN(n5895) );
  NAND2X0 U8593 ( .IN1(n10055), .IN2(n6737), .QN(n5894) );
  NAND2X0 U8407 ( .IN1(n4103), .IN2(n5776), .QN(P1_N1119) );
  NAND2X0 U8408 ( .IN1(n7028), .IN2(n4105), .QN(n5776) );
  NAND2X0 U8409 ( .IN1(n4106), .IN2(n5777), .QN(P1_N1118) );
  NAND2X0 U8410 ( .IN1(n7028), .IN2(n4108), .QN(n5777) );
  NAND2X0 U8411 ( .IN1(n4109), .IN2(n5778), .QN(P1_N1117) );
  NAND2X0 U8412 ( .IN1(n7028), .IN2(n4111), .QN(n5778) );
  NAND2X0 U8413 ( .IN1(n4112), .IN2(n5779), .QN(P1_N1116) );
  NAND2X0 U8414 ( .IN1(n7028), .IN2(n4114), .QN(n5779) );
  NAND2X0 U8415 ( .IN1(n4115), .IN2(n5780), .QN(P1_N1115) );
  NAND2X0 U8416 ( .IN1(n7028), .IN2(n4117), .QN(n5780) );
  NAND2X0 U8417 ( .IN1(n4118), .IN2(n5781), .QN(P1_N1114) );
  NAND2X0 U8418 ( .IN1(n7024), .IN2(n4120), .QN(n5781) );
  NAND2X0 U8419 ( .IN1(n4121), .IN2(n5782), .QN(P1_N1113) );
  NAND2X0 U8420 ( .IN1(n7024), .IN2(n4123), .QN(n5782) );
  NAND2X0 U8421 ( .IN1(n4124), .IN2(n5783), .QN(P1_N1112) );
  NAND2X0 U8422 ( .IN1(n7024), .IN2(n4126), .QN(n5783) );
  NAND2X0 U8423 ( .IN1(n4127), .IN2(n5784), .QN(P1_N1111) );
  NAND2X0 U8424 ( .IN1(n7463), .IN2(n4129), .QN(n5784) );
  NAND2X0 U8425 ( .IN1(n4130), .IN2(n5785), .QN(P1_N1110) );
  NAND2X0 U8426 ( .IN1(n7463), .IN2(n4132), .QN(n5785) );
  NAND2X0 U8427 ( .IN1(n4133), .IN2(n5786), .QN(P1_N1109) );
  NAND2X0 U8428 ( .IN1(n7463), .IN2(n4135), .QN(n5786) );
  NAND2X0 U8429 ( .IN1(n4136), .IN2(n5787), .QN(P1_N1108) );
  NAND2X0 U8430 ( .IN1(n7463), .IN2(n4138), .QN(n5787) );
  NAND2X0 U8431 ( .IN1(n4139), .IN2(n5788), .QN(P1_N1107) );
  NAND2X0 U8432 ( .IN1(n7026), .IN2(n4141), .QN(n5788) );
  NAND2X0 U8433 ( .IN1(n4142), .IN2(n5789), .QN(P1_N1106) );
  NAND2X0 U8434 ( .IN1(n7026), .IN2(n4144), .QN(n5789) );
  NAND2X0 U8435 ( .IN1(n4145), .IN2(n5790), .QN(P1_N1105) );
  NAND2X0 U8436 ( .IN1(n7026), .IN2(n4147), .QN(n5790) );
  NAND2X0 U8437 ( .IN1(n4148), .IN2(n5791), .QN(P1_N1104) );
  NAND2X0 U8438 ( .IN1(n7026), .IN2(n4150), .QN(n5791) );
  NAND2X0 U8439 ( .IN1(n4151), .IN2(n5792), .QN(P1_N1103) );
  NAND2X0 U8440 ( .IN1(n7022), .IN2(n4153), .QN(n5792) );
  NAND2X0 U8441 ( .IN1(n4154), .IN2(n5793), .QN(P1_N1102) );
  NAND2X0 U8442 ( .IN1(n7022), .IN2(n4156), .QN(n5793) );
  NAND2X0 U8443 ( .IN1(n5794), .IN2(n5795), .QN(P1_N682) );
  NAND2X0 U8444 ( .IN1(n171), .IN2(n7340), .QN(n5795) );
  AND2X1 U8445 ( .IN1(n5796), .IN2(n5797), .Q(n5794) );
  NAND2X0 U8446 ( .IN1(n6996), .IN2(P1_N344), .QN(n5797) );
  NAND2X0 U8447 ( .IN1(n192), .IN2(n7337), .QN(n5796) );
  NAND2X0 U8448 ( .IN1(n5798), .IN2(n5799), .QN(P1_N681) );
  NAND2X0 U8449 ( .IN1(n172), .IN2(n7340), .QN(n5799) );
  AND2X1 U8450 ( .IN1(n5800), .IN2(n5801), .Q(n5798) );
  NAND2X0 U8451 ( .IN1(P1_N345), .IN2(n6996), .QN(n5801) );
  NAND2X0 U8452 ( .IN1(n193), .IN2(n7337), .QN(n5800) );
  NAND2X0 U8453 ( .IN1(n5802), .IN2(n5803), .QN(P1_N680) );
  NAND2X0 U8454 ( .IN1(n173), .IN2(n7340), .QN(n5803) );
  AND2X1 U8455 ( .IN1(n5804), .IN2(n5805), .Q(n5802) );
  NAND2X0 U8456 ( .IN1(P1_N346), .IN2(n6996), .QN(n5805) );
  NAND2X0 U8457 ( .IN1(n194), .IN2(n7337), .QN(n5804) );
  NAND2X0 U8458 ( .IN1(n5806), .IN2(n5807), .QN(P1_N679) );
  NAND2X0 U8459 ( .IN1(n174), .IN2(n7340), .QN(n5807) );
  AND2X1 U8460 ( .IN1(n5808), .IN2(n5809), .Q(n5806) );
  NAND2X0 U8461 ( .IN1(P1_N347), .IN2(n6996), .QN(n5809) );
  NAND2X0 U8462 ( .IN1(n195), .IN2(n7337), .QN(n5808) );
  NAND2X0 U8463 ( .IN1(n5810), .IN2(n5811), .QN(P1_N678) );
  NAND2X0 U8464 ( .IN1(n175), .IN2(n7340), .QN(n5811) );
  AND2X1 U8465 ( .IN1(n5812), .IN2(n5813), .Q(n5810) );
  NAND2X0 U8466 ( .IN1(P1_N348), .IN2(n6996), .QN(n5813) );
  NAND2X0 U8467 ( .IN1(n196), .IN2(n7337), .QN(n5812) );
  NAND2X0 U8468 ( .IN1(n5814), .IN2(n5815), .QN(P1_N677) );
  NAND2X0 U8469 ( .IN1(n176), .IN2(n7340), .QN(n5815) );
  AND2X1 U8470 ( .IN1(n5816), .IN2(n5817), .Q(n5814) );
  NAND2X0 U8471 ( .IN1(P1_N349), .IN2(n6996), .QN(n5817) );
  NAND2X0 U8472 ( .IN1(n197), .IN2(n7337), .QN(n5816) );
  NAND2X0 U8473 ( .IN1(n5818), .IN2(n5819), .QN(P1_N676) );
  NAND2X0 U8474 ( .IN1(n177), .IN2(n7340), .QN(n5819) );
  AND2X1 U8475 ( .IN1(n5820), .IN2(n5821), .Q(n5818) );
  NAND2X0 U8476 ( .IN1(P1_N350), .IN2(n6996), .QN(n5821) );
  NAND2X0 U8477 ( .IN1(n198), .IN2(n7337), .QN(n5820) );
  NAND2X0 U8478 ( .IN1(n5822), .IN2(n5823), .QN(P1_N675) );
  NAND2X0 U8479 ( .IN1(n178), .IN2(n7340), .QN(n5823) );
  AND2X1 U8480 ( .IN1(n5824), .IN2(n5825), .Q(n5822) );
  NAND2X0 U8481 ( .IN1(P1_N351), .IN2(n6996), .QN(n5825) );
  NAND2X0 U8482 ( .IN1(n199), .IN2(n7337), .QN(n5824) );
  NAND2X0 U8483 ( .IN1(n5826), .IN2(n5827), .QN(P1_N674) );
  NAND2X0 U8484 ( .IN1(n179), .IN2(n7340), .QN(n5827) );
  AND2X1 U8485 ( .IN1(n5828), .IN2(n5829), .Q(n5826) );
  NAND2X0 U8486 ( .IN1(P1_N352), .IN2(n6996), .QN(n5829) );
  NAND2X0 U8487 ( .IN1(n200), .IN2(n7337), .QN(n5828) );
  NAND2X0 U8488 ( .IN1(n5830), .IN2(n5831), .QN(P1_N673) );
  NAND2X0 U8489 ( .IN1(n180), .IN2(n7340), .QN(n5831) );
  AND2X1 U8490 ( .IN1(n5832), .IN2(n5833), .Q(n5830) );
  NAND2X0 U8491 ( .IN1(P1_N353), .IN2(n6996), .QN(n5833) );
  NAND2X0 U8492 ( .IN1(n201), .IN2(n7337), .QN(n5832) );
  NAND2X0 U8493 ( .IN1(n5834), .IN2(n5835), .QN(P1_N672) );
  NAND2X0 U8494 ( .IN1(n181), .IN2(n7340), .QN(n5835) );
  AND2X1 U8495 ( .IN1(n5836), .IN2(n5837), .Q(n5834) );
  NAND2X0 U8496 ( .IN1(P1_N354), .IN2(n6996), .QN(n5837) );
  NAND2X0 U8497 ( .IN1(n202), .IN2(n7337), .QN(n5836) );
  NAND2X0 U8498 ( .IN1(n5838), .IN2(n5839), .QN(P1_N671) );
  NAND2X0 U8499 ( .IN1(n182), .IN2(n7340), .QN(n5839) );
  NAND2X0 U8308 ( .IN1(n5721), .IN2(n5722), .QN(P1_N1307) );
  NAND2X0 U8309 ( .IN1(P1_N1124), .IN2(n5709), .QN(n5722) );
  NAND2X0 U8310 ( .IN1(P1_N386), .IN2(P1_N5572), .QN(n5721) );
  NAND2X0 U8311 ( .IN1(n5723), .IN2(n5724), .QN(P1_N1306) );
  NAND2X0 U8312 ( .IN1(P1_N1123), .IN2(n5709), .QN(n5724) );
  NAND2X0 U8313 ( .IN1(P1_N385), .IN2(P1_N5572), .QN(n5723) );
  NAND2X0 U8314 ( .IN1(n5725), .IN2(n5726), .QN(P1_N1305) );
  NAND2X0 U8315 ( .IN1(P1_N1122), .IN2(n5709), .QN(n5726) );
  NAND2X0 U8316 ( .IN1(P1_N384), .IN2(P1_N5572), .QN(n5725) );
  NAND2X0 U8317 ( .IN1(n5727), .IN2(n5728), .QN(P1_N1304) );
  NAND2X0 U8318 ( .IN1(n5709), .IN2(P1_N1121), .QN(n5728) );
  NAND2X0 U8319 ( .IN1(P1_N383), .IN2(P1_N5572), .QN(n5727) );
  NAND2X0 U8320 ( .IN1(n5729), .IN2(n5730), .QN(P1_N1303) );
  NAND2X0 U8321 ( .IN1(n5709), .IN2(P1_N1120), .QN(n5730) );
  NAND2X0 U8322 ( .IN1(P1_N382), .IN2(P1_N5572), .QN(n5729) );
  NAND2X0 U8323 ( .IN1(n5731), .IN2(n5732), .QN(P1_N1302) );
  NAND2X0 U8324 ( .IN1(n5709), .IN2(P1_N1119), .QN(n5732) );
  NAND2X0 U8325 ( .IN1(P1_N381), .IN2(P1_N5572), .QN(n5731) );
  NAND2X0 U8326 ( .IN1(n5733), .IN2(n5734), .QN(P1_N1301) );
  NAND2X0 U8327 ( .IN1(n5709), .IN2(P1_N1118), .QN(n5734) );
  NAND2X0 U8328 ( .IN1(P1_N380), .IN2(P1_N5572), .QN(n5733) );
  NAND2X0 U8329 ( .IN1(n5735), .IN2(n5736), .QN(P1_N1300) );
  NAND2X0 U8330 ( .IN1(n5709), .IN2(P1_N1117), .QN(n5736) );
  NAND2X0 U8331 ( .IN1(P1_N379), .IN2(P1_N5572), .QN(n5735) );
  NAND2X0 U8332 ( .IN1(n5737), .IN2(n5738), .QN(P1_N1299) );
  NAND2X0 U8333 ( .IN1(n5709), .IN2(P1_N1116), .QN(n5738) );
  NAND2X0 U8334 ( .IN1(P1_N378), .IN2(P1_N5572), .QN(n5737) );
  NAND2X0 U8335 ( .IN1(n5739), .IN2(n5740), .QN(P1_N1298) );
  NAND2X0 U8336 ( .IN1(n5709), .IN2(P1_N1115), .QN(n5740) );
  NAND2X0 U8337 ( .IN1(P1_N377), .IN2(P1_N5572), .QN(n5739) );
  NAND2X0 U8338 ( .IN1(n5741), .IN2(n5742), .QN(P1_N1297) );
  NAND2X0 U8339 ( .IN1(n5709), .IN2(P1_N1114), .QN(n5742) );
  NAND2X0 U8340 ( .IN1(P1_N376), .IN2(P1_N5572), .QN(n5741) );
  NAND2X0 U8341 ( .IN1(n5743), .IN2(n5744), .QN(P1_N1296) );
  NAND2X0 U8342 ( .IN1(n5709), .IN2(P1_N1113), .QN(n5744) );
  NAND2X0 U8343 ( .IN1(P1_N375), .IN2(P1_N5572), .QN(n5743) );
  NAND2X0 U8344 ( .IN1(n5745), .IN2(n5746), .QN(P1_N1295) );
  NAND2X0 U8345 ( .IN1(n5709), .IN2(P1_N1112), .QN(n5746) );
  NAND2X0 U8346 ( .IN1(P1_N374), .IN2(P1_N5572), .QN(n5745) );
  NAND2X0 U8347 ( .IN1(n5747), .IN2(n5748), .QN(P1_N1294) );
  NAND2X0 U8348 ( .IN1(n5709), .IN2(P1_N1111), .QN(n5748) );
  NAND2X0 U8349 ( .IN1(P1_N373), .IN2(P1_N5572), .QN(n5747) );
  NAND2X0 U8350 ( .IN1(n5749), .IN2(n5750), .QN(P1_N1293) );
  NAND2X0 U8351 ( .IN1(n5709), .IN2(P1_N1110), .QN(n5750) );
  NAND2X0 U8352 ( .IN1(P1_N372), .IN2(P1_N5572), .QN(n5749) );
  NAND2X0 U8353 ( .IN1(n5751), .IN2(n5752), .QN(P1_N1292) );
  NAND2X0 U8354 ( .IN1(n5709), .IN2(P1_N1109), .QN(n5752) );
  NAND2X0 U8355 ( .IN1(P1_N371), .IN2(P1_N5572), .QN(n5751) );
  NAND2X0 U8356 ( .IN1(n5753), .IN2(n5754), .QN(P1_N1291) );
  NAND2X0 U8357 ( .IN1(n5709), .IN2(P1_N1108), .QN(n5754) );
  NAND2X0 U8358 ( .IN1(P1_N370), .IN2(P1_N5572), .QN(n5753) );
  NAND2X0 U8359 ( .IN1(n5755), .IN2(n5756), .QN(P1_N1290) );
  NAND2X0 U8360 ( .IN1(n5709), .IN2(P1_N1107), .QN(n5756) );
  NAND2X0 U8361 ( .IN1(P1_N369), .IN2(P1_N5572), .QN(n5755) );
  NAND2X0 U8362 ( .IN1(n5757), .IN2(n5758), .QN(P1_N1289) );
  NAND2X0 U8363 ( .IN1(n5709), .IN2(P1_N1106), .QN(n5758) );
  NAND2X0 U8364 ( .IN1(P1_N368), .IN2(P1_N5572), .QN(n5757) );
  NAND2X0 U8365 ( .IN1(n5759), .IN2(n5760), .QN(P1_N1288) );
  NAND2X0 U8366 ( .IN1(n5709), .IN2(P1_N1105), .QN(n5760) );
  NAND2X0 U8367 ( .IN1(n18451), .IN2(P1_N5572), .QN(n5759) );
  NAND2X0 U8368 ( .IN1(n5761), .IN2(n5762), .QN(P1_N1287) );
  NAND2X0 U8369 ( .IN1(n5709), .IN2(P1_N1104), .QN(n5762) );
  NAND2X0 U8370 ( .IN1(n6623), .IN2(P1_N5572), .QN(n5761) );
  NAND2X0 U8371 ( .IN1(n5763), .IN2(n5764), .QN(P1_N1286) );
  NAND2X0 U8372 ( .IN1(n5709), .IN2(P1_N1103), .QN(n5764) );
  NAND2X0 U8373 ( .IN1(n6622), .IN2(P1_N5572), .QN(n5763) );
  NAND2X0 U8374 ( .IN1(n5765), .IN2(n5766), .QN(P1_N1285) );
  NAND2X0 U8375 ( .IN1(n5709), .IN2(P1_N1102), .QN(n5766) );
  NAND2X0 U8378 ( .IN1(n6621), .IN2(P1_N5572), .QN(n5765) );
  NAND2X0 U8383 ( .IN1(n7356), .IN2(n5769), .QN(P1_N1252) );
  NAND2X0 U8384 ( .IN1(n7355), .IN2(n5770), .QN(P1_N1250) );
  NOR2X0 U8385 ( .QN(P1_N1314), .IN1(n5770), .IN2(n5769) );
  INVX0 U8386 ( .ZN(n5769), .INP(n7355) );
  INVX0 U8387 ( .ZN(n5770), .INP(n7356) );
  NOR2X0 U8388 ( .QN(P1_N1131), .IN1(n7328), .IN2(n7029) );
  NAND2X0 U8390 ( .IN1(n5772), .IN2(n5773), .QN(n4181) );
  NAND2X0 U8391 ( .IN1(N36), .IN2(N5), .QN(n5773) );
  NAND2X0 U8392 ( .IN1(n10099), .IN2(n6739), .QN(n5772) );
  NOR2X0 U8393 ( .QN(P1_N1130), .IN1(n7029), .IN2(n7326) );
  NOR2X0 U8394 ( .QN(P1_N1129), .IN1(n7029), .IN2(n7324) );
  NOR2X0 U8395 ( .QN(P1_N1128), .IN1(n7029), .IN2(n7322) );
  NOR2X0 U8396 ( .QN(P1_N1127), .IN1(n7029), .IN2(n7320) );
  NOR2X0 U8397 ( .QN(P1_N1126), .IN1(n7029), .IN2(n7318) );
  NOR2X0 U8398 ( .QN(P1_N1125), .IN1(n7027), .IN2(n7316) );
  NOR2X0 U8399 ( .QN(P1_N1124), .IN1(n7027), .IN2(n7314) );
  NOR2X0 U8400 ( .QN(P1_N1123), .IN1(n7027), .IN2(n7312) );
  NOR2X0 U8401 ( .QN(P1_N1122), .IN1(n7023), .IN2(n7310) );
  NAND2X0 U8403 ( .IN1(n4097), .IN2(n5774), .QN(P1_N1121) );
  NAND2X0 U8404 ( .IN1(n7019), .IN2(n4099), .QN(n5774) );
  NAND2X0 U8405 ( .IN1(n4100), .IN2(n5775), .QN(P1_N1120) );
  NAND2X0 U8406 ( .IN1(n7028), .IN2(n4102), .QN(n5775) );
  NAND2X0 U8207 ( .IN1(P1_N370), .IN2(P1_N5573), .QN(n5667) );
  NAND2X0 U8208 ( .IN1(n5669), .IN2(n5670), .QN(P1_N1545) );
  NAND2X0 U8209 ( .IN1(n5623), .IN2(P1_N1362), .QN(n5670) );
  NAND2X0 U8210 ( .IN1(P1_N369), .IN2(P1_N5573), .QN(n5669) );
  NAND2X0 U8211 ( .IN1(n5671), .IN2(n5672), .QN(P1_N1544) );
  NAND2X0 U8212 ( .IN1(n5623), .IN2(P1_N1361), .QN(n5672) );
  NAND2X0 U8213 ( .IN1(P1_N368), .IN2(P1_N5573), .QN(n5671) );
  NAND2X0 U8214 ( .IN1(n5673), .IN2(n5674), .QN(P1_N1543) );
  NAND2X0 U8215 ( .IN1(n5623), .IN2(P1_N1360), .QN(n5674) );
  NAND2X0 U8216 ( .IN1(n18451), .IN2(P1_N5573), .QN(n5673) );
  NAND2X0 U8217 ( .IN1(n5675), .IN2(n5676), .QN(P1_N1542) );
  NAND2X0 U8218 ( .IN1(n5623), .IN2(P1_N1359), .QN(n5676) );
  NAND2X0 U8219 ( .IN1(n6623), .IN2(P1_N5573), .QN(n5675) );
  NAND2X0 U8220 ( .IN1(n5677), .IN2(n5678), .QN(P1_N1541) );
  NAND2X0 U8221 ( .IN1(n5623), .IN2(P1_N1358), .QN(n5678) );
  NAND2X0 U8222 ( .IN1(n6622), .IN2(P1_N5573), .QN(n5677) );
  NAND2X0 U8223 ( .IN1(n5679), .IN2(n5680), .QN(P1_N1540) );
  NAND2X0 U8224 ( .IN1(n5623), .IN2(P1_N1357), .QN(n5680) );
  NAND2X0 U8227 ( .IN1(n6621), .IN2(P1_N5573), .QN(n5679) );
  NAND2X0 U8232 ( .IN1(n7358), .IN2(n5683), .QN(P1_N1507) );
  NAND2X0 U8233 ( .IN1(n7357), .IN2(n5684), .QN(P1_N1505) );
  NOR2X0 U8234 ( .QN(P1_N1569), .IN1(n5684), .IN2(n5683) );
  INVX0 U8235 ( .ZN(n5683), .INP(n7357) );
  INVX0 U8236 ( .ZN(n5684), .INP(n7358) );
  NOR2X0 U8237 ( .QN(P1_N1386), .IN1(n7328), .IN2(n7029) );
  NOR2X0 U8238 ( .QN(P1_N1385), .IN1(n7029), .IN2(n7326) );
  NOR2X0 U8239 ( .QN(P1_N1384), .IN1(n7029), .IN2(n7324) );
  NOR2X0 U8240 ( .QN(P1_N1383), .IN1(n7029), .IN2(n7322) );
  NOR2X0 U8241 ( .QN(P1_N1382), .IN1(n7029), .IN2(n7320) );
  NOR2X0 U8242 ( .QN(P1_N1381), .IN1(n7029), .IN2(n7318) );
  NOR2X0 U8243 ( .QN(P1_N1380), .IN1(n7027), .IN2(n7316) );
  NOR2X0 U8244 ( .QN(P1_N1379), .IN1(n7027), .IN2(n7314) );
  NOR2X0 U8245 ( .QN(P1_N1378), .IN1(n7027), .IN2(n7312) );
  NOR2X0 U8246 ( .QN(P1_N1377), .IN1(n7023), .IN2(n7310) );
  NAND2X0 U8248 ( .IN1(n4097), .IN2(n5686), .QN(P1_N1376) );
  NAND2X0 U8249 ( .IN1(n7019), .IN2(n4099), .QN(n5686) );
  NAND2X0 U8250 ( .IN1(n4100), .IN2(n5687), .QN(P1_N1375) );
  NAND2X0 U8251 ( .IN1(n7028), .IN2(n4102), .QN(n5687) );
  NAND2X0 U8252 ( .IN1(n4103), .IN2(n5688), .QN(P1_N1374) );
  NAND2X0 U8253 ( .IN1(n7028), .IN2(n4105), .QN(n5688) );
  NAND2X0 U8254 ( .IN1(n4106), .IN2(n5689), .QN(P1_N1373) );
  NAND2X0 U8255 ( .IN1(n7028), .IN2(n4108), .QN(n5689) );
  NAND2X0 U8256 ( .IN1(n4109), .IN2(n5690), .QN(P1_N1372) );
  NAND2X0 U8257 ( .IN1(n7028), .IN2(n4111), .QN(n5690) );
  NAND2X0 U8258 ( .IN1(n4112), .IN2(n5691), .QN(P1_N1371) );
  NAND2X0 U8259 ( .IN1(n7028), .IN2(n4114), .QN(n5691) );
  NAND2X0 U8260 ( .IN1(n4115), .IN2(n5692), .QN(P1_N1370) );
  NAND2X0 U8261 ( .IN1(n7024), .IN2(n4117), .QN(n5692) );
  NAND2X0 U8262 ( .IN1(n4118), .IN2(n5693), .QN(P1_N1369) );
  NAND2X0 U8263 ( .IN1(n7024), .IN2(n4120), .QN(n5693) );
  NAND2X0 U8264 ( .IN1(n4121), .IN2(n5694), .QN(P1_N1368) );
  NAND2X0 U8265 ( .IN1(n7024), .IN2(n4123), .QN(n5694) );
  NAND2X0 U8266 ( .IN1(n4124), .IN2(n5695), .QN(P1_N1367) );
  NAND2X0 U8267 ( .IN1(n7024), .IN2(n4126), .QN(n5695) );
  NAND2X0 U8268 ( .IN1(n4127), .IN2(n5696), .QN(P1_N1366) );
  NAND2X0 U8269 ( .IN1(n7463), .IN2(n4129), .QN(n5696) );
  NAND2X0 U8270 ( .IN1(n4130), .IN2(n5697), .QN(P1_N1365) );
  NAND2X0 U8271 ( .IN1(n7463), .IN2(n4132), .QN(n5697) );
  NAND2X0 U8272 ( .IN1(n4133), .IN2(n5698), .QN(P1_N1364) );
  NAND2X0 U8273 ( .IN1(n7463), .IN2(n4135), .QN(n5698) );
  NAND2X0 U8274 ( .IN1(n4136), .IN2(n5699), .QN(P1_N1363) );
  NAND2X0 U8275 ( .IN1(n7463), .IN2(n4138), .QN(n5699) );
  NAND2X0 U8276 ( .IN1(n4139), .IN2(n5700), .QN(P1_N1362) );
  NAND2X0 U8277 ( .IN1(n7026), .IN2(n4141), .QN(n5700) );
  NAND2X0 U8278 ( .IN1(n4142), .IN2(n5701), .QN(P1_N1361) );
  NAND2X0 U8279 ( .IN1(n7026), .IN2(n4144), .QN(n5701) );
  NAND2X0 U8280 ( .IN1(n4145), .IN2(n5702), .QN(P1_N1360) );
  NAND2X0 U8281 ( .IN1(n7026), .IN2(n4147), .QN(n5702) );
  NAND2X0 U8282 ( .IN1(n4148), .IN2(n5703), .QN(P1_N1359) );
  NAND2X0 U8283 ( .IN1(n7026), .IN2(n4150), .QN(n5703) );
  NAND2X0 U8284 ( .IN1(n4151), .IN2(n5704), .QN(P1_N1358) );
  NAND2X0 U8285 ( .IN1(n7022), .IN2(n4153), .QN(n5704) );
  NAND2X0 U8286 ( .IN1(n4154), .IN2(n5705), .QN(P1_N1357) );
  NAND2X0 U8287 ( .IN1(n7022), .IN2(n4156), .QN(n5705) );
  NAND2X0 U8290 ( .IN1(n5707), .IN2(n5708), .QN(P1_N1313) );
  NAND2X0 U8291 ( .IN1(P1_N1130), .IN2(n5709), .QN(n5708) );
  NAND2X0 U8292 ( .IN1(P1_N392), .IN2(P1_N5572), .QN(n5707) );
  NAND2X0 U8293 ( .IN1(n5711), .IN2(n5712), .QN(P1_N1312) );
  NAND2X0 U8294 ( .IN1(P1_N1129), .IN2(n5709), .QN(n5712) );
  NAND2X0 U8295 ( .IN1(P1_N391), .IN2(P1_N5572), .QN(n5711) );
  NAND2X0 U8296 ( .IN1(n5713), .IN2(n5714), .QN(P1_N1311) );
  NAND2X0 U8297 ( .IN1(P1_N1128), .IN2(n5709), .QN(n5714) );
  NAND2X0 U8298 ( .IN1(P1_N390), .IN2(P1_N5572), .QN(n5713) );
  NAND2X0 U8299 ( .IN1(n5715), .IN2(n5716), .QN(P1_N1310) );
  NAND2X0 U8300 ( .IN1(P1_N1127), .IN2(n5709), .QN(n5716) );
  NAND2X0 U8301 ( .IN1(P1_N389), .IN2(P1_N5572), .QN(n5715) );
  NAND2X0 U8302 ( .IN1(n5717), .IN2(n5718), .QN(P1_N1309) );
  NAND2X0 U8303 ( .IN1(P1_N1126), .IN2(n5709), .QN(n5718) );
  NAND2X0 U8304 ( .IN1(P1_N388), .IN2(P1_N5572), .QN(n5717) );
  NAND2X0 U8305 ( .IN1(n5719), .IN2(n5720), .QN(P1_N1308) );
  NAND2X0 U8306 ( .IN1(P1_N1125), .IN2(n5709), .QN(n5720) );
  NAND2X0 U8307 ( .IN1(P1_N387), .IN2(P1_N5572), .QN(n5719) );
  NAND2X0 U8112 ( .IN1(n7024), .IN2(n4120), .QN(n5607) );
  NAND2X0 U8113 ( .IN1(n4121), .IN2(n5608), .QN(P1_N1623) );
  NAND2X0 U8114 ( .IN1(n7024), .IN2(n4123), .QN(n5608) );
  NAND2X0 U8115 ( .IN1(n4124), .IN2(n5609), .QN(P1_N1622) );
  NAND2X0 U8116 ( .IN1(n7024), .IN2(n4126), .QN(n5609) );
  NAND2X0 U8117 ( .IN1(n4127), .IN2(n5610), .QN(P1_N1621) );
  NAND2X0 U8118 ( .IN1(n7463), .IN2(n4129), .QN(n5610) );
  NAND2X0 U8119 ( .IN1(n4130), .IN2(n5611), .QN(P1_N1620) );
  NAND2X0 U8120 ( .IN1(n7463), .IN2(n4132), .QN(n5611) );
  NAND2X0 U8121 ( .IN1(n4133), .IN2(n5612), .QN(P1_N1619) );
  NAND2X0 U8122 ( .IN1(n7463), .IN2(n4135), .QN(n5612) );
  NAND2X0 U8123 ( .IN1(n4136), .IN2(n5613), .QN(P1_N1618) );
  NAND2X0 U8124 ( .IN1(n7463), .IN2(n4138), .QN(n5613) );
  NAND2X0 U8125 ( .IN1(n4139), .IN2(n5614), .QN(P1_N1617) );
  NAND2X0 U8126 ( .IN1(n7026), .IN2(n4141), .QN(n5614) );
  NAND2X0 U8127 ( .IN1(n4142), .IN2(n5615), .QN(P1_N1616) );
  NAND2X0 U8128 ( .IN1(n7026), .IN2(n4144), .QN(n5615) );
  NAND2X0 U8129 ( .IN1(n4145), .IN2(n5616), .QN(P1_N1615) );
  NAND2X0 U8130 ( .IN1(n7026), .IN2(n4147), .QN(n5616) );
  NAND2X0 U8131 ( .IN1(n4148), .IN2(n5617), .QN(P1_N1614) );
  NAND2X0 U8132 ( .IN1(n7022), .IN2(n4150), .QN(n5617) );
  NAND2X0 U8133 ( .IN1(n4151), .IN2(n5618), .QN(P1_N1613) );
  NAND2X0 U8134 ( .IN1(n7022), .IN2(n4153), .QN(n5618) );
  NAND2X0 U8135 ( .IN1(n4154), .IN2(n5619), .QN(P1_N1612) );
  NAND2X0 U8136 ( .IN1(n7022), .IN2(n4156), .QN(n5619) );
  NAND2X0 U8139 ( .IN1(n5621), .IN2(n5622), .QN(P1_N1568) );
  NAND2X0 U8140 ( .IN1(P1_N1385), .IN2(n5623), .QN(n5622) );
  NAND2X0 U8141 ( .IN1(P1_N392), .IN2(P1_N5573), .QN(n5621) );
  NAND2X0 U8142 ( .IN1(n5625), .IN2(n5626), .QN(P1_N1567) );
  NAND2X0 U8143 ( .IN1(P1_N1384), .IN2(n5623), .QN(n5626) );
  NAND2X0 U8144 ( .IN1(P1_N391), .IN2(P1_N5573), .QN(n5625) );
  NAND2X0 U8145 ( .IN1(n5627), .IN2(n5628), .QN(P1_N1566) );
  NAND2X0 U8146 ( .IN1(P1_N1383), .IN2(n5623), .QN(n5628) );
  NAND2X0 U8147 ( .IN1(P1_N390), .IN2(P1_N5573), .QN(n5627) );
  NAND2X0 U8148 ( .IN1(n5629), .IN2(n5630), .QN(P1_N1565) );
  NAND2X0 U8149 ( .IN1(P1_N1382), .IN2(n5623), .QN(n5630) );
  NAND2X0 U8150 ( .IN1(P1_N389), .IN2(P1_N5573), .QN(n5629) );
  NAND2X0 U8151 ( .IN1(n5631), .IN2(n5632), .QN(P1_N1564) );
  NAND2X0 U8152 ( .IN1(P1_N1381), .IN2(n5623), .QN(n5632) );
  NAND2X0 U8153 ( .IN1(P1_N388), .IN2(P1_N5573), .QN(n5631) );
  NAND2X0 U8154 ( .IN1(n5633), .IN2(n5634), .QN(P1_N1563) );
  NAND2X0 U8155 ( .IN1(P1_N1380), .IN2(n5623), .QN(n5634) );
  NAND2X0 U8156 ( .IN1(P1_N387), .IN2(P1_N5573), .QN(n5633) );
  NAND2X0 U8157 ( .IN1(n5635), .IN2(n5636), .QN(P1_N1562) );
  NAND2X0 U8158 ( .IN1(P1_N1379), .IN2(n5623), .QN(n5636) );
  NAND2X0 U8159 ( .IN1(P1_N386), .IN2(P1_N5573), .QN(n5635) );
  NAND2X0 U8160 ( .IN1(n5637), .IN2(n5638), .QN(P1_N1561) );
  NAND2X0 U8161 ( .IN1(P1_N1378), .IN2(n5623), .QN(n5638) );
  NAND2X0 U8162 ( .IN1(P1_N385), .IN2(P1_N5573), .QN(n5637) );
  NAND2X0 U8163 ( .IN1(n5639), .IN2(n5640), .QN(P1_N1560) );
  NAND2X0 U8164 ( .IN1(P1_N1377), .IN2(n5623), .QN(n5640) );
  NAND2X0 U8165 ( .IN1(P1_N384), .IN2(P1_N5573), .QN(n5639) );
  NAND2X0 U8166 ( .IN1(n5641), .IN2(n5642), .QN(P1_N1559) );
  NAND2X0 U8167 ( .IN1(n5623), .IN2(P1_N1376), .QN(n5642) );
  NAND2X0 U8168 ( .IN1(P1_N383), .IN2(P1_N5573), .QN(n5641) );
  NAND2X0 U8169 ( .IN1(n5643), .IN2(n5644), .QN(P1_N1558) );
  NAND2X0 U8170 ( .IN1(n5623), .IN2(P1_N1375), .QN(n5644) );
  NAND2X0 U8171 ( .IN1(P1_N382), .IN2(P1_N5573), .QN(n5643) );
  NAND2X0 U8172 ( .IN1(n5645), .IN2(n5646), .QN(P1_N1557) );
  NAND2X0 U8173 ( .IN1(n5623), .IN2(P1_N1374), .QN(n5646) );
  NAND2X0 U8174 ( .IN1(P1_N381), .IN2(P1_N5573), .QN(n5645) );
  NAND2X0 U8175 ( .IN1(n5647), .IN2(n5648), .QN(P1_N1556) );
  NAND2X0 U8176 ( .IN1(n5623), .IN2(P1_N1373), .QN(n5648) );
  NAND2X0 U8177 ( .IN1(P1_N380), .IN2(P1_N5573), .QN(n5647) );
  NAND2X0 U8178 ( .IN1(n5649), .IN2(n5650), .QN(P1_N1555) );
  NAND2X0 U8179 ( .IN1(n5623), .IN2(P1_N1372), .QN(n5650) );
  NAND2X0 U8180 ( .IN1(P1_N379), .IN2(P1_N5573), .QN(n5649) );
  NAND2X0 U8181 ( .IN1(n5651), .IN2(n5652), .QN(P1_N1554) );
  NAND2X0 U8182 ( .IN1(n5623), .IN2(P1_N1371), .QN(n5652) );
  NAND2X0 U8183 ( .IN1(P1_N378), .IN2(P1_N5573), .QN(n5651) );
  NAND2X0 U8184 ( .IN1(n5653), .IN2(n5654), .QN(P1_N1553) );
  NAND2X0 U8185 ( .IN1(n5623), .IN2(P1_N1370), .QN(n5654) );
  NAND2X0 U8186 ( .IN1(P1_N377), .IN2(P1_N5573), .QN(n5653) );
  NAND2X0 U8187 ( .IN1(n5655), .IN2(n5656), .QN(P1_N1552) );
  NAND2X0 U8188 ( .IN1(n5623), .IN2(P1_N1369), .QN(n5656) );
  NAND2X0 U8189 ( .IN1(P1_N376), .IN2(P1_N5573), .QN(n5655) );
  NAND2X0 U8190 ( .IN1(n5657), .IN2(n5658), .QN(P1_N1551) );
  NAND2X0 U8191 ( .IN1(n5623), .IN2(P1_N1368), .QN(n5658) );
  NAND2X0 U8192 ( .IN1(P1_N375), .IN2(P1_N5573), .QN(n5657) );
  NAND2X0 U8193 ( .IN1(n5659), .IN2(n5660), .QN(P1_N1550) );
  NAND2X0 U8194 ( .IN1(n5623), .IN2(P1_N1367), .QN(n5660) );
  NAND2X0 U8195 ( .IN1(P1_N374), .IN2(P1_N5573), .QN(n5659) );
  NAND2X0 U8196 ( .IN1(n5661), .IN2(n5662), .QN(P1_N1549) );
  NAND2X0 U8197 ( .IN1(n5623), .IN2(P1_N1366), .QN(n5662) );
  NAND2X0 U8198 ( .IN1(P1_N373), .IN2(P1_N5573), .QN(n5661) );
  NAND2X0 U8199 ( .IN1(n5663), .IN2(n5664), .QN(P1_N1548) );
  NAND2X0 U8200 ( .IN1(n5623), .IN2(P1_N1365), .QN(n5664) );
  NAND2X0 U8201 ( .IN1(P1_N372), .IN2(P1_N5573), .QN(n5663) );
  NAND2X0 U8202 ( .IN1(n5665), .IN2(n5666), .QN(P1_N1547) );
  NAND2X0 U8203 ( .IN1(n5623), .IN2(P1_N1364), .QN(n5666) );
  NAND2X0 U8204 ( .IN1(P1_N371), .IN2(P1_N5573), .QN(n5665) );
  NAND2X0 U8205 ( .IN1(n5667), .IN2(n5668), .QN(P1_N1546) );
  NAND2X0 U8206 ( .IN1(n5623), .IN2(P1_N1363), .QN(n5668) );
  NAND2X0 U8013 ( .IN1(P1_N1865), .IN2(n5511), .QN(n5546) );
  NAND2X0 U8014 ( .IN1(P1_N375), .IN2(P1_N5577), .QN(n5545) );
  NAND2X0 U8015 ( .IN1(n5547), .IN2(n5548), .QN(P1_N1923) );
  NAND2X0 U8016 ( .IN1(P1_N1864), .IN2(n5511), .QN(n5548) );
  NAND2X0 U8017 ( .IN1(P1_N374), .IN2(P1_N5577), .QN(n5547) );
  NAND2X0 U8018 ( .IN1(n5549), .IN2(n5550), .QN(P1_N1922) );
  NAND2X0 U8019 ( .IN1(P1_N1863), .IN2(n5511), .QN(n5550) );
  NAND2X0 U8020 ( .IN1(P1_N373), .IN2(P1_N5577), .QN(n5549) );
  NAND2X0 U8021 ( .IN1(n5551), .IN2(n5552), .QN(P1_N1921) );
  NAND2X0 U8022 ( .IN1(P1_N1862), .IN2(n5511), .QN(n5552) );
  NAND2X0 U8023 ( .IN1(P1_N372), .IN2(P1_N5577), .QN(n5551) );
  NAND2X0 U8024 ( .IN1(n5553), .IN2(n5554), .QN(P1_N1920) );
  NAND2X0 U8025 ( .IN1(P1_N1861), .IN2(n5511), .QN(n5554) );
  NAND2X0 U8026 ( .IN1(P1_N371), .IN2(P1_N5577), .QN(n5553) );
  NAND2X0 U8027 ( .IN1(n5555), .IN2(n5556), .QN(P1_N1919) );
  NAND2X0 U8028 ( .IN1(P1_N1860), .IN2(n5511), .QN(n5556) );
  NAND2X0 U8029 ( .IN1(P1_N370), .IN2(P1_N5577), .QN(n5555) );
  NAND2X0 U8030 ( .IN1(n5557), .IN2(n5558), .QN(P1_N1918) );
  NAND2X0 U8031 ( .IN1(P1_N1859), .IN2(n5511), .QN(n5558) );
  NAND2X0 U8032 ( .IN1(P1_N369), .IN2(P1_N5577), .QN(n5557) );
  NAND2X0 U8033 ( .IN1(n5559), .IN2(n5560), .QN(P1_N1917) );
  NAND2X0 U8034 ( .IN1(P1_N1858), .IN2(n5511), .QN(n5560) );
  NAND2X0 U8035 ( .IN1(P1_N368), .IN2(P1_N5577), .QN(n5559) );
  NAND2X0 U8036 ( .IN1(n5561), .IN2(n5562), .QN(P1_N1916) );
  NAND2X0 U8037 ( .IN1(P1_N1857), .IN2(n5511), .QN(n5562) );
  NAND2X0 U8038 ( .IN1(n18451), .IN2(P1_N5577), .QN(n5561) );
  NAND2X0 U8039 ( .IN1(n5563), .IN2(n5564), .QN(P1_N1915) );
  NAND2X0 U8040 ( .IN1(P1_N1856), .IN2(n5511), .QN(n5564) );
  NAND2X0 U8041 ( .IN1(n6623), .IN2(P1_N5577), .QN(n5563) );
  NAND2X0 U8042 ( .IN1(n5565), .IN2(n5566), .QN(P1_N1914) );
  NAND2X0 U8043 ( .IN1(P1_N1855), .IN2(n5511), .QN(n5566) );
  NAND2X0 U8044 ( .IN1(n6622), .IN2(P1_N5577), .QN(n5565) );
  NAND2X0 U8045 ( .IN1(n5567), .IN2(n5568), .QN(P1_N1913) );
  NAND2X0 U8046 ( .IN1(P1_N1854), .IN2(n5511), .QN(n5568) );
  NAND2X0 U8049 ( .IN1(n6621), .IN2(P1_N5577), .QN(n5567) );
  AND2X1 U8054 ( .IN1(P1_N134), .IN2(n5571), .Q(P1_N190) );
  NAND2X0 U8055 ( .IN1(n5572), .IN2(n5573), .QN(n5571) );
  NOR2X0 U8056 ( .QN(n5573), .IN1(n5574), .IN2(n5575) );
  NAND2X0 U8057 ( .IN1(n5576), .IN2(n5577), .QN(n5575) );
  AND2X1 U8058 ( .IN1(n5578), .IN2(n5579), .Q(n5577) );
  NOR2X0 U8059 ( .QN(n5579), .IN1(P1_N156), .IN2(P1_N155) );
  NOR2X0 U8060 ( .QN(n5578), .IN1(P1_N154), .IN2(P1_N153) );
  NOR2X0 U8061 ( .QN(n5576), .IN1(P1_N150), .IN2(n5580) );
  OR2X1 U8062 ( .IN2(P1_N151), .IN1(P1_N152), .Q(n5580) );
  NAND2X0 U8063 ( .IN1(n5581), .IN2(n5582), .QN(n5574) );
  AND2X1 U8064 ( .IN1(n5583), .IN2(n5584), .Q(n5582) );
  NOR2X0 U8065 ( .QN(n5584), .IN1(P1_N163), .IN2(P1_N162) );
  NOR2X0 U8066 ( .QN(n5583), .IN1(P1_N161), .IN2(P1_N160) );
  NOR2X0 U8067 ( .QN(n5581), .IN1(P1_N157), .IN2(n5585) );
  OR2X1 U8068 ( .IN2(P1_N158), .IN1(P1_N159), .Q(n5585) );
  NOR2X0 U8069 ( .QN(n5572), .IN1(n5586), .IN2(n5587) );
  NAND2X0 U8070 ( .IN1(n5588), .IN2(n5589), .QN(n5587) );
  NOR2X0 U8071 ( .QN(n5589), .IN1(P1_N140), .IN2(n5590) );
  OR2X1 U8072 ( .IN2(P1_N141), .IN1(P1_N142), .Q(n5590) );
  NOR2X0 U8073 ( .QN(n5588), .IN1(P1_N137), .IN2(n5591) );
  OR2X1 U8074 ( .IN2(P1_N138), .IN1(P1_N139), .Q(n5591) );
  NAND2X0 U8075 ( .IN1(n5592), .IN2(n5593), .QN(n5586) );
  AND2X1 U8076 ( .IN1(n5594), .IN2(n5595), .Q(n5593) );
  NOR2X0 U8077 ( .QN(n5595), .IN1(P1_N149), .IN2(P1_N148) );
  NOR2X0 U8078 ( .QN(n5594), .IN1(P1_N147), .IN2(P1_N146) );
  NOR2X0 U8079 ( .QN(n5592), .IN1(P1_N143), .IN2(n5596) );
  OR2X1 U8080 ( .IN2(P1_N144), .IN1(P1_N145), .Q(n5596) );
  NAND2X0 U8081 ( .IN1(n7360), .IN2(n5597), .QN(P1_N1761) );
  NAND2X0 U8082 ( .IN1(n7359), .IN2(n5598), .QN(P1_N1759) );
  NOR2X0 U8083 ( .QN(P1_N1942), .IN1(n5598), .IN2(n5597) );
  INVX0 U8084 ( .ZN(n5597), .INP(n7359) );
  INVX0 U8085 ( .ZN(n5598), .INP(n7360) );
  NOR2X0 U8086 ( .QN(P1_N1641), .IN1(n7328), .IN2(n7023) );
  NOR2X0 U8087 ( .QN(P1_N1640), .IN1(n7326), .IN2(n7023) );
  NOR2X0 U8088 ( .QN(P1_N1639), .IN1(n7324), .IN2(n7021) );
  NOR2X0 U8089 ( .QN(P1_N1638), .IN1(n7322), .IN2(n7021) );
  NOR2X0 U8090 ( .QN(P1_N1637), .IN1(n7320), .IN2(n7021) );
  NOR2X0 U8091 ( .QN(P1_N1636), .IN1(n7318), .IN2(n7021) );
  NOR2X0 U8092 ( .QN(P1_N1635), .IN1(n7316), .IN2(n7029) );
  NOR2X0 U8093 ( .QN(P1_N1634), .IN1(n7314), .IN2(n7027) );
  NOR2X0 U8094 ( .QN(P1_N1633), .IN1(n7312), .IN2(n7027) );
  NOR2X0 U8095 ( .QN(P1_N1632), .IN1(n7310), .IN2(n7029) );
  NAND2X0 U8097 ( .IN1(n4097), .IN2(n5600), .QN(P1_N1631) );
  NAND2X0 U8098 ( .IN1(n7019), .IN2(n4099), .QN(n5600) );
  NAND2X0 U8099 ( .IN1(n4100), .IN2(n5601), .QN(P1_N1630) );
  NAND2X0 U8100 ( .IN1(n7019), .IN2(n4102), .QN(n5601) );
  NAND2X0 U8101 ( .IN1(n4103), .IN2(n5602), .QN(P1_N1629) );
  NAND2X0 U8102 ( .IN1(n7028), .IN2(n4105), .QN(n5602) );
  NAND2X0 U8103 ( .IN1(n4106), .IN2(n5603), .QN(P1_N1628) );
  NAND2X0 U8104 ( .IN1(n7028), .IN2(n4108), .QN(n5603) );
  NAND2X0 U8105 ( .IN1(n4109), .IN2(n5604), .QN(P1_N1627) );
  NAND2X0 U8106 ( .IN1(n7028), .IN2(n4111), .QN(n5604) );
  NAND2X0 U8107 ( .IN1(n4112), .IN2(n5605), .QN(P1_N1626) );
  NAND2X0 U8108 ( .IN1(n7024), .IN2(n4114), .QN(n5605) );
  NAND2X0 U8109 ( .IN1(n4115), .IN2(n5606), .QN(P1_N1625) );
  NAND2X0 U8110 ( .IN1(n7024), .IN2(n4117), .QN(n5606) );
  NAND2X0 U8111 ( .IN1(n4118), .IN2(n5607), .QN(P1_N1624) );
  NOR2X0 U7917 ( .QN(P1_N2005), .IN1(n7310), .IN2(n7021) );
  NAND2X0 U7919 ( .IN1(n4097), .IN2(n5488), .QN(P1_N2004) );
  NAND2X0 U7920 ( .IN1(n7019), .IN2(n4099), .QN(n5488) );
  NAND2X0 U7921 ( .IN1(n4100), .IN2(n5489), .QN(P1_N2003) );
  NAND2X0 U7922 ( .IN1(n7028), .IN2(n4102), .QN(n5489) );
  NAND2X0 U7923 ( .IN1(n4103), .IN2(n5490), .QN(P1_N2002) );
  NAND2X0 U7924 ( .IN1(n7028), .IN2(n4105), .QN(n5490) );
  NAND2X0 U7925 ( .IN1(n4106), .IN2(n5491), .QN(P1_N2001) );
  NAND2X0 U7926 ( .IN1(n7028), .IN2(n4108), .QN(n5491) );
  NAND2X0 U7927 ( .IN1(n4109), .IN2(n5492), .QN(P1_N2000) );
  NAND2X0 U7928 ( .IN1(n7028), .IN2(n4111), .QN(n5492) );
  NAND2X0 U7929 ( .IN1(n4112), .IN2(n5493), .QN(P1_N1999) );
  NAND2X0 U7930 ( .IN1(n7024), .IN2(n4114), .QN(n5493) );
  NAND2X0 U7931 ( .IN1(n4115), .IN2(n5494), .QN(P1_N1998) );
  NAND2X0 U7932 ( .IN1(n7024), .IN2(n4117), .QN(n5494) );
  NAND2X0 U7933 ( .IN1(n4118), .IN2(n5495), .QN(P1_N1997) );
  NAND2X0 U7934 ( .IN1(n7024), .IN2(n4120), .QN(n5495) );
  NAND2X0 U7935 ( .IN1(n4121), .IN2(n5496), .QN(P1_N1996) );
  NAND2X0 U7936 ( .IN1(n7024), .IN2(n4123), .QN(n5496) );
  NAND2X0 U7937 ( .IN1(n4124), .IN2(n5497), .QN(P1_N1995) );
  NAND2X0 U7938 ( .IN1(n7024), .IN2(n4126), .QN(n5497) );
  NAND2X0 U7939 ( .IN1(n4127), .IN2(n5498), .QN(P1_N1994) );
  NAND2X0 U7940 ( .IN1(n7463), .IN2(n4129), .QN(n5498) );
  NAND2X0 U7941 ( .IN1(n4130), .IN2(n5499), .QN(P1_N1993) );
  NAND2X0 U7942 ( .IN1(n7463), .IN2(n4132), .QN(n5499) );
  NAND2X0 U7943 ( .IN1(n4133), .IN2(n5500), .QN(P1_N1992) );
  NAND2X0 U7944 ( .IN1(n7463), .IN2(n4135), .QN(n5500) );
  NAND2X0 U7945 ( .IN1(n4136), .IN2(n5501), .QN(P1_N1991) );
  NAND2X0 U7946 ( .IN1(n7463), .IN2(n4138), .QN(n5501) );
  NAND2X0 U7947 ( .IN1(n4139), .IN2(n5502), .QN(P1_N1990) );
  NAND2X0 U7948 ( .IN1(n7026), .IN2(n4141), .QN(n5502) );
  NAND2X0 U7949 ( .IN1(n4142), .IN2(n5503), .QN(P1_N1989) );
  NAND2X0 U7950 ( .IN1(n7026), .IN2(n4144), .QN(n5503) );
  NAND2X0 U7951 ( .IN1(n4145), .IN2(n5504), .QN(P1_N1988) );
  NAND2X0 U7952 ( .IN1(n7026), .IN2(n4147), .QN(n5504) );
  NAND2X0 U7953 ( .IN1(n4148), .IN2(n5505), .QN(P1_N1987) );
  NAND2X0 U7954 ( .IN1(n7022), .IN2(n4150), .QN(n5505) );
  NAND2X0 U7955 ( .IN1(n4151), .IN2(n5506), .QN(P1_N1986) );
  NAND2X0 U7956 ( .IN1(n7022), .IN2(n4153), .QN(n5506) );
  NAND2X0 U7957 ( .IN1(n4154), .IN2(n5507), .QN(P1_N1985) );
  NAND2X0 U7958 ( .IN1(n7022), .IN2(n4156), .QN(n5507) );
  NAND2X0 U7961 ( .IN1(n5509), .IN2(n5510), .QN(P1_N1941) );
  NAND2X0 U7962 ( .IN1(P1_N1882), .IN2(n5511), .QN(n5510) );
  NAND2X0 U7963 ( .IN1(P1_N392), .IN2(P1_N5577), .QN(n5509) );
  NAND2X0 U7964 ( .IN1(n5513), .IN2(n5514), .QN(P1_N1940) );
  NAND2X0 U7965 ( .IN1(P1_N1881), .IN2(n5511), .QN(n5514) );
  NAND2X0 U7966 ( .IN1(P1_N391), .IN2(P1_N5577), .QN(n5513) );
  NAND2X0 U7967 ( .IN1(n5515), .IN2(n5516), .QN(P1_N1939) );
  NAND2X0 U7968 ( .IN1(P1_N1880), .IN2(n5511), .QN(n5516) );
  NAND2X0 U7969 ( .IN1(P1_N390), .IN2(P1_N5577), .QN(n5515) );
  NAND2X0 U7970 ( .IN1(n5517), .IN2(n5518), .QN(P1_N1938) );
  NAND2X0 U7971 ( .IN1(P1_N1879), .IN2(n5511), .QN(n5518) );
  NAND2X0 U7972 ( .IN1(P1_N389), .IN2(P1_N5577), .QN(n5517) );
  NAND2X0 U7973 ( .IN1(n5519), .IN2(n5520), .QN(P1_N1937) );
  NAND2X0 U7974 ( .IN1(P1_N1878), .IN2(n5511), .QN(n5520) );
  NAND2X0 U7975 ( .IN1(P1_N388), .IN2(P1_N5577), .QN(n5519) );
  NAND2X0 U7976 ( .IN1(n5521), .IN2(n5522), .QN(P1_N1936) );
  NAND2X0 U7977 ( .IN1(P1_N1877), .IN2(n5511), .QN(n5522) );
  NAND2X0 U7978 ( .IN1(P1_N387), .IN2(P1_N5577), .QN(n5521) );
  NAND2X0 U7979 ( .IN1(n5523), .IN2(n5524), .QN(P1_N1935) );
  NAND2X0 U7980 ( .IN1(P1_N1876), .IN2(n5511), .QN(n5524) );
  NAND2X0 U7981 ( .IN1(P1_N386), .IN2(P1_N5577), .QN(n5523) );
  NAND2X0 U7982 ( .IN1(n5525), .IN2(n5526), .QN(P1_N1934) );
  NAND2X0 U7983 ( .IN1(P1_N1875), .IN2(n5511), .QN(n5526) );
  NAND2X0 U7984 ( .IN1(P1_N385), .IN2(P1_N5577), .QN(n5525) );
  NAND2X0 U7985 ( .IN1(n5527), .IN2(n5528), .QN(P1_N1933) );
  NAND2X0 U7986 ( .IN1(P1_N1874), .IN2(n5511), .QN(n5528) );
  NAND2X0 U7987 ( .IN1(P1_N384), .IN2(P1_N5577), .QN(n5527) );
  NAND2X0 U7988 ( .IN1(n5529), .IN2(n5530), .QN(P1_N1932) );
  NAND2X0 U7989 ( .IN1(P1_N1873), .IN2(n5511), .QN(n5530) );
  NAND2X0 U7990 ( .IN1(P1_N383), .IN2(P1_N5577), .QN(n5529) );
  NAND2X0 U7991 ( .IN1(n5531), .IN2(n5532), .QN(P1_N1931) );
  NAND2X0 U7992 ( .IN1(P1_N1872), .IN2(n5511), .QN(n5532) );
  NAND2X0 U7993 ( .IN1(P1_N382), .IN2(P1_N5577), .QN(n5531) );
  NAND2X0 U7994 ( .IN1(n5533), .IN2(n5534), .QN(P1_N1930) );
  NAND2X0 U7995 ( .IN1(P1_N1871), .IN2(n5511), .QN(n5534) );
  NAND2X0 U7996 ( .IN1(P1_N381), .IN2(P1_N5577), .QN(n5533) );
  NAND2X0 U7997 ( .IN1(n5535), .IN2(n5536), .QN(P1_N1929) );
  NAND2X0 U7998 ( .IN1(P1_N1870), .IN2(n5511), .QN(n5536) );
  NAND2X0 U7999 ( .IN1(P1_N380), .IN2(P1_N5577), .QN(n5535) );
  NAND2X0 U8000 ( .IN1(n5537), .IN2(n5538), .QN(P1_N1928) );
  NAND2X0 U8001 ( .IN1(P1_N1869), .IN2(n5511), .QN(n5538) );
  NAND2X0 U8002 ( .IN1(P1_N379), .IN2(P1_N5577), .QN(n5537) );
  NAND2X0 U8003 ( .IN1(n5539), .IN2(n5540), .QN(P1_N1927) );
  NAND2X0 U8004 ( .IN1(P1_N1868), .IN2(n5511), .QN(n5540) );
  NAND2X0 U8005 ( .IN1(P1_N378), .IN2(P1_N5577), .QN(n5539) );
  NAND2X0 U8006 ( .IN1(n5541), .IN2(n5542), .QN(P1_N1926) );
  NAND2X0 U8007 ( .IN1(P1_N1867), .IN2(n5511), .QN(n5542) );
  NAND2X0 U8008 ( .IN1(P1_N377), .IN2(P1_N5577), .QN(n5541) );
  NAND2X0 U8009 ( .IN1(n5543), .IN2(n5544), .QN(P1_N1925) );
  NAND2X0 U8010 ( .IN1(P1_N1866), .IN2(n5511), .QN(n5544) );
  NAND2X0 U8011 ( .IN1(P1_N376), .IN2(P1_N5577), .QN(n5543) );
  NAND2X0 U8012 ( .IN1(n5545), .IN2(n5546), .QN(P1_N1924) );
  NAND2X0 U7819 ( .IN1(n5431), .IN2(n5432), .QN(P1_N2311) );
  NAND2X0 U7820 ( .IN1(P1_N2252), .IN2(n5425), .QN(n5432) );
  NAND2X0 U7821 ( .IN1(P1_N389), .IN2(P1_N5578), .QN(n5431) );
  NAND2X0 U7822 ( .IN1(n5433), .IN2(n5434), .QN(P1_N2310) );
  NAND2X0 U7823 ( .IN1(P1_N2251), .IN2(n5425), .QN(n5434) );
  NAND2X0 U7824 ( .IN1(P1_N388), .IN2(P1_N5578), .QN(n5433) );
  NAND2X0 U7825 ( .IN1(n5435), .IN2(n5436), .QN(P1_N2309) );
  NAND2X0 U7826 ( .IN1(P1_N2250), .IN2(n5425), .QN(n5436) );
  NAND2X0 U7827 ( .IN1(P1_N387), .IN2(P1_N5578), .QN(n5435) );
  NAND2X0 U7828 ( .IN1(n5437), .IN2(n5438), .QN(P1_N2308) );
  NAND2X0 U7829 ( .IN1(P1_N2249), .IN2(n5425), .QN(n5438) );
  NAND2X0 U7830 ( .IN1(P1_N386), .IN2(P1_N5578), .QN(n5437) );
  NAND2X0 U7831 ( .IN1(n5439), .IN2(n5440), .QN(P1_N2307) );
  NAND2X0 U7832 ( .IN1(P1_N2248), .IN2(n5425), .QN(n5440) );
  NAND2X0 U7833 ( .IN1(P1_N385), .IN2(P1_N5578), .QN(n5439) );
  NAND2X0 U7834 ( .IN1(n5441), .IN2(n5442), .QN(P1_N2306) );
  NAND2X0 U7835 ( .IN1(P1_N2247), .IN2(n5425), .QN(n5442) );
  NAND2X0 U7836 ( .IN1(P1_N384), .IN2(P1_N5578), .QN(n5441) );
  NAND2X0 U7837 ( .IN1(n5443), .IN2(n5444), .QN(P1_N2305) );
  NAND2X0 U7838 ( .IN1(P1_N2246), .IN2(n5425), .QN(n5444) );
  NAND2X0 U7839 ( .IN1(P1_N383), .IN2(P1_N5578), .QN(n5443) );
  NAND2X0 U7840 ( .IN1(n5445), .IN2(n5446), .QN(P1_N2304) );
  NAND2X0 U7841 ( .IN1(P1_N2245), .IN2(n5425), .QN(n5446) );
  NAND2X0 U7842 ( .IN1(P1_N382), .IN2(P1_N5578), .QN(n5445) );
  NAND2X0 U7843 ( .IN1(n5447), .IN2(n5448), .QN(P1_N2303) );
  NAND2X0 U7844 ( .IN1(P1_N2244), .IN2(n5425), .QN(n5448) );
  NAND2X0 U7845 ( .IN1(P1_N381), .IN2(P1_N5578), .QN(n5447) );
  NAND2X0 U7846 ( .IN1(n5449), .IN2(n5450), .QN(P1_N2302) );
  NAND2X0 U7847 ( .IN1(P1_N2243), .IN2(n5425), .QN(n5450) );
  NAND2X0 U7848 ( .IN1(P1_N380), .IN2(P1_N5578), .QN(n5449) );
  NAND2X0 U7849 ( .IN1(n5451), .IN2(n5452), .QN(P1_N2301) );
  NAND2X0 U7850 ( .IN1(P1_N2242), .IN2(n5425), .QN(n5452) );
  NAND2X0 U7851 ( .IN1(P1_N379), .IN2(P1_N5578), .QN(n5451) );
  NAND2X0 U7852 ( .IN1(n5453), .IN2(n5454), .QN(P1_N2300) );
  NAND2X0 U7853 ( .IN1(P1_N2241), .IN2(n5425), .QN(n5454) );
  NAND2X0 U7854 ( .IN1(P1_N378), .IN2(P1_N5578), .QN(n5453) );
  NAND2X0 U7855 ( .IN1(n5455), .IN2(n5456), .QN(P1_N2299) );
  NAND2X0 U7856 ( .IN1(P1_N2240), .IN2(n5425), .QN(n5456) );
  NAND2X0 U7857 ( .IN1(P1_N377), .IN2(P1_N5578), .QN(n5455) );
  NAND2X0 U7858 ( .IN1(n5457), .IN2(n5458), .QN(P1_N2298) );
  NAND2X0 U7859 ( .IN1(P1_N2239), .IN2(n5425), .QN(n5458) );
  NAND2X0 U7860 ( .IN1(P1_N376), .IN2(P1_N5578), .QN(n5457) );
  NAND2X0 U7861 ( .IN1(n5459), .IN2(n5460), .QN(P1_N2297) );
  NAND2X0 U7862 ( .IN1(P1_N2238), .IN2(n5425), .QN(n5460) );
  NAND2X0 U7863 ( .IN1(P1_N375), .IN2(P1_N5578), .QN(n5459) );
  NAND2X0 U7864 ( .IN1(n5461), .IN2(n5462), .QN(P1_N2296) );
  NAND2X0 U7865 ( .IN1(P1_N2237), .IN2(n5425), .QN(n5462) );
  NAND2X0 U7866 ( .IN1(P1_N374), .IN2(P1_N5578), .QN(n5461) );
  NAND2X0 U7867 ( .IN1(n5463), .IN2(n5464), .QN(P1_N2295) );
  NAND2X0 U7868 ( .IN1(P1_N2236), .IN2(n5425), .QN(n5464) );
  NAND2X0 U7869 ( .IN1(P1_N373), .IN2(P1_N5578), .QN(n5463) );
  NAND2X0 U7870 ( .IN1(n5465), .IN2(n5466), .QN(P1_N2294) );
  NAND2X0 U7871 ( .IN1(P1_N2235), .IN2(n5425), .QN(n5466) );
  NAND2X0 U7872 ( .IN1(P1_N372), .IN2(P1_N5578), .QN(n5465) );
  NAND2X0 U7873 ( .IN1(n5467), .IN2(n5468), .QN(P1_N2293) );
  NAND2X0 U7874 ( .IN1(P1_N2234), .IN2(n5425), .QN(n5468) );
  NAND2X0 U7875 ( .IN1(P1_N371), .IN2(P1_N5578), .QN(n5467) );
  NAND2X0 U7876 ( .IN1(n5469), .IN2(n5470), .QN(P1_N2292) );
  NAND2X0 U7877 ( .IN1(P1_N2233), .IN2(n5425), .QN(n5470) );
  NAND2X0 U7878 ( .IN1(P1_N370), .IN2(P1_N5578), .QN(n5469) );
  NAND2X0 U7879 ( .IN1(n5471), .IN2(n5472), .QN(P1_N2291) );
  NAND2X0 U7880 ( .IN1(P1_N2232), .IN2(n5425), .QN(n5472) );
  NAND2X0 U7881 ( .IN1(P1_N369), .IN2(P1_N5578), .QN(n5471) );
  NAND2X0 U7882 ( .IN1(n5473), .IN2(n5474), .QN(P1_N2290) );
  NAND2X0 U7883 ( .IN1(P1_N2231), .IN2(n5425), .QN(n5474) );
  NAND2X0 U7884 ( .IN1(P1_N368), .IN2(P1_N5578), .QN(n5473) );
  NAND2X0 U7885 ( .IN1(n5475), .IN2(n5476), .QN(P1_N2289) );
  NAND2X0 U7886 ( .IN1(P1_N2230), .IN2(n5425), .QN(n5476) );
  NAND2X0 U7887 ( .IN1(n18451), .IN2(P1_N5578), .QN(n5475) );
  NAND2X0 U7888 ( .IN1(n5477), .IN2(n5478), .QN(P1_N2288) );
  NAND2X0 U7889 ( .IN1(P1_N2229), .IN2(n5425), .QN(n5478) );
  NAND2X0 U7890 ( .IN1(n6623), .IN2(P1_N5578), .QN(n5477) );
  NAND2X0 U7891 ( .IN1(n5479), .IN2(n5480), .QN(P1_N2287) );
  NAND2X0 U7892 ( .IN1(P1_N2228), .IN2(n5425), .QN(n5480) );
  NAND2X0 U7893 ( .IN1(n6622), .IN2(P1_N5578), .QN(n5479) );
  NAND2X0 U7894 ( .IN1(n5481), .IN2(n5482), .QN(P1_N2286) );
  NAND2X0 U7895 ( .IN1(P1_N2227), .IN2(n5425), .QN(n5482) );
  NAND2X0 U7898 ( .IN1(n6621), .IN2(P1_N5578), .QN(n5481) );
  NAND2X0 U7903 ( .IN1(n7362), .IN2(n5485), .QN(P1_N2134) );
  NAND2X0 U7904 ( .IN1(n7361), .IN2(n5486), .QN(P1_N2132) );
  NOR2X0 U7905 ( .QN(P1_N2315), .IN1(n5486), .IN2(n5485) );
  INVX0 U7906 ( .ZN(n5485), .INP(n7361) );
  INVX0 U7907 ( .ZN(n5486), .INP(n7362) );
  NOR2X0 U7908 ( .QN(P1_N2014), .IN1(n7328), .IN2(n7023) );
  NOR2X0 U7909 ( .QN(P1_N2013), .IN1(n7326), .IN2(n7023) );
  NOR2X0 U7910 ( .QN(P1_N2012), .IN1(n7324), .IN2(n7021) );
  NOR2X0 U7911 ( .QN(P1_N2011), .IN1(n7322), .IN2(n7021) );
  NOR2X0 U7912 ( .QN(P1_N2010), .IN1(n7320), .IN2(n7021) );
  NOR2X0 U7913 ( .QN(P1_N2009), .IN1(n7318), .IN2(n7021) );
  NOR2X0 U7914 ( .QN(P1_N2008), .IN1(n7316), .IN2(n7029) );
  NOR2X0 U7915 ( .QN(P1_N2007), .IN1(n7314), .IN2(n7027) );
  NOR2X0 U7916 ( .QN(P1_N2006), .IN1(n7312), .IN2(n7027) );
  NAND2X0 U7718 ( .IN1(n6622), .IN2(P1_N5579), .QN(n5370) );
  NAND2X0 U7719 ( .IN1(n5372), .IN2(n5373), .QN(P1_N2659) );
  NAND2X0 U7720 ( .IN1(P1_N2600), .IN2(n5316), .QN(n5373) );
  NAND2X0 U7723 ( .IN1(n6621), .IN2(P1_N5579), .QN(n5372) );
  NAND2X0 U7728 ( .IN1(n7364), .IN2(n5376), .QN(P1_N2507) );
  NAND2X0 U7729 ( .IN1(n7363), .IN2(n5377), .QN(P1_N2505) );
  NOR2X0 U7730 ( .QN(P1_N2688), .IN1(n5377), .IN2(n5376) );
  INVX0 U7731 ( .ZN(n5376), .INP(n7363) );
  INVX0 U7732 ( .ZN(n5377), .INP(n7364) );
  AND2X1 U7733 ( .IN1(P1_N193), .IN2(n5378), .Q(P1_N244) );
  NAND2X0 U7734 ( .IN1(n5379), .IN2(n5380), .QN(n5378) );
  NOR2X0 U7735 ( .QN(n5380), .IN1(n5381), .IN2(n5382) );
  NAND2X0 U7736 ( .IN1(n5383), .IN2(n5384), .QN(n5382) );
  NOR2X0 U7737 ( .QN(n5384), .IN1(P1_N212), .IN2(n5385) );
  OR2X1 U7738 ( .IN2(P1_N213), .IN1(P1_N214), .Q(n5385) );
  NOR2X0 U7739 ( .QN(n5383), .IN1(P1_N209), .IN2(n5386) );
  OR2X1 U7740 ( .IN2(P1_N210), .IN1(P1_N211), .Q(n5386) );
  NAND2X0 U7741 ( .IN1(n5387), .IN2(n5388), .QN(n5381) );
  NOR2X0 U7742 ( .QN(n5388), .IN1(P1_N218), .IN2(n5389) );
  OR2X1 U7743 ( .IN2(P1_N219), .IN1(P1_N220), .Q(n5389) );
  NOR2X0 U7744 ( .QN(n5387), .IN1(P1_N215), .IN2(n5390) );
  OR2X1 U7745 ( .IN2(P1_N216), .IN1(P1_N217), .Q(n5390) );
  NOR2X0 U7746 ( .QN(n5379), .IN1(n5391), .IN2(n5392) );
  NAND2X0 U7747 ( .IN1(n5393), .IN2(n5394), .QN(n5392) );
  NOR2X0 U7748 ( .QN(n5394), .IN1(P1_N200), .IN2(n5395) );
  OR2X1 U7749 ( .IN2(P1_N201), .IN1(P1_N202), .Q(n5395) );
  NOR2X0 U7750 ( .QN(n5393), .IN1(P1_N197), .IN2(n5396) );
  OR2X1 U7751 ( .IN2(P1_N198), .IN1(P1_N199), .Q(n5396) );
  NAND2X0 U7752 ( .IN1(n5397), .IN2(n5398), .QN(n5391) );
  NOR2X0 U7753 ( .QN(n5398), .IN1(P1_N206), .IN2(n5399) );
  OR2X1 U7754 ( .IN2(P1_N207), .IN1(P1_N208), .Q(n5399) );
  NOR2X0 U7755 ( .QN(n5397), .IN1(P1_N203), .IN2(n5400) );
  OR2X1 U7756 ( .IN2(P1_N204), .IN1(P1_N205), .Q(n5400) );
  NOR2X0 U7757 ( .QN(P1_N2387), .IN1(n7328), .IN2(n7023) );
  NOR2X0 U7758 ( .QN(P1_N2386), .IN1(n7326), .IN2(n7023) );
  NOR2X0 U7759 ( .QN(P1_N2385), .IN1(n7324), .IN2(n7021) );
  NOR2X0 U7760 ( .QN(P1_N2384), .IN1(n7322), .IN2(n7021) );
  NOR2X0 U7761 ( .QN(P1_N2383), .IN1(n7320), .IN2(n7021) );
  NOR2X0 U7762 ( .QN(P1_N2382), .IN1(n7318), .IN2(n7021) );
  NOR2X0 U7763 ( .QN(P1_N2381), .IN1(n7316), .IN2(n7029) );
  NOR2X0 U7764 ( .QN(P1_N2380), .IN1(n7314), .IN2(n7027) );
  NOR2X0 U7765 ( .QN(P1_N2379), .IN1(n7312), .IN2(n7027) );
  NOR2X0 U7766 ( .QN(P1_N2378), .IN1(n7310), .IN2(n7027) );
  NAND2X0 U7768 ( .IN1(n4097), .IN2(n5402), .QN(P1_N2377) );
  NAND2X0 U7769 ( .IN1(n7019), .IN2(n4099), .QN(n5402) );
  NAND2X0 U7770 ( .IN1(n4100), .IN2(n5403), .QN(P1_N2376) );
  NAND2X0 U7771 ( .IN1(n7019), .IN2(n4102), .QN(n5403) );
  NAND2X0 U7772 ( .IN1(n4103), .IN2(n5404), .QN(P1_N2375) );
  NAND2X0 U7773 ( .IN1(n7028), .IN2(n4105), .QN(n5404) );
  NAND2X0 U7774 ( .IN1(n4106), .IN2(n5405), .QN(P1_N2374) );
  NAND2X0 U7775 ( .IN1(n7028), .IN2(n4108), .QN(n5405) );
  NAND2X0 U7776 ( .IN1(n4109), .IN2(n5406), .QN(P1_N2373) );
  NAND2X0 U7777 ( .IN1(n7028), .IN2(n4111), .QN(n5406) );
  NAND2X0 U7778 ( .IN1(n4112), .IN2(n5407), .QN(P1_N2372) );
  NAND2X0 U7779 ( .IN1(n7024), .IN2(n4114), .QN(n5407) );
  NAND2X0 U7780 ( .IN1(n4115), .IN2(n5408), .QN(P1_N2371) );
  NAND2X0 U7781 ( .IN1(n7024), .IN2(n4117), .QN(n5408) );
  NAND2X0 U7782 ( .IN1(n4118), .IN2(n5409), .QN(P1_N2370) );
  NAND2X0 U7783 ( .IN1(n7024), .IN2(n4120), .QN(n5409) );
  NAND2X0 U7784 ( .IN1(n4121), .IN2(n5410), .QN(P1_N2369) );
  NAND2X0 U7785 ( .IN1(n7024), .IN2(n4123), .QN(n5410) );
  NAND2X0 U7786 ( .IN1(n4124), .IN2(n5411), .QN(P1_N2368) );
  NAND2X0 U7787 ( .IN1(n7024), .IN2(n4126), .QN(n5411) );
  NAND2X0 U7788 ( .IN1(n4127), .IN2(n5412), .QN(P1_N2367) );
  NAND2X0 U7789 ( .IN1(n7463), .IN2(n4129), .QN(n5412) );
  NAND2X0 U7790 ( .IN1(n4130), .IN2(n5413), .QN(P1_N2366) );
  NAND2X0 U7791 ( .IN1(n7463), .IN2(n4132), .QN(n5413) );
  NAND2X0 U7792 ( .IN1(n4133), .IN2(n5414), .QN(P1_N2365) );
  NAND2X0 U7793 ( .IN1(n7463), .IN2(n4135), .QN(n5414) );
  NAND2X0 U7794 ( .IN1(n4136), .IN2(n5415), .QN(P1_N2364) );
  NAND2X0 U7795 ( .IN1(n7463), .IN2(n4138), .QN(n5415) );
  NAND2X0 U7796 ( .IN1(n4139), .IN2(n5416), .QN(P1_N2363) );
  NAND2X0 U7797 ( .IN1(n7026), .IN2(n4141), .QN(n5416) );
  NAND2X0 U7798 ( .IN1(n4142), .IN2(n5417), .QN(P1_N2362) );
  NAND2X0 U7799 ( .IN1(n7026), .IN2(n4144), .QN(n5417) );
  NAND2X0 U7800 ( .IN1(n4145), .IN2(n5418), .QN(P1_N2361) );
  NAND2X0 U7801 ( .IN1(n7026), .IN2(n4147), .QN(n5418) );
  NAND2X0 U7802 ( .IN1(n4148), .IN2(n5419), .QN(P1_N2360) );
  NAND2X0 U7803 ( .IN1(n7022), .IN2(n4150), .QN(n5419) );
  NAND2X0 U7804 ( .IN1(n4151), .IN2(n5420), .QN(P1_N2359) );
  NAND2X0 U7805 ( .IN1(n7022), .IN2(n4153), .QN(n5420) );
  NAND2X0 U7806 ( .IN1(n4154), .IN2(n5421), .QN(P1_N2358) );
  NAND2X0 U7807 ( .IN1(n7022), .IN2(n4156), .QN(n5421) );
  NAND2X0 U7810 ( .IN1(n5423), .IN2(n5424), .QN(P1_N2314) );
  NAND2X0 U7811 ( .IN1(P1_N2255), .IN2(n5425), .QN(n5424) );
  NAND2X0 U7812 ( .IN1(P1_N392), .IN2(P1_N5578), .QN(n5423) );
  NAND2X0 U7813 ( .IN1(n5427), .IN2(n5428), .QN(P1_N2313) );
  NAND2X0 U7814 ( .IN1(P1_N2254), .IN2(n5425), .QN(n5428) );
  NAND2X0 U7815 ( .IN1(P1_N391), .IN2(P1_N5578), .QN(n5427) );
  NAND2X0 U7816 ( .IN1(n5429), .IN2(n5430), .QN(P1_N2312) );
  NAND2X0 U7817 ( .IN1(P1_N2253), .IN2(n5425), .QN(n5430) );
  NAND2X0 U7818 ( .IN1(P1_N390), .IN2(P1_N5578), .QN(n5429) );
  NAND2X0 U7623 ( .IN1(n4142), .IN2(n5308), .QN(P1_N2735) );
  NAND2X0 U7624 ( .IN1(n7026), .IN2(n4144), .QN(n5308) );
  NAND2X0 U7625 ( .IN1(n4145), .IN2(n5309), .QN(P1_N2734) );
  NAND2X0 U7626 ( .IN1(n7026), .IN2(n4147), .QN(n5309) );
  NAND2X0 U7627 ( .IN1(n4148), .IN2(n5310), .QN(P1_N2733) );
  NAND2X0 U7628 ( .IN1(n7022), .IN2(n4150), .QN(n5310) );
  NAND2X0 U7629 ( .IN1(n4151), .IN2(n5311), .QN(P1_N2732) );
  NAND2X0 U7630 ( .IN1(n7022), .IN2(n4153), .QN(n5311) );
  NAND2X0 U7631 ( .IN1(n4154), .IN2(n5312), .QN(P1_N2731) );
  NAND2X0 U7632 ( .IN1(n7022), .IN2(n4156), .QN(n5312) );
  NAND2X0 U7635 ( .IN1(n5314), .IN2(n5315), .QN(P1_N2687) );
  NAND2X0 U7636 ( .IN1(P1_N2628), .IN2(n5316), .QN(n5315) );
  NAND2X0 U7637 ( .IN1(P1_N392), .IN2(P1_N5579), .QN(n5314) );
  NAND2X0 U7638 ( .IN1(n5318), .IN2(n5319), .QN(P1_N2686) );
  NAND2X0 U7639 ( .IN1(P1_N2627), .IN2(n5316), .QN(n5319) );
  NAND2X0 U7640 ( .IN1(P1_N391), .IN2(P1_N5579), .QN(n5318) );
  NAND2X0 U7641 ( .IN1(n5320), .IN2(n5321), .QN(P1_N2685) );
  NAND2X0 U7642 ( .IN1(P1_N2626), .IN2(n5316), .QN(n5321) );
  NAND2X0 U7643 ( .IN1(P1_N390), .IN2(P1_N5579), .QN(n5320) );
  NAND2X0 U7644 ( .IN1(n5322), .IN2(n5323), .QN(P1_N2684) );
  NAND2X0 U7645 ( .IN1(P1_N2625), .IN2(n5316), .QN(n5323) );
  NAND2X0 U7646 ( .IN1(P1_N389), .IN2(P1_N5579), .QN(n5322) );
  NAND2X0 U7647 ( .IN1(n5324), .IN2(n5325), .QN(P1_N2683) );
  NAND2X0 U7648 ( .IN1(P1_N2624), .IN2(n5316), .QN(n5325) );
  NAND2X0 U7649 ( .IN1(P1_N388), .IN2(P1_N5579), .QN(n5324) );
  NAND2X0 U7650 ( .IN1(n5326), .IN2(n5327), .QN(P1_N2682) );
  NAND2X0 U7651 ( .IN1(P1_N2623), .IN2(n5316), .QN(n5327) );
  NAND2X0 U7652 ( .IN1(P1_N387), .IN2(P1_N5579), .QN(n5326) );
  NAND2X0 U7653 ( .IN1(n5328), .IN2(n5329), .QN(P1_N2681) );
  NAND2X0 U7654 ( .IN1(P1_N2622), .IN2(n5316), .QN(n5329) );
  NAND2X0 U7655 ( .IN1(P1_N386), .IN2(P1_N5579), .QN(n5328) );
  NAND2X0 U7656 ( .IN1(n5330), .IN2(n5331), .QN(P1_N2680) );
  NAND2X0 U7657 ( .IN1(P1_N2621), .IN2(n5316), .QN(n5331) );
  NAND2X0 U7658 ( .IN1(P1_N385), .IN2(P1_N5579), .QN(n5330) );
  NAND2X0 U7659 ( .IN1(n5332), .IN2(n5333), .QN(P1_N2679) );
  NAND2X0 U7660 ( .IN1(P1_N2620), .IN2(n5316), .QN(n5333) );
  NAND2X0 U7661 ( .IN1(P1_N384), .IN2(P1_N5579), .QN(n5332) );
  NAND2X0 U7662 ( .IN1(n5334), .IN2(n5335), .QN(P1_N2678) );
  NAND2X0 U7663 ( .IN1(P1_N2619), .IN2(n5316), .QN(n5335) );
  NAND2X0 U7664 ( .IN1(P1_N383), .IN2(P1_N5579), .QN(n5334) );
  NAND2X0 U7665 ( .IN1(n5336), .IN2(n5337), .QN(P1_N2677) );
  NAND2X0 U7666 ( .IN1(P1_N2618), .IN2(n5316), .QN(n5337) );
  NAND2X0 U7667 ( .IN1(P1_N382), .IN2(P1_N5579), .QN(n5336) );
  NAND2X0 U7668 ( .IN1(n5338), .IN2(n5339), .QN(P1_N2676) );
  NAND2X0 U7669 ( .IN1(P1_N2617), .IN2(n5316), .QN(n5339) );
  NAND2X0 U7670 ( .IN1(P1_N381), .IN2(P1_N5579), .QN(n5338) );
  NAND2X0 U7671 ( .IN1(n5340), .IN2(n5341), .QN(P1_N2675) );
  NAND2X0 U7672 ( .IN1(P1_N2616), .IN2(n5316), .QN(n5341) );
  NAND2X0 U7673 ( .IN1(P1_N380), .IN2(P1_N5579), .QN(n5340) );
  NAND2X0 U7674 ( .IN1(n5342), .IN2(n5343), .QN(P1_N2674) );
  NAND2X0 U7675 ( .IN1(P1_N2615), .IN2(n5316), .QN(n5343) );
  NAND2X0 U7676 ( .IN1(P1_N379), .IN2(P1_N5579), .QN(n5342) );
  NAND2X0 U7677 ( .IN1(n5344), .IN2(n5345), .QN(P1_N2673) );
  NAND2X0 U7678 ( .IN1(P1_N2614), .IN2(n5316), .QN(n5345) );
  NAND2X0 U7679 ( .IN1(P1_N378), .IN2(P1_N5579), .QN(n5344) );
  NAND2X0 U7680 ( .IN1(n5346), .IN2(n5347), .QN(P1_N2672) );
  NAND2X0 U7681 ( .IN1(P1_N2613), .IN2(n5316), .QN(n5347) );
  NAND2X0 U7682 ( .IN1(P1_N377), .IN2(P1_N5579), .QN(n5346) );
  NAND2X0 U7683 ( .IN1(n5348), .IN2(n5349), .QN(P1_N2671) );
  NAND2X0 U7684 ( .IN1(P1_N2612), .IN2(n5316), .QN(n5349) );
  NAND2X0 U7685 ( .IN1(P1_N376), .IN2(P1_N5579), .QN(n5348) );
  NAND2X0 U7686 ( .IN1(n5350), .IN2(n5351), .QN(P1_N2670) );
  NAND2X0 U7687 ( .IN1(P1_N2611), .IN2(n5316), .QN(n5351) );
  NAND2X0 U7688 ( .IN1(P1_N375), .IN2(P1_N5579), .QN(n5350) );
  NAND2X0 U7689 ( .IN1(n5352), .IN2(n5353), .QN(P1_N2669) );
  NAND2X0 U7690 ( .IN1(P1_N2610), .IN2(n5316), .QN(n5353) );
  NAND2X0 U7691 ( .IN1(P1_N374), .IN2(P1_N5579), .QN(n5352) );
  NAND2X0 U7692 ( .IN1(n5354), .IN2(n5355), .QN(P1_N2668) );
  NAND2X0 U7693 ( .IN1(P1_N2609), .IN2(n5316), .QN(n5355) );
  NAND2X0 U7694 ( .IN1(P1_N373), .IN2(P1_N5579), .QN(n5354) );
  NAND2X0 U7695 ( .IN1(n5356), .IN2(n5357), .QN(P1_N2667) );
  NAND2X0 U7696 ( .IN1(P1_N2608), .IN2(n5316), .QN(n5357) );
  NAND2X0 U7697 ( .IN1(P1_N372), .IN2(P1_N5579), .QN(n5356) );
  NAND2X0 U7698 ( .IN1(n5358), .IN2(n5359), .QN(P1_N2666) );
  NAND2X0 U7699 ( .IN1(P1_N2607), .IN2(n5316), .QN(n5359) );
  NAND2X0 U7700 ( .IN1(P1_N371), .IN2(P1_N5579), .QN(n5358) );
  NAND2X0 U7701 ( .IN1(n5360), .IN2(n5361), .QN(P1_N2665) );
  NAND2X0 U7702 ( .IN1(P1_N2606), .IN2(n5316), .QN(n5361) );
  NAND2X0 U7703 ( .IN1(P1_N370), .IN2(P1_N5579), .QN(n5360) );
  NAND2X0 U7704 ( .IN1(n5362), .IN2(n5363), .QN(P1_N2664) );
  NAND2X0 U7705 ( .IN1(P1_N2605), .IN2(n5316), .QN(n5363) );
  NAND2X0 U7706 ( .IN1(P1_N369), .IN2(P1_N5579), .QN(n5362) );
  NAND2X0 U7707 ( .IN1(n5364), .IN2(n5365), .QN(P1_N2663) );
  NAND2X0 U7708 ( .IN1(P1_N2604), .IN2(n5316), .QN(n5365) );
  NAND2X0 U7709 ( .IN1(P1_N368), .IN2(P1_N5579), .QN(n5364) );
  NAND2X0 U7710 ( .IN1(n5366), .IN2(n5367), .QN(P1_N2662) );
  NAND2X0 U7711 ( .IN1(P1_N2603), .IN2(n5316), .QN(n5367) );
  NAND2X0 U7712 ( .IN1(n18451), .IN2(P1_N5579), .QN(n5366) );
  NAND2X0 U7713 ( .IN1(n5368), .IN2(n5369), .QN(P1_N2661) );
  NAND2X0 U7714 ( .IN1(P1_N2602), .IN2(n5316), .QN(n5369) );
  NAND2X0 U7715 ( .IN1(n6623), .IN2(P1_N5579), .QN(n5368) );
  NAND2X0 U7716 ( .IN1(n5370), .IN2(n5371), .QN(P1_N2660) );
  NAND2X0 U7717 ( .IN1(P1_N2601), .IN2(n5316), .QN(n5371) );
  NAND2X0 U7524 ( .IN1(P1_N373), .IN2(P1_N5580), .QN(n5250) );
  NAND2X0 U7525 ( .IN1(n5252), .IN2(n5253), .QN(P1_N3040) );
  NAND2X0 U7526 ( .IN1(P1_N2981), .IN2(n5212), .QN(n5253) );
  NAND2X0 U7527 ( .IN1(P1_N372), .IN2(P1_N5580), .QN(n5252) );
  NAND2X0 U7528 ( .IN1(n5254), .IN2(n5255), .QN(P1_N3039) );
  NAND2X0 U7529 ( .IN1(P1_N2980), .IN2(n5212), .QN(n5255) );
  NAND2X0 U7530 ( .IN1(P1_N371), .IN2(P1_N5580), .QN(n5254) );
  NAND2X0 U7531 ( .IN1(n5256), .IN2(n5257), .QN(P1_N3038) );
  NAND2X0 U7532 ( .IN1(P1_N2979), .IN2(n5212), .QN(n5257) );
  NAND2X0 U7533 ( .IN1(P1_N370), .IN2(P1_N5580), .QN(n5256) );
  NAND2X0 U7534 ( .IN1(n5258), .IN2(n5259), .QN(P1_N3037) );
  NAND2X0 U7535 ( .IN1(P1_N2978), .IN2(n5212), .QN(n5259) );
  NAND2X0 U7536 ( .IN1(P1_N369), .IN2(P1_N5580), .QN(n5258) );
  NAND2X0 U7537 ( .IN1(n5260), .IN2(n5261), .QN(P1_N3036) );
  NAND2X0 U7538 ( .IN1(P1_N2977), .IN2(n5212), .QN(n5261) );
  NAND2X0 U7539 ( .IN1(P1_N368), .IN2(P1_N5580), .QN(n5260) );
  NAND2X0 U7540 ( .IN1(n5262), .IN2(n5263), .QN(P1_N3035) );
  NAND2X0 U7541 ( .IN1(P1_N2976), .IN2(n5212), .QN(n5263) );
  NAND2X0 U7542 ( .IN1(n18451), .IN2(P1_N5580), .QN(n5262) );
  NAND2X0 U7543 ( .IN1(n5264), .IN2(n5265), .QN(P1_N3034) );
  NAND2X0 U7544 ( .IN1(P1_N2975), .IN2(n5212), .QN(n5265) );
  NAND2X0 U7545 ( .IN1(n6623), .IN2(P1_N5580), .QN(n5264) );
  NAND2X0 U7546 ( .IN1(n5266), .IN2(n5267), .QN(P1_N3033) );
  NAND2X0 U7547 ( .IN1(P1_N2974), .IN2(n5212), .QN(n5267) );
  NAND2X0 U7548 ( .IN1(n6622), .IN2(P1_N5580), .QN(n5266) );
  NAND2X0 U7549 ( .IN1(n5268), .IN2(n5269), .QN(P1_N3032) );
  NAND2X0 U7550 ( .IN1(P1_N2973), .IN2(n5212), .QN(n5269) );
  NAND2X0 U7553 ( .IN1(n6621), .IN2(P1_N5580), .QN(n5268) );
  AND2X1 U7558 ( .IN1(P1_N248), .IN2(n5272), .Q(P1_N290) );
  NAND2X0 U7559 ( .IN1(n5273), .IN2(n5274), .QN(n5272) );
  NOR2X0 U7560 ( .QN(n5274), .IN1(n5275), .IN2(n5276) );
  NAND2X0 U7561 ( .IN1(n5277), .IN2(n5278), .QN(n5276) );
  NOR2X0 U7562 ( .QN(n5278), .IN1(P1_N264), .IN2(n5279) );
  OR2X1 U7563 ( .IN2(P1_N265), .IN1(P1_N266), .Q(n5279) );
  NOR2X0 U7564 ( .QN(n5277), .IN1(P1_N263), .IN2(P1_N262) );
  NAND2X0 U7565 ( .IN1(n5280), .IN2(n5281), .QN(n5275) );
  NOR2X0 U7566 ( .QN(n5281), .IN1(P1_N269), .IN2(n5282) );
  OR2X1 U7567 ( .IN2(P1_N270), .IN1(P1_N271), .Q(n5282) );
  NOR2X0 U7568 ( .QN(n5280), .IN1(P1_N268), .IN2(P1_N267) );
  NOR2X0 U7569 ( .QN(n5273), .IN1(n5283), .IN2(n5284) );
  NAND2X0 U7570 ( .IN1(n5285), .IN2(n5286), .QN(n5284) );
  NOR2X0 U7571 ( .QN(n5286), .IN1(P1_N256), .IN2(P1_N255) );
  NOR2X0 U7572 ( .QN(n5285), .IN1(P1_N254), .IN2(P1_N253) );
  NAND2X0 U7573 ( .IN1(n5287), .IN2(n5288), .QN(n5283) );
  NOR2X0 U7574 ( .QN(n5288), .IN1(P1_N259), .IN2(n5289) );
  OR2X1 U7575 ( .IN2(P1_N260), .IN1(P1_N261), .Q(n5289) );
  NOR2X0 U7576 ( .QN(n5287), .IN1(P1_N258), .IN2(P1_N257) );
  NAND2X0 U7577 ( .IN1(n7366), .IN2(n5290), .QN(P1_N2880) );
  NAND2X0 U7578 ( .IN1(n7365), .IN2(n5291), .QN(P1_N2878) );
  NOR2X0 U7579 ( .QN(P1_N3061), .IN1(n5291), .IN2(n5290) );
  INVX0 U7580 ( .ZN(n5290), .INP(n7365) );
  INVX0 U7581 ( .ZN(n5291), .INP(n7366) );
  NOR2X0 U7582 ( .QN(P1_N2760), .IN1(n7328), .IN2(n7023) );
  NOR2X0 U7583 ( .QN(P1_N2759), .IN1(n7326), .IN2(n7023) );
  NOR2X0 U7584 ( .QN(P1_N2758), .IN1(n7324), .IN2(n7021) );
  NOR2X0 U7585 ( .QN(P1_N2757), .IN1(n7322), .IN2(n7021) );
  NOR2X0 U7586 ( .QN(P1_N2756), .IN1(n7320), .IN2(n7021) );
  NOR2X0 U7587 ( .QN(P1_N2755), .IN1(n7318), .IN2(n7021) );
  NOR2X0 U7588 ( .QN(P1_N2754), .IN1(n7316), .IN2(n7029) );
  NOR2X0 U7589 ( .QN(P1_N2753), .IN1(n7314), .IN2(n7027) );
  NOR2X0 U7590 ( .QN(P1_N2752), .IN1(n7312), .IN2(n7027) );
  NOR2X0 U7591 ( .QN(P1_N2751), .IN1(n7310), .IN2(n7029) );
  NAND2X0 U7593 ( .IN1(n4097), .IN2(n5293), .QN(P1_N2750) );
  NAND2X0 U7594 ( .IN1(n7019), .IN2(n4099), .QN(n5293) );
  NAND2X0 U7595 ( .IN1(n4100), .IN2(n5294), .QN(P1_N2749) );
  NAND2X0 U7596 ( .IN1(n7019), .IN2(n4102), .QN(n5294) );
  NAND2X0 U7597 ( .IN1(n4103), .IN2(n5295), .QN(P1_N2748) );
  NAND2X0 U7598 ( .IN1(n7028), .IN2(n4105), .QN(n5295) );
  NAND2X0 U7599 ( .IN1(n4106), .IN2(n5296), .QN(P1_N2747) );
  NAND2X0 U7600 ( .IN1(n7028), .IN2(n4108), .QN(n5296) );
  NAND2X0 U7601 ( .IN1(n4109), .IN2(n5297), .QN(P1_N2746) );
  NAND2X0 U7602 ( .IN1(n7028), .IN2(n4111), .QN(n5297) );
  NAND2X0 U7603 ( .IN1(n4112), .IN2(n5298), .QN(P1_N2745) );
  NAND2X0 U7604 ( .IN1(n7024), .IN2(n4114), .QN(n5298) );
  NAND2X0 U7605 ( .IN1(n4115), .IN2(n5299), .QN(P1_N2744) );
  NAND2X0 U7606 ( .IN1(n7024), .IN2(n4117), .QN(n5299) );
  NAND2X0 U7607 ( .IN1(n4118), .IN2(n5300), .QN(P1_N2743) );
  NAND2X0 U7608 ( .IN1(n7024), .IN2(n4120), .QN(n5300) );
  NAND2X0 U7609 ( .IN1(n4121), .IN2(n5301), .QN(P1_N2742) );
  NAND2X0 U7610 ( .IN1(n7024), .IN2(n4123), .QN(n5301) );
  NAND2X0 U7611 ( .IN1(n4124), .IN2(n5302), .QN(P1_N2741) );
  NAND2X0 U7612 ( .IN1(n7024), .IN2(n4126), .QN(n5302) );
  NAND2X0 U7613 ( .IN1(n4127), .IN2(n5303), .QN(P1_N2740) );
  NAND2X0 U7614 ( .IN1(n7463), .IN2(n4129), .QN(n5303) );
  NAND2X0 U7615 ( .IN1(n4130), .IN2(n5304), .QN(P1_N2739) );
  NAND2X0 U7616 ( .IN1(n7463), .IN2(n4132), .QN(n5304) );
  NAND2X0 U7617 ( .IN1(n4133), .IN2(n5305), .QN(P1_N2738) );
  NAND2X0 U7618 ( .IN1(n7463), .IN2(n4135), .QN(n5305) );
  NAND2X0 U7619 ( .IN1(n4136), .IN2(n5306), .QN(P1_N2737) );
  NAND2X0 U7620 ( .IN1(n7463), .IN2(n4138), .QN(n5306) );
  NAND2X0 U7621 ( .IN1(n4139), .IN2(n5307), .QN(P1_N2736) );
  NAND2X0 U7622 ( .IN1(n7026), .IN2(n4141), .QN(n5307) );
  NAND2X0 U7429 ( .IN1(n4106), .IN2(n5192), .QN(P1_N3120) );
  NAND2X0 U7430 ( .IN1(n7028), .IN2(n4108), .QN(n5192) );
  NAND2X0 U7431 ( .IN1(n4109), .IN2(n5193), .QN(P1_N3119) );
  NAND2X0 U7432 ( .IN1(n7028), .IN2(n4111), .QN(n5193) );
  NAND2X0 U7433 ( .IN1(n4112), .IN2(n5194), .QN(P1_N3118) );
  NAND2X0 U7434 ( .IN1(n7024), .IN2(n4114), .QN(n5194) );
  NAND2X0 U7435 ( .IN1(n4115), .IN2(n5195), .QN(P1_N3117) );
  NAND2X0 U7436 ( .IN1(n7024), .IN2(n4117), .QN(n5195) );
  NAND2X0 U7437 ( .IN1(n4118), .IN2(n5196), .QN(P1_N3116) );
  NAND2X0 U7438 ( .IN1(n7024), .IN2(n4120), .QN(n5196) );
  NAND2X0 U7439 ( .IN1(n4121), .IN2(n5197), .QN(P1_N3115) );
  NAND2X0 U7440 ( .IN1(n7024), .IN2(n4123), .QN(n5197) );
  NAND2X0 U7441 ( .IN1(n4124), .IN2(n5198), .QN(P1_N3114) );
  NAND2X0 U7442 ( .IN1(n7024), .IN2(n4126), .QN(n5198) );
  NAND2X0 U7443 ( .IN1(n4127), .IN2(n5199), .QN(P1_N3113) );
  NAND2X0 U7444 ( .IN1(n7463), .IN2(n4129), .QN(n5199) );
  NAND2X0 U7445 ( .IN1(n4130), .IN2(n5200), .QN(P1_N3112) );
  NAND2X0 U7446 ( .IN1(n7463), .IN2(n4132), .QN(n5200) );
  NAND2X0 U7447 ( .IN1(n4133), .IN2(n5201), .QN(P1_N3111) );
  NAND2X0 U7448 ( .IN1(n7463), .IN2(n4135), .QN(n5201) );
  NAND2X0 U7449 ( .IN1(n4136), .IN2(n5202), .QN(P1_N3110) );
  NAND2X0 U7450 ( .IN1(n7463), .IN2(n4138), .QN(n5202) );
  NAND2X0 U7451 ( .IN1(n4139), .IN2(n5203), .QN(P1_N3109) );
  NAND2X0 U7452 ( .IN1(n7026), .IN2(n4141), .QN(n5203) );
  NAND2X0 U7453 ( .IN1(n4142), .IN2(n5204), .QN(P1_N3108) );
  NAND2X0 U7454 ( .IN1(n7026), .IN2(n4144), .QN(n5204) );
  NAND2X0 U7455 ( .IN1(n4145), .IN2(n5205), .QN(P1_N3107) );
  NAND2X0 U7456 ( .IN1(n7026), .IN2(n4147), .QN(n5205) );
  NAND2X0 U7457 ( .IN1(n4148), .IN2(n5206), .QN(P1_N3106) );
  NAND2X0 U7458 ( .IN1(n7022), .IN2(n4150), .QN(n5206) );
  NAND2X0 U7459 ( .IN1(n4151), .IN2(n5207), .QN(P1_N3105) );
  NAND2X0 U7460 ( .IN1(n7022), .IN2(n4153), .QN(n5207) );
  NAND2X0 U7461 ( .IN1(n4154), .IN2(n5208), .QN(P1_N3104) );
  NAND2X0 U7462 ( .IN1(n7022), .IN2(n4156), .QN(n5208) );
  NAND2X0 U7465 ( .IN1(n5210), .IN2(n5211), .QN(P1_N3060) );
  NAND2X0 U7466 ( .IN1(P1_N3001), .IN2(n5212), .QN(n5211) );
  NAND2X0 U7467 ( .IN1(P1_N392), .IN2(P1_N5580), .QN(n5210) );
  NAND2X0 U7468 ( .IN1(n5214), .IN2(n5215), .QN(P1_N3059) );
  NAND2X0 U7469 ( .IN1(P1_N3000), .IN2(n5212), .QN(n5215) );
  NAND2X0 U7470 ( .IN1(P1_N391), .IN2(P1_N5580), .QN(n5214) );
  NAND2X0 U7471 ( .IN1(n5216), .IN2(n5217), .QN(P1_N3058) );
  NAND2X0 U7472 ( .IN1(P1_N2999), .IN2(n5212), .QN(n5217) );
  NAND2X0 U7473 ( .IN1(P1_N390), .IN2(P1_N5580), .QN(n5216) );
  NAND2X0 U7474 ( .IN1(n5218), .IN2(n5219), .QN(P1_N3057) );
  NAND2X0 U7475 ( .IN1(P1_N2998), .IN2(n5212), .QN(n5219) );
  NAND2X0 U7476 ( .IN1(P1_N389), .IN2(P1_N5580), .QN(n5218) );
  NAND2X0 U7477 ( .IN1(n5220), .IN2(n5221), .QN(P1_N3056) );
  NAND2X0 U7478 ( .IN1(P1_N2997), .IN2(n5212), .QN(n5221) );
  NAND2X0 U7479 ( .IN1(P1_N388), .IN2(P1_N5580), .QN(n5220) );
  NAND2X0 U7480 ( .IN1(n5222), .IN2(n5223), .QN(P1_N3055) );
  NAND2X0 U7481 ( .IN1(P1_N2996), .IN2(n5212), .QN(n5223) );
  NAND2X0 U7482 ( .IN1(P1_N387), .IN2(P1_N5580), .QN(n5222) );
  NAND2X0 U7483 ( .IN1(n5224), .IN2(n5225), .QN(P1_N3054) );
  NAND2X0 U7484 ( .IN1(P1_N2995), .IN2(n5212), .QN(n5225) );
  NAND2X0 U7485 ( .IN1(P1_N386), .IN2(P1_N5580), .QN(n5224) );
  NAND2X0 U7486 ( .IN1(n5226), .IN2(n5227), .QN(P1_N3053) );
  NAND2X0 U7487 ( .IN1(P1_N2994), .IN2(n5212), .QN(n5227) );
  NAND2X0 U7488 ( .IN1(P1_N385), .IN2(P1_N5580), .QN(n5226) );
  NAND2X0 U7489 ( .IN1(n5228), .IN2(n5229), .QN(P1_N3052) );
  NAND2X0 U7490 ( .IN1(P1_N2993), .IN2(n5212), .QN(n5229) );
  NAND2X0 U7491 ( .IN1(P1_N384), .IN2(P1_N5580), .QN(n5228) );
  NAND2X0 U7492 ( .IN1(n5230), .IN2(n5231), .QN(P1_N3051) );
  NAND2X0 U7493 ( .IN1(P1_N2992), .IN2(n5212), .QN(n5231) );
  NAND2X0 U7494 ( .IN1(P1_N383), .IN2(P1_N5580), .QN(n5230) );
  NAND2X0 U7495 ( .IN1(n5232), .IN2(n5233), .QN(P1_N3050) );
  NAND2X0 U7496 ( .IN1(P1_N2991), .IN2(n5212), .QN(n5233) );
  NAND2X0 U7497 ( .IN1(P1_N382), .IN2(P1_N5580), .QN(n5232) );
  NAND2X0 U7498 ( .IN1(n5234), .IN2(n5235), .QN(P1_N3049) );
  NAND2X0 U7499 ( .IN1(P1_N2990), .IN2(n5212), .QN(n5235) );
  NAND2X0 U7500 ( .IN1(P1_N381), .IN2(P1_N5580), .QN(n5234) );
  NAND2X0 U7501 ( .IN1(n5236), .IN2(n5237), .QN(P1_N3048) );
  NAND2X0 U7502 ( .IN1(P1_N2989), .IN2(n5212), .QN(n5237) );
  NAND2X0 U7503 ( .IN1(P1_N380), .IN2(P1_N5580), .QN(n5236) );
  NAND2X0 U7504 ( .IN1(n5238), .IN2(n5239), .QN(P1_N3047) );
  NAND2X0 U7505 ( .IN1(P1_N2988), .IN2(n5212), .QN(n5239) );
  NAND2X0 U7506 ( .IN1(P1_N379), .IN2(P1_N5580), .QN(n5238) );
  NAND2X0 U7507 ( .IN1(n5240), .IN2(n5241), .QN(P1_N3046) );
  NAND2X0 U7508 ( .IN1(P1_N2987), .IN2(n5212), .QN(n5241) );
  NAND2X0 U7509 ( .IN1(P1_N378), .IN2(P1_N5580), .QN(n5240) );
  NAND2X0 U7510 ( .IN1(n5242), .IN2(n5243), .QN(P1_N3045) );
  NAND2X0 U7511 ( .IN1(P1_N2986), .IN2(n5212), .QN(n5243) );
  NAND2X0 U7512 ( .IN1(P1_N377), .IN2(P1_N5580), .QN(n5242) );
  NAND2X0 U7513 ( .IN1(n5244), .IN2(n5245), .QN(P1_N3044) );
  NAND2X0 U7514 ( .IN1(P1_N2985), .IN2(n5212), .QN(n5245) );
  NAND2X0 U7515 ( .IN1(P1_N376), .IN2(P1_N5580), .QN(n5244) );
  NAND2X0 U7516 ( .IN1(n5246), .IN2(n5247), .QN(P1_N3043) );
  NAND2X0 U7517 ( .IN1(P1_N2984), .IN2(n5212), .QN(n5247) );
  NAND2X0 U7518 ( .IN1(P1_N375), .IN2(P1_N5580), .QN(n5246) );
  NAND2X0 U7519 ( .IN1(n5248), .IN2(n5249), .QN(P1_N3042) );
  NAND2X0 U7520 ( .IN1(P1_N2983), .IN2(n5212), .QN(n5249) );
  NAND2X0 U7521 ( .IN1(P1_N374), .IN2(P1_N5580), .QN(n5248) );
  NAND2X0 U7522 ( .IN1(n5250), .IN2(n5251), .QN(P1_N3041) );
  NAND2X0 U7523 ( .IN1(P1_N2982), .IN2(n5212), .QN(n5251) );
  NAND2X0 U7330 ( .IN1(n5130), .IN2(n5131), .QN(P1_N3420) );
  NAND2X0 U7331 ( .IN1(P1_N3361), .IN2(n5104), .QN(n5131) );
  NAND2X0 U7332 ( .IN1(P1_N379), .IN2(P1_N5581), .QN(n5130) );
  AND2X1 U7333 ( .IN1(P1_N295), .IN2(n5132), .Q(P1_N342) );
  NAND2X0 U7334 ( .IN1(n5133), .IN2(n5134), .QN(n5132) );
  NOR2X0 U7335 ( .QN(n5134), .IN1(n5135), .IN2(n5136) );
  NAND2X0 U7336 ( .IN1(n5137), .IN2(n5138), .QN(n5136) );
  NOR2X0 U7337 ( .QN(n5138), .IN1(P1_N311), .IN2(n5139) );
  OR2X1 U7338 ( .IN2(P1_N312), .IN1(P1_N313), .Q(n5139) );
  NOR2X0 U7339 ( .QN(n5137), .IN1(P1_N308), .IN2(n5140) );
  OR2X1 U7340 ( .IN2(P1_N309), .IN1(P1_N310), .Q(n5140) );
  NAND2X0 U7341 ( .IN1(n5141), .IN2(n5142), .QN(n5135) );
  NOR2X0 U7342 ( .QN(n5142), .IN1(P1_N317), .IN2(n5143) );
  OR2X1 U7343 ( .IN2(P1_N318), .IN1(P1_N319), .Q(n5143) );
  NOR2X0 U7344 ( .QN(n5141), .IN1(P1_N314), .IN2(n5144) );
  OR2X1 U7345 ( .IN2(P1_N315), .IN1(P1_N316), .Q(n5144) );
  NOR2X0 U7346 ( .QN(n5133), .IN1(n5145), .IN2(n5146) );
  NAND2X0 U7347 ( .IN1(n5147), .IN2(n5148), .QN(n5146) );
  NOR2X0 U7348 ( .QN(n5148), .IN1(P1_N299), .IN2(n5149) );
  OR2X1 U7349 ( .IN2(P1_N300), .IN1(P1_N301), .Q(n5149) );
  NOR2X0 U7350 ( .QN(n5147), .IN1(P1_N298), .IN2(P1_N297) );
  NAND2X0 U7351 ( .IN1(n5150), .IN2(n5151), .QN(n5145) );
  NOR2X0 U7352 ( .QN(n5151), .IN1(P1_N305), .IN2(n5152) );
  OR2X1 U7353 ( .IN2(P1_N306), .IN1(P1_N307), .Q(n5152) );
  NOR2X0 U7354 ( .QN(n5150), .IN1(P1_N302), .IN2(n5153) );
  OR2X1 U7355 ( .IN2(P1_N303), .IN1(P1_N304), .Q(n5153) );
  NAND2X0 U7356 ( .IN1(n5154), .IN2(n5155), .QN(P1_N3419) );
  NAND2X0 U7357 ( .IN1(P1_N3360), .IN2(n5104), .QN(n5155) );
  NAND2X0 U7358 ( .IN1(P1_N378), .IN2(P1_N5581), .QN(n5154) );
  NAND2X0 U7359 ( .IN1(n5156), .IN2(n5157), .QN(P1_N3418) );
  NAND2X0 U7360 ( .IN1(P1_N3359), .IN2(n5104), .QN(n5157) );
  NAND2X0 U7361 ( .IN1(P1_N377), .IN2(P1_N5581), .QN(n5156) );
  NAND2X0 U7362 ( .IN1(n5158), .IN2(n5159), .QN(P1_N3417) );
  NAND2X0 U7363 ( .IN1(P1_N3358), .IN2(n5104), .QN(n5159) );
  NAND2X0 U7364 ( .IN1(P1_N376), .IN2(P1_N5581), .QN(n5158) );
  NAND2X0 U7365 ( .IN1(n5160), .IN2(n5161), .QN(P1_N3416) );
  NAND2X0 U7366 ( .IN1(P1_N3357), .IN2(n5104), .QN(n5161) );
  NAND2X0 U7367 ( .IN1(P1_N375), .IN2(P1_N5581), .QN(n5160) );
  NAND2X0 U7368 ( .IN1(n5162), .IN2(n5163), .QN(P1_N3415) );
  NAND2X0 U7369 ( .IN1(P1_N3356), .IN2(n5104), .QN(n5163) );
  NAND2X0 U7370 ( .IN1(P1_N374), .IN2(P1_N5581), .QN(n5162) );
  NAND2X0 U7371 ( .IN1(n5164), .IN2(n5165), .QN(P1_N3414) );
  NAND2X0 U7372 ( .IN1(P1_N3355), .IN2(n5104), .QN(n5165) );
  NAND2X0 U7373 ( .IN1(P1_N373), .IN2(P1_N5581), .QN(n5164) );
  NAND2X0 U7374 ( .IN1(n5166), .IN2(n5167), .QN(P1_N3413) );
  NAND2X0 U7375 ( .IN1(P1_N3354), .IN2(n5104), .QN(n5167) );
  NAND2X0 U7376 ( .IN1(P1_N372), .IN2(P1_N5581), .QN(n5166) );
  NAND2X0 U7377 ( .IN1(n5168), .IN2(n5169), .QN(P1_N3412) );
  NAND2X0 U7378 ( .IN1(P1_N3353), .IN2(n5104), .QN(n5169) );
  NAND2X0 U7379 ( .IN1(P1_N371), .IN2(P1_N5581), .QN(n5168) );
  NAND2X0 U7380 ( .IN1(n5170), .IN2(n5171), .QN(P1_N3411) );
  NAND2X0 U7381 ( .IN1(P1_N3352), .IN2(n5104), .QN(n5171) );
  NAND2X0 U7382 ( .IN1(P1_N370), .IN2(P1_N5581), .QN(n5170) );
  NAND2X0 U7383 ( .IN1(n5172), .IN2(n5173), .QN(P1_N3410) );
  NAND2X0 U7384 ( .IN1(P1_N3351), .IN2(n5104), .QN(n5173) );
  NAND2X0 U7385 ( .IN1(P1_N369), .IN2(P1_N5581), .QN(n5172) );
  NAND2X0 U7386 ( .IN1(n5174), .IN2(n5175), .QN(P1_N3409) );
  NAND2X0 U7387 ( .IN1(P1_N3350), .IN2(n5104), .QN(n5175) );
  NAND2X0 U7388 ( .IN1(P1_N368), .IN2(P1_N5581), .QN(n5174) );
  NAND2X0 U7389 ( .IN1(n5176), .IN2(n5177), .QN(P1_N3408) );
  NAND2X0 U7390 ( .IN1(P1_N3349), .IN2(n5104), .QN(n5177) );
  NAND2X0 U7391 ( .IN1(n18451), .IN2(P1_N5581), .QN(n5176) );
  NAND2X0 U7392 ( .IN1(n5178), .IN2(n5179), .QN(P1_N3407) );
  NAND2X0 U7393 ( .IN1(P1_N3348), .IN2(n5104), .QN(n5179) );
  NAND2X0 U7394 ( .IN1(n6623), .IN2(P1_N5581), .QN(n5178) );
  NAND2X0 U7395 ( .IN1(n5180), .IN2(n5181), .QN(P1_N3406) );
  NAND2X0 U7396 ( .IN1(P1_N3347), .IN2(n5104), .QN(n5181) );
  NAND2X0 U7397 ( .IN1(n6622), .IN2(P1_N5581), .QN(n5180) );
  NAND2X0 U7398 ( .IN1(n5182), .IN2(n5183), .QN(P1_N3405) );
  NAND2X0 U7399 ( .IN1(P1_N3346), .IN2(n5104), .QN(n5183) );
  NAND2X0 U7402 ( .IN1(n6621), .IN2(P1_N5581), .QN(n5182) );
  NAND2X0 U7407 ( .IN1(n7368), .IN2(n5186), .QN(P1_N3253) );
  NAND2X0 U7408 ( .IN1(n7367), .IN2(n5187), .QN(P1_N3251) );
  NOR2X0 U7409 ( .QN(P1_N3434), .IN1(n5187), .IN2(n5186) );
  INVX0 U7410 ( .ZN(n5186), .INP(n7367) );
  INVX0 U7411 ( .ZN(n5187), .INP(n7368) );
  NOR2X0 U7412 ( .QN(P1_N3133), .IN1(n7328), .IN2(n7023) );
  NOR2X0 U7413 ( .QN(P1_N3132), .IN1(n7326), .IN2(n7023) );
  NOR2X0 U7414 ( .QN(P1_N3131), .IN1(n7324), .IN2(n7021) );
  NOR2X0 U7415 ( .QN(P1_N3130), .IN1(n7322), .IN2(n7021) );
  NOR2X0 U7416 ( .QN(P1_N3129), .IN1(n7320), .IN2(n7021) );
  NOR2X0 U7417 ( .QN(P1_N3128), .IN1(n7318), .IN2(n7021) );
  NOR2X0 U7418 ( .QN(P1_N3127), .IN1(n7316), .IN2(n7027) );
  NOR2X0 U7419 ( .QN(P1_N3126), .IN1(n7314), .IN2(n7027) );
  NOR2X0 U7420 ( .QN(P1_N3125), .IN1(n7312), .IN2(n7027) );
  NOR2X0 U7421 ( .QN(P1_N3124), .IN1(n7310), .IN2(n7027) );
  NAND2X0 U7423 ( .IN1(n4097), .IN2(n5189), .QN(P1_N3123) );
  NAND2X0 U7424 ( .IN1(n7019), .IN2(n4099), .QN(n5189) );
  NAND2X0 U7425 ( .IN1(n4100), .IN2(n5190), .QN(P1_N3122) );
  NAND2X0 U7426 ( .IN1(n7028), .IN2(n4102), .QN(n5190) );
  NAND2X0 U7427 ( .IN1(n4103), .IN2(n5191), .QN(P1_N3121) );
  NAND2X0 U7428 ( .IN1(n7028), .IN2(n4105), .QN(n5191) );
  NAND2X0 U7234 ( .IN1(n7369), .IN2(n5079), .QN(P1_N3624) );
  NOR2X0 U7235 ( .QN(P1_N3807), .IN1(n5079), .IN2(n5078) );
  INVX0 U7236 ( .ZN(n5078), .INP(n7369) );
  INVX0 U7237 ( .ZN(n5079), .INP(n7370) );
  NOR2X0 U7238 ( .QN(P1_N3506), .IN1(n7328), .IN2(n7023) );
  NOR2X0 U7239 ( .QN(P1_N3505), .IN1(n7326), .IN2(n7023) );
  NOR2X0 U7240 ( .QN(P1_N3504), .IN1(n7324), .IN2(n7021) );
  NOR2X0 U7241 ( .QN(P1_N3503), .IN1(n7322), .IN2(n7021) );
  NOR2X0 U7242 ( .QN(P1_N3502), .IN1(n7320), .IN2(n7021) );
  NOR2X0 U7243 ( .QN(P1_N3501), .IN1(n7318), .IN2(n7021) );
  NOR2X0 U7244 ( .QN(P1_N3500), .IN1(n7316), .IN2(n7029) );
  NOR2X0 U7245 ( .QN(P1_N3499), .IN1(n7314), .IN2(n7027) );
  NOR2X0 U7246 ( .QN(P1_N3498), .IN1(n7312), .IN2(n7027) );
  NOR2X0 U7247 ( .QN(P1_N3497), .IN1(n7310), .IN2(n7029) );
  NAND2X0 U7249 ( .IN1(n4097), .IN2(n5081), .QN(P1_N3496) );
  NAND2X0 U7250 ( .IN1(n7019), .IN2(n4099), .QN(n5081) );
  NAND2X0 U7251 ( .IN1(n4100), .IN2(n5082), .QN(P1_N3495) );
  NAND2X0 U7252 ( .IN1(n7028), .IN2(n4102), .QN(n5082) );
  NAND2X0 U7253 ( .IN1(n4103), .IN2(n5083), .QN(P1_N3494) );
  NAND2X0 U7254 ( .IN1(n7028), .IN2(n4105), .QN(n5083) );
  NAND2X0 U7255 ( .IN1(n4106), .IN2(n5084), .QN(P1_N3493) );
  NAND2X0 U7256 ( .IN1(n7028), .IN2(n4108), .QN(n5084) );
  NAND2X0 U7257 ( .IN1(n4109), .IN2(n5085), .QN(P1_N3492) );
  NAND2X0 U7258 ( .IN1(n7028), .IN2(n4111), .QN(n5085) );
  NAND2X0 U7259 ( .IN1(n4112), .IN2(n5086), .QN(P1_N3491) );
  NAND2X0 U7260 ( .IN1(n7024), .IN2(n4114), .QN(n5086) );
  NAND2X0 U7261 ( .IN1(n4115), .IN2(n5087), .QN(P1_N3490) );
  NAND2X0 U7262 ( .IN1(n7024), .IN2(n4117), .QN(n5087) );
  NAND2X0 U7263 ( .IN1(n4118), .IN2(n5088), .QN(P1_N3489) );
  NAND2X0 U7264 ( .IN1(n7024), .IN2(n4120), .QN(n5088) );
  NAND2X0 U7265 ( .IN1(n4121), .IN2(n5089), .QN(P1_N3488) );
  NAND2X0 U7266 ( .IN1(n7024), .IN2(n4123), .QN(n5089) );
  NAND2X0 U7267 ( .IN1(n4124), .IN2(n5090), .QN(P1_N3487) );
  NAND2X0 U7268 ( .IN1(n7024), .IN2(n4126), .QN(n5090) );
  NAND2X0 U7269 ( .IN1(n4127), .IN2(n5091), .QN(P1_N3486) );
  NAND2X0 U7270 ( .IN1(n7463), .IN2(n4129), .QN(n5091) );
  NAND2X0 U7271 ( .IN1(n4130), .IN2(n5092), .QN(P1_N3485) );
  NAND2X0 U7272 ( .IN1(n7463), .IN2(n4132), .QN(n5092) );
  NAND2X0 U7273 ( .IN1(n4133), .IN2(n5093), .QN(P1_N3484) );
  NAND2X0 U7274 ( .IN1(n7463), .IN2(n4135), .QN(n5093) );
  NAND2X0 U7275 ( .IN1(n4136), .IN2(n5094), .QN(P1_N3483) );
  NAND2X0 U7276 ( .IN1(n7463), .IN2(n4138), .QN(n5094) );
  NAND2X0 U7277 ( .IN1(n4139), .IN2(n5095), .QN(P1_N3482) );
  NAND2X0 U7278 ( .IN1(n7026), .IN2(n4141), .QN(n5095) );
  NAND2X0 U7279 ( .IN1(n4142), .IN2(n5096), .QN(P1_N3481) );
  NAND2X0 U7280 ( .IN1(n7026), .IN2(n4144), .QN(n5096) );
  NAND2X0 U7281 ( .IN1(n4145), .IN2(n5097), .QN(P1_N3480) );
  NAND2X0 U7282 ( .IN1(n7026), .IN2(n4147), .QN(n5097) );
  NAND2X0 U7283 ( .IN1(n4148), .IN2(n5098), .QN(P1_N3479) );
  NAND2X0 U7284 ( .IN1(n7022), .IN2(n4150), .QN(n5098) );
  NAND2X0 U7285 ( .IN1(n4151), .IN2(n5099), .QN(P1_N3478) );
  NAND2X0 U7286 ( .IN1(n7022), .IN2(n4153), .QN(n5099) );
  NAND2X0 U7287 ( .IN1(n4154), .IN2(n5100), .QN(P1_N3477) );
  NAND2X0 U7288 ( .IN1(n7022), .IN2(n4156), .QN(n5100) );
  NAND2X0 U7291 ( .IN1(n5102), .IN2(n5103), .QN(P1_N3433) );
  NAND2X0 U7292 ( .IN1(P1_N3374), .IN2(n5104), .QN(n5103) );
  NAND2X0 U7293 ( .IN1(P1_N392), .IN2(P1_N5581), .QN(n5102) );
  NAND2X0 U7294 ( .IN1(n5106), .IN2(n5107), .QN(P1_N3432) );
  NAND2X0 U7295 ( .IN1(P1_N3373), .IN2(n5104), .QN(n5107) );
  NAND2X0 U7296 ( .IN1(P1_N391), .IN2(P1_N5581), .QN(n5106) );
  NAND2X0 U7297 ( .IN1(n5108), .IN2(n5109), .QN(P1_N3431) );
  NAND2X0 U7298 ( .IN1(P1_N3372), .IN2(n5104), .QN(n5109) );
  NAND2X0 U7299 ( .IN1(P1_N390), .IN2(P1_N5581), .QN(n5108) );
  NAND2X0 U7300 ( .IN1(n5110), .IN2(n5111), .QN(P1_N3430) );
  NAND2X0 U7301 ( .IN1(P1_N3371), .IN2(n5104), .QN(n5111) );
  NAND2X0 U7302 ( .IN1(P1_N389), .IN2(P1_N5581), .QN(n5110) );
  NAND2X0 U7303 ( .IN1(n5112), .IN2(n5113), .QN(P1_N3429) );
  NAND2X0 U7304 ( .IN1(P1_N3370), .IN2(n5104), .QN(n5113) );
  NAND2X0 U7305 ( .IN1(P1_N388), .IN2(P1_N5581), .QN(n5112) );
  NAND2X0 U7306 ( .IN1(n5114), .IN2(n5115), .QN(P1_N3428) );
  NAND2X0 U7307 ( .IN1(P1_N3369), .IN2(n5104), .QN(n5115) );
  NAND2X0 U7308 ( .IN1(P1_N387), .IN2(P1_N5581), .QN(n5114) );
  NAND2X0 U7309 ( .IN1(n5116), .IN2(n5117), .QN(P1_N3427) );
  NAND2X0 U7310 ( .IN1(P1_N3368), .IN2(n5104), .QN(n5117) );
  NAND2X0 U7311 ( .IN1(P1_N386), .IN2(P1_N5581), .QN(n5116) );
  NAND2X0 U7312 ( .IN1(n5118), .IN2(n5119), .QN(P1_N3426) );
  NAND2X0 U7313 ( .IN1(P1_N3367), .IN2(n5104), .QN(n5119) );
  NAND2X0 U7314 ( .IN1(P1_N385), .IN2(P1_N5581), .QN(n5118) );
  NAND2X0 U7315 ( .IN1(n5120), .IN2(n5121), .QN(P1_N3425) );
  NAND2X0 U7316 ( .IN1(P1_N3366), .IN2(n5104), .QN(n5121) );
  NAND2X0 U7317 ( .IN1(P1_N384), .IN2(P1_N5581), .QN(n5120) );
  NAND2X0 U7318 ( .IN1(n5122), .IN2(n5123), .QN(P1_N3424) );
  NAND2X0 U7319 ( .IN1(P1_N3365), .IN2(n5104), .QN(n5123) );
  NAND2X0 U7320 ( .IN1(P1_N383), .IN2(P1_N5581), .QN(n5122) );
  NAND2X0 U7321 ( .IN1(n5124), .IN2(n5125), .QN(P1_N3423) );
  NAND2X0 U7322 ( .IN1(P1_N3364), .IN2(n5104), .QN(n5125) );
  NAND2X0 U7323 ( .IN1(P1_N382), .IN2(P1_N5581), .QN(n5124) );
  NAND2X0 U7324 ( .IN1(n5126), .IN2(n5127), .QN(P1_N3422) );
  NAND2X0 U7325 ( .IN1(P1_N3363), .IN2(n5104), .QN(n5127) );
  NAND2X0 U7326 ( .IN1(P1_N381), .IN2(P1_N5581), .QN(n5126) );
  NAND2X0 U7327 ( .IN1(n5128), .IN2(n5129), .QN(P1_N3421) );
  NAND2X0 U7328 ( .IN1(P1_N3362), .IN2(n5104), .QN(n5129) );
  NAND2X0 U7329 ( .IN1(P1_N380), .IN2(P1_N5581), .QN(n5128) );
  NAND2X0 U7134 ( .IN1(n4151), .IN2(n5013), .QN(P1_N3851) );
  NAND2X0 U7135 ( .IN1(n7022), .IN2(n4153), .QN(n5013) );
  NAND2X0 U7136 ( .IN1(n4154), .IN2(n5014), .QN(P1_N3850) );
  NAND2X0 U7137 ( .IN1(n7022), .IN2(n4156), .QN(n5014) );
  NAND2X0 U7140 ( .IN1(n5016), .IN2(n5017), .QN(P1_N3806) );
  NAND2X0 U7141 ( .IN1(P1_N3747), .IN2(n5018), .QN(n5017) );
  NAND2X0 U7142 ( .IN1(P1_N392), .IN2(P1_N5582), .QN(n5016) );
  NAND2X0 U7143 ( .IN1(n5020), .IN2(n5021), .QN(P1_N3805) );
  NAND2X0 U7144 ( .IN1(P1_N3746), .IN2(n5018), .QN(n5021) );
  NAND2X0 U7145 ( .IN1(P1_N391), .IN2(P1_N5582), .QN(n5020) );
  NAND2X0 U7146 ( .IN1(n5022), .IN2(n5023), .QN(P1_N3804) );
  NAND2X0 U7147 ( .IN1(P1_N3745), .IN2(n5018), .QN(n5023) );
  NAND2X0 U7148 ( .IN1(P1_N390), .IN2(P1_N5582), .QN(n5022) );
  NAND2X0 U7149 ( .IN1(n5024), .IN2(n5025), .QN(P1_N3803) );
  NAND2X0 U7150 ( .IN1(P1_N3744), .IN2(n5018), .QN(n5025) );
  NAND2X0 U7151 ( .IN1(P1_N389), .IN2(P1_N5582), .QN(n5024) );
  NAND2X0 U7152 ( .IN1(n5026), .IN2(n5027), .QN(P1_N3802) );
  NAND2X0 U7153 ( .IN1(P1_N3743), .IN2(n5018), .QN(n5027) );
  NAND2X0 U7154 ( .IN1(P1_N388), .IN2(P1_N5582), .QN(n5026) );
  NAND2X0 U7155 ( .IN1(n5028), .IN2(n5029), .QN(P1_N3801) );
  NAND2X0 U7156 ( .IN1(P1_N3742), .IN2(n5018), .QN(n5029) );
  NAND2X0 U7157 ( .IN1(P1_N387), .IN2(P1_N5582), .QN(n5028) );
  NAND2X0 U7158 ( .IN1(n5030), .IN2(n5031), .QN(P1_N3800) );
  NAND2X0 U7159 ( .IN1(P1_N3741), .IN2(n5018), .QN(n5031) );
  NAND2X0 U7160 ( .IN1(P1_N386), .IN2(P1_N5582), .QN(n5030) );
  NAND2X0 U7161 ( .IN1(n5032), .IN2(n5033), .QN(P1_N3799) );
  NAND2X0 U7162 ( .IN1(P1_N3740), .IN2(n5018), .QN(n5033) );
  NAND2X0 U7163 ( .IN1(P1_N385), .IN2(P1_N5582), .QN(n5032) );
  NAND2X0 U7164 ( .IN1(n5034), .IN2(n5035), .QN(P1_N3798) );
  NAND2X0 U7165 ( .IN1(P1_N3739), .IN2(n5018), .QN(n5035) );
  NAND2X0 U7166 ( .IN1(P1_N384), .IN2(P1_N5582), .QN(n5034) );
  NAND2X0 U7167 ( .IN1(n5036), .IN2(n5037), .QN(P1_N3797) );
  NAND2X0 U7168 ( .IN1(P1_N3738), .IN2(n5018), .QN(n5037) );
  NAND2X0 U7169 ( .IN1(P1_N383), .IN2(P1_N5582), .QN(n5036) );
  NAND2X0 U7170 ( .IN1(n5038), .IN2(n5039), .QN(P1_N3796) );
  NAND2X0 U7171 ( .IN1(P1_N3737), .IN2(n5018), .QN(n5039) );
  NAND2X0 U7172 ( .IN1(P1_N382), .IN2(P1_N5582), .QN(n5038) );
  NAND2X0 U7173 ( .IN1(n5040), .IN2(n5041), .QN(P1_N3795) );
  NAND2X0 U7174 ( .IN1(P1_N3736), .IN2(n5018), .QN(n5041) );
  NAND2X0 U7175 ( .IN1(P1_N381), .IN2(P1_N5582), .QN(n5040) );
  NAND2X0 U7176 ( .IN1(n5042), .IN2(n5043), .QN(P1_N3794) );
  NAND2X0 U7177 ( .IN1(P1_N3735), .IN2(n5018), .QN(n5043) );
  NAND2X0 U7178 ( .IN1(P1_N380), .IN2(P1_N5582), .QN(n5042) );
  NAND2X0 U7179 ( .IN1(n5044), .IN2(n5045), .QN(P1_N3793) );
  NAND2X0 U7180 ( .IN1(P1_N3734), .IN2(n5018), .QN(n5045) );
  NAND2X0 U7181 ( .IN1(P1_N379), .IN2(P1_N5582), .QN(n5044) );
  NAND2X0 U7182 ( .IN1(n5046), .IN2(n5047), .QN(P1_N3792) );
  NAND2X0 U7183 ( .IN1(P1_N3733), .IN2(n5018), .QN(n5047) );
  NAND2X0 U7184 ( .IN1(P1_N378), .IN2(P1_N5582), .QN(n5046) );
  NAND2X0 U7185 ( .IN1(n5048), .IN2(n5049), .QN(P1_N3791) );
  NAND2X0 U7186 ( .IN1(P1_N3732), .IN2(n5018), .QN(n5049) );
  NAND2X0 U7187 ( .IN1(P1_N377), .IN2(P1_N5582), .QN(n5048) );
  NAND2X0 U7188 ( .IN1(n5050), .IN2(n5051), .QN(P1_N3790) );
  NAND2X0 U7189 ( .IN1(P1_N3731), .IN2(n5018), .QN(n5051) );
  NAND2X0 U7190 ( .IN1(P1_N376), .IN2(P1_N5582), .QN(n5050) );
  NAND2X0 U7191 ( .IN1(n5052), .IN2(n5053), .QN(P1_N3789) );
  NAND2X0 U7192 ( .IN1(P1_N3730), .IN2(n5018), .QN(n5053) );
  NAND2X0 U7193 ( .IN1(P1_N375), .IN2(P1_N5582), .QN(n5052) );
  NAND2X0 U7194 ( .IN1(n5054), .IN2(n5055), .QN(P1_N3788) );
  NAND2X0 U7195 ( .IN1(P1_N3729), .IN2(n5018), .QN(n5055) );
  NAND2X0 U7196 ( .IN1(P1_N374), .IN2(P1_N5582), .QN(n5054) );
  NAND2X0 U7197 ( .IN1(n5056), .IN2(n5057), .QN(P1_N3787) );
  NAND2X0 U7198 ( .IN1(P1_N3728), .IN2(n5018), .QN(n5057) );
  NAND2X0 U7199 ( .IN1(P1_N373), .IN2(P1_N5582), .QN(n5056) );
  NAND2X0 U7200 ( .IN1(n5058), .IN2(n5059), .QN(P1_N3786) );
  NAND2X0 U7201 ( .IN1(P1_N3727), .IN2(n5018), .QN(n5059) );
  NAND2X0 U7202 ( .IN1(P1_N372), .IN2(P1_N5582), .QN(n5058) );
  NAND2X0 U7203 ( .IN1(n5060), .IN2(n5061), .QN(P1_N3785) );
  NAND2X0 U7204 ( .IN1(P1_N3726), .IN2(n5018), .QN(n5061) );
  NAND2X0 U7205 ( .IN1(P1_N371), .IN2(P1_N5582), .QN(n5060) );
  NAND2X0 U7206 ( .IN1(n5062), .IN2(n5063), .QN(P1_N3784) );
  NAND2X0 U7207 ( .IN1(P1_N3725), .IN2(n5018), .QN(n5063) );
  NAND2X0 U7208 ( .IN1(P1_N370), .IN2(P1_N5582), .QN(n5062) );
  NAND2X0 U7209 ( .IN1(n5064), .IN2(n5065), .QN(P1_N3783) );
  NAND2X0 U7210 ( .IN1(P1_N3724), .IN2(n5018), .QN(n5065) );
  NAND2X0 U7211 ( .IN1(P1_N369), .IN2(P1_N5582), .QN(n5064) );
  NAND2X0 U7212 ( .IN1(n5066), .IN2(n5067), .QN(P1_N3782) );
  NAND2X0 U7213 ( .IN1(P1_N3723), .IN2(n5018), .QN(n5067) );
  NAND2X0 U7214 ( .IN1(P1_N368), .IN2(P1_N5582), .QN(n5066) );
  NAND2X0 U7215 ( .IN1(n5068), .IN2(n5069), .QN(P1_N3781) );
  NAND2X0 U7216 ( .IN1(P1_N3722), .IN2(n5018), .QN(n5069) );
  NAND2X0 U7217 ( .IN1(n18451), .IN2(P1_N5582), .QN(n5068) );
  NAND2X0 U7218 ( .IN1(n5070), .IN2(n5071), .QN(P1_N3780) );
  NAND2X0 U7219 ( .IN1(P1_N3721), .IN2(n5018), .QN(n5071) );
  NAND2X0 U7220 ( .IN1(n6623), .IN2(P1_N5582), .QN(n5070) );
  NAND2X0 U7221 ( .IN1(n5072), .IN2(n5073), .QN(P1_N3779) );
  NAND2X0 U7222 ( .IN1(P1_N3720), .IN2(n5018), .QN(n5073) );
  NAND2X0 U7223 ( .IN1(n6622), .IN2(P1_N5582), .QN(n5072) );
  NAND2X0 U7224 ( .IN1(n5074), .IN2(n5075), .QN(P1_N3778) );
  NAND2X0 U7225 ( .IN1(P1_N3719), .IN2(n5018), .QN(n5075) );
  NAND2X0 U7228 ( .IN1(n6621), .IN2(P1_N5582), .QN(n5074) );
  NAND2X0 U7233 ( .IN1(n7370), .IN2(n5078), .QN(P1_N3626) );
  NAND2X0 U7035 ( .IN1(P1_N4105), .IN2(n4932), .QN(n4963) );
  NAND2X0 U7036 ( .IN1(P1_N377), .IN2(P1_N5583), .QN(n4962) );
  NAND2X0 U7037 ( .IN1(n4964), .IN2(n4965), .QN(P1_N4163) );
  NAND2X0 U7038 ( .IN1(P1_N4104), .IN2(n4932), .QN(n4965) );
  NAND2X0 U7039 ( .IN1(P1_N376), .IN2(P1_N5583), .QN(n4964) );
  NAND2X0 U7040 ( .IN1(n4966), .IN2(n4967), .QN(P1_N4162) );
  NAND2X0 U7041 ( .IN1(P1_N4103), .IN2(n4932), .QN(n4967) );
  NAND2X0 U7042 ( .IN1(P1_N375), .IN2(P1_N5583), .QN(n4966) );
  NAND2X0 U7043 ( .IN1(n4968), .IN2(n4969), .QN(P1_N4161) );
  NAND2X0 U7044 ( .IN1(P1_N4102), .IN2(n4932), .QN(n4969) );
  NAND2X0 U7045 ( .IN1(P1_N374), .IN2(P1_N5583), .QN(n4968) );
  NAND2X0 U7046 ( .IN1(n4970), .IN2(n4971), .QN(P1_N4160) );
  NAND2X0 U7047 ( .IN1(P1_N4101), .IN2(n4932), .QN(n4971) );
  NAND2X0 U7048 ( .IN1(P1_N373), .IN2(P1_N5583), .QN(n4970) );
  NAND2X0 U7049 ( .IN1(n4972), .IN2(n4973), .QN(P1_N4159) );
  NAND2X0 U7050 ( .IN1(P1_N4100), .IN2(n4932), .QN(n4973) );
  NAND2X0 U7051 ( .IN1(P1_N372), .IN2(P1_N5583), .QN(n4972) );
  NAND2X0 U7052 ( .IN1(n4974), .IN2(n4975), .QN(P1_N4158) );
  NAND2X0 U7053 ( .IN1(P1_N4099), .IN2(n4932), .QN(n4975) );
  NAND2X0 U7054 ( .IN1(P1_N371), .IN2(P1_N5583), .QN(n4974) );
  NAND2X0 U7055 ( .IN1(n4976), .IN2(n4977), .QN(P1_N4157) );
  NAND2X0 U7056 ( .IN1(P1_N4098), .IN2(n4932), .QN(n4977) );
  NAND2X0 U7057 ( .IN1(P1_N370), .IN2(P1_N5583), .QN(n4976) );
  NAND2X0 U7058 ( .IN1(n4978), .IN2(n4979), .QN(P1_N4156) );
  NAND2X0 U7059 ( .IN1(P1_N4097), .IN2(n4932), .QN(n4979) );
  NAND2X0 U7060 ( .IN1(P1_N369), .IN2(P1_N5583), .QN(n4978) );
  NAND2X0 U7061 ( .IN1(n4980), .IN2(n4981), .QN(P1_N4155) );
  NAND2X0 U7062 ( .IN1(P1_N4096), .IN2(n4932), .QN(n4981) );
  NAND2X0 U7063 ( .IN1(P1_N368), .IN2(P1_N5583), .QN(n4980) );
  NAND2X0 U7064 ( .IN1(n4982), .IN2(n4983), .QN(P1_N4154) );
  NAND2X0 U7065 ( .IN1(P1_N4095), .IN2(n4932), .QN(n4983) );
  NAND2X0 U7066 ( .IN1(n18451), .IN2(P1_N5583), .QN(n4982) );
  NAND2X0 U7067 ( .IN1(n4984), .IN2(n4985), .QN(P1_N4153) );
  NAND2X0 U7068 ( .IN1(P1_N4094), .IN2(n4932), .QN(n4985) );
  NAND2X0 U7069 ( .IN1(n6623), .IN2(P1_N5583), .QN(n4984) );
  NAND2X0 U7070 ( .IN1(n4986), .IN2(n4987), .QN(P1_N4152) );
  NAND2X0 U7071 ( .IN1(P1_N4093), .IN2(n4932), .QN(n4987) );
  NAND2X0 U7072 ( .IN1(n6622), .IN2(P1_N5583), .QN(n4986) );
  NAND2X0 U7073 ( .IN1(n4988), .IN2(n4989), .QN(P1_N4151) );
  NAND2X0 U7074 ( .IN1(P1_N4092), .IN2(n4932), .QN(n4989) );
  NAND2X0 U7077 ( .IN1(n6621), .IN2(P1_N5583), .QN(n4988) );
  NAND2X0 U7082 ( .IN1(n7372), .IN2(n4992), .QN(P1_N3999) );
  NAND2X0 U7083 ( .IN1(n7371), .IN2(n4993), .QN(P1_N3997) );
  NOR2X0 U7084 ( .QN(P1_N4180), .IN1(n4993), .IN2(n4992) );
  INVX0 U7085 ( .ZN(n4992), .INP(n7371) );
  INVX0 U7086 ( .ZN(n4993), .INP(n7372) );
  NOR2X0 U7087 ( .QN(P1_N3879), .IN1(n7328), .IN2(n7023) );
  NOR2X0 U7088 ( .QN(P1_N3878), .IN1(n7326), .IN2(n7023) );
  NOR2X0 U7089 ( .QN(P1_N3877), .IN1(n7324), .IN2(n7021) );
  NOR2X0 U7090 ( .QN(P1_N3876), .IN1(n7322), .IN2(n7021) );
  NOR2X0 U7091 ( .QN(P1_N3875), .IN1(n7320), .IN2(n7021) );
  NOR2X0 U7092 ( .QN(P1_N3874), .IN1(n7318), .IN2(n7029) );
  NOR2X0 U7093 ( .QN(P1_N3873), .IN1(n7316), .IN2(n7029) );
  NOR2X0 U7094 ( .QN(P1_N3872), .IN1(n7314), .IN2(n7027) );
  NOR2X0 U7095 ( .QN(P1_N3871), .IN1(n7312), .IN2(n7027) );
  NOR2X0 U7096 ( .QN(P1_N3870), .IN1(n7310), .IN2(n7027) );
  NAND2X0 U7098 ( .IN1(n4097), .IN2(n4995), .QN(P1_N3869) );
  NAND2X0 U7099 ( .IN1(n7019), .IN2(n4099), .QN(n4995) );
  NAND2X0 U7100 ( .IN1(n4100), .IN2(n4996), .QN(P1_N3868) );
  NAND2X0 U7101 ( .IN1(n7028), .IN2(n4102), .QN(n4996) );
  NAND2X0 U7102 ( .IN1(n4103), .IN2(n4997), .QN(P1_N3867) );
  NAND2X0 U7103 ( .IN1(n7028), .IN2(n4105), .QN(n4997) );
  NAND2X0 U7104 ( .IN1(n4106), .IN2(n4998), .QN(P1_N3866) );
  NAND2X0 U7105 ( .IN1(n7028), .IN2(n4108), .QN(n4998) );
  NAND2X0 U7106 ( .IN1(n4109), .IN2(n4999), .QN(P1_N3865) );
  NAND2X0 U7107 ( .IN1(n7028), .IN2(n4111), .QN(n4999) );
  NAND2X0 U7108 ( .IN1(n4112), .IN2(n5000), .QN(P1_N3864) );
  NAND2X0 U7109 ( .IN1(n7024), .IN2(n4114), .QN(n5000) );
  NAND2X0 U7110 ( .IN1(n4115), .IN2(n5001), .QN(P1_N3863) );
  NAND2X0 U7111 ( .IN1(n7024), .IN2(n4117), .QN(n5001) );
  NAND2X0 U7112 ( .IN1(n4118), .IN2(n5002), .QN(P1_N3862) );
  NAND2X0 U7113 ( .IN1(n7024), .IN2(n4120), .QN(n5002) );
  NAND2X0 U7114 ( .IN1(n4121), .IN2(n5003), .QN(P1_N3861) );
  NAND2X0 U7115 ( .IN1(n7024), .IN2(n4123), .QN(n5003) );
  NAND2X0 U7116 ( .IN1(n4124), .IN2(n5004), .QN(P1_N3860) );
  NAND2X0 U7117 ( .IN1(n7024), .IN2(n4126), .QN(n5004) );
  NAND2X0 U7118 ( .IN1(n4127), .IN2(n5005), .QN(P1_N3859) );
  NAND2X0 U7119 ( .IN1(n7463), .IN2(n4129), .QN(n5005) );
  NAND2X0 U7120 ( .IN1(n4130), .IN2(n5006), .QN(P1_N3858) );
  NAND2X0 U7121 ( .IN1(n7463), .IN2(n4132), .QN(n5006) );
  NAND2X0 U7122 ( .IN1(n4133), .IN2(n5007), .QN(P1_N3857) );
  NAND2X0 U7123 ( .IN1(n7463), .IN2(n4135), .QN(n5007) );
  NAND2X0 U7124 ( .IN1(n4136), .IN2(n5008), .QN(P1_N3856) );
  NAND2X0 U7125 ( .IN1(n7463), .IN2(n4138), .QN(n5008) );
  NAND2X0 U7126 ( .IN1(n4139), .IN2(n5009), .QN(P1_N3855) );
  NAND2X0 U7127 ( .IN1(n7026), .IN2(n4141), .QN(n5009) );
  NAND2X0 U7128 ( .IN1(n4142), .IN2(n5010), .QN(P1_N3854) );
  NAND2X0 U7129 ( .IN1(n7026), .IN2(n4144), .QN(n5010) );
  NAND2X0 U7130 ( .IN1(n4145), .IN2(n5011), .QN(P1_N3853) );
  NAND2X0 U7131 ( .IN1(n7026), .IN2(n4147), .QN(n5011) );
  NAND2X0 U7132 ( .IN1(n4148), .IN2(n5012), .QN(P1_N3852) );
  NAND2X0 U7133 ( .IN1(n7022), .IN2(n4150), .QN(n5012) );
  NOR2X0 U6939 ( .QN(P1_N4249), .IN1(n7322), .IN2(n7021) );
  NOR2X0 U6940 ( .QN(P1_N4248), .IN1(n7320), .IN2(n7021) );
  NOR2X0 U6941 ( .QN(P1_N4247), .IN1(n7318), .IN2(n7021) );
  NOR2X0 U6942 ( .QN(P1_N4246), .IN1(n7316), .IN2(n7029) );
  NOR2X0 U6943 ( .QN(P1_N4245), .IN1(n7314), .IN2(n7027) );
  NOR2X0 U6944 ( .QN(P1_N4244), .IN1(n7312), .IN2(n7027) );
  NOR2X0 U6945 ( .QN(P1_N4243), .IN1(n7310), .IN2(n7021) );
  NAND2X0 U6947 ( .IN1(n4097), .IN2(n4909), .QN(P1_N4242) );
  NAND2X0 U6948 ( .IN1(n7019), .IN2(n4099), .QN(n4909) );
  NAND2X0 U6949 ( .IN1(n4100), .IN2(n4910), .QN(P1_N4241) );
  NAND2X0 U6950 ( .IN1(n7019), .IN2(n4102), .QN(n4910) );
  NAND2X0 U6951 ( .IN1(n4103), .IN2(n4911), .QN(P1_N4240) );
  NAND2X0 U6952 ( .IN1(n7028), .IN2(n4105), .QN(n4911) );
  NAND2X0 U6953 ( .IN1(n4106), .IN2(n4912), .QN(P1_N4239) );
  NAND2X0 U6954 ( .IN1(n7028), .IN2(n4108), .QN(n4912) );
  NAND2X0 U6955 ( .IN1(n4109), .IN2(n4913), .QN(P1_N4238) );
  NAND2X0 U6956 ( .IN1(n7028), .IN2(n4111), .QN(n4913) );
  NAND2X0 U6957 ( .IN1(n4112), .IN2(n4914), .QN(P1_N4237) );
  NAND2X0 U6958 ( .IN1(n7024), .IN2(n4114), .QN(n4914) );
  NAND2X0 U6959 ( .IN1(n4115), .IN2(n4915), .QN(P1_N4236) );
  NAND2X0 U6960 ( .IN1(n7024), .IN2(n4117), .QN(n4915) );
  NAND2X0 U6961 ( .IN1(n4118), .IN2(n4916), .QN(P1_N4235) );
  NAND2X0 U6962 ( .IN1(n7024), .IN2(n4120), .QN(n4916) );
  NAND2X0 U6963 ( .IN1(n4121), .IN2(n4917), .QN(P1_N4234) );
  NAND2X0 U6964 ( .IN1(n7024), .IN2(n4123), .QN(n4917) );
  NAND2X0 U6965 ( .IN1(n4124), .IN2(n4918), .QN(P1_N4233) );
  NAND2X0 U6966 ( .IN1(n7024), .IN2(n4126), .QN(n4918) );
  NAND2X0 U6967 ( .IN1(n4127), .IN2(n4919), .QN(P1_N4232) );
  NAND2X0 U6968 ( .IN1(n7463), .IN2(n4129), .QN(n4919) );
  NAND2X0 U6969 ( .IN1(n4130), .IN2(n4920), .QN(P1_N4231) );
  NAND2X0 U6970 ( .IN1(n7463), .IN2(n4132), .QN(n4920) );
  NAND2X0 U6971 ( .IN1(n4133), .IN2(n4921), .QN(P1_N4230) );
  NAND2X0 U6972 ( .IN1(n7463), .IN2(n4135), .QN(n4921) );
  NAND2X0 U6973 ( .IN1(n4136), .IN2(n4922), .QN(P1_N4229) );
  NAND2X0 U6974 ( .IN1(n7463), .IN2(n4138), .QN(n4922) );
  NAND2X0 U6975 ( .IN1(n4139), .IN2(n4923), .QN(P1_N4228) );
  NAND2X0 U6976 ( .IN1(n7026), .IN2(n4141), .QN(n4923) );
  NAND2X0 U6977 ( .IN1(n4142), .IN2(n4924), .QN(P1_N4227) );
  NAND2X0 U6978 ( .IN1(n7026), .IN2(n4144), .QN(n4924) );
  NAND2X0 U6979 ( .IN1(n4145), .IN2(n4925), .QN(P1_N4226) );
  NAND2X0 U6980 ( .IN1(n7026), .IN2(n4147), .QN(n4925) );
  NAND2X0 U6981 ( .IN1(n4148), .IN2(n4926), .QN(P1_N4225) );
  NAND2X0 U6982 ( .IN1(n7022), .IN2(n4150), .QN(n4926) );
  NAND2X0 U6983 ( .IN1(n4151), .IN2(n4927), .QN(P1_N4224) );
  NAND2X0 U6984 ( .IN1(n7022), .IN2(n4153), .QN(n4927) );
  NAND2X0 U6985 ( .IN1(n4154), .IN2(n4928), .QN(P1_N4223) );
  NAND2X0 U6986 ( .IN1(n7022), .IN2(n4156), .QN(n4928) );
  NAND2X0 U6989 ( .IN1(n4930), .IN2(n4931), .QN(P1_N4179) );
  NAND2X0 U6990 ( .IN1(P1_N4120), .IN2(n4932), .QN(n4931) );
  NAND2X0 U6991 ( .IN1(P1_N392), .IN2(P1_N5583), .QN(n4930) );
  NAND2X0 U6992 ( .IN1(n4934), .IN2(n4935), .QN(P1_N4178) );
  NAND2X0 U6993 ( .IN1(P1_N4119), .IN2(n4932), .QN(n4935) );
  NAND2X0 U6994 ( .IN1(P1_N391), .IN2(P1_N5583), .QN(n4934) );
  NAND2X0 U6995 ( .IN1(n4936), .IN2(n4937), .QN(P1_N4177) );
  NAND2X0 U6996 ( .IN1(P1_N4118), .IN2(n4932), .QN(n4937) );
  NAND2X0 U6997 ( .IN1(P1_N390), .IN2(P1_N5583), .QN(n4936) );
  NAND2X0 U6998 ( .IN1(n4938), .IN2(n4939), .QN(P1_N4176) );
  NAND2X0 U6999 ( .IN1(P1_N4117), .IN2(n4932), .QN(n4939) );
  NAND2X0 U7000 ( .IN1(P1_N389), .IN2(P1_N5583), .QN(n4938) );
  NAND2X0 U7001 ( .IN1(n4940), .IN2(n4941), .QN(P1_N4175) );
  NAND2X0 U7002 ( .IN1(P1_N4116), .IN2(n4932), .QN(n4941) );
  NAND2X0 U7003 ( .IN1(P1_N388), .IN2(P1_N5583), .QN(n4940) );
  NAND2X0 U7004 ( .IN1(n4942), .IN2(n4943), .QN(P1_N4174) );
  NAND2X0 U7005 ( .IN1(P1_N4115), .IN2(n4932), .QN(n4943) );
  NAND2X0 U7006 ( .IN1(P1_N387), .IN2(P1_N5583), .QN(n4942) );
  NAND2X0 U7007 ( .IN1(n4944), .IN2(n4945), .QN(P1_N4173) );
  NAND2X0 U7008 ( .IN1(P1_N4114), .IN2(n4932), .QN(n4945) );
  NAND2X0 U7009 ( .IN1(P1_N386), .IN2(P1_N5583), .QN(n4944) );
  NAND2X0 U7010 ( .IN1(n4946), .IN2(n4947), .QN(P1_N4172) );
  NAND2X0 U7011 ( .IN1(P1_N4113), .IN2(n4932), .QN(n4947) );
  NAND2X0 U7012 ( .IN1(P1_N385), .IN2(P1_N5583), .QN(n4946) );
  NAND2X0 U7013 ( .IN1(n4948), .IN2(n4949), .QN(P1_N4171) );
  NAND2X0 U7014 ( .IN1(P1_N4112), .IN2(n4932), .QN(n4949) );
  NAND2X0 U7015 ( .IN1(P1_N384), .IN2(P1_N5583), .QN(n4948) );
  NAND2X0 U7016 ( .IN1(n4950), .IN2(n4951), .QN(P1_N4170) );
  NAND2X0 U7017 ( .IN1(P1_N4111), .IN2(n4932), .QN(n4951) );
  NAND2X0 U7018 ( .IN1(P1_N383), .IN2(P1_N5583), .QN(n4950) );
  NAND2X0 U7019 ( .IN1(n4952), .IN2(n4953), .QN(P1_N4169) );
  NAND2X0 U7020 ( .IN1(P1_N4110), .IN2(n4932), .QN(n4953) );
  NAND2X0 U7021 ( .IN1(P1_N382), .IN2(P1_N5583), .QN(n4952) );
  NAND2X0 U7022 ( .IN1(n4954), .IN2(n4955), .QN(P1_N4168) );
  NAND2X0 U7023 ( .IN1(P1_N4109), .IN2(n4932), .QN(n4955) );
  NAND2X0 U7024 ( .IN1(P1_N381), .IN2(P1_N5583), .QN(n4954) );
  NAND2X0 U7025 ( .IN1(n4956), .IN2(n4957), .QN(P1_N4167) );
  NAND2X0 U7026 ( .IN1(P1_N4108), .IN2(n4932), .QN(n4957) );
  NAND2X0 U7027 ( .IN1(P1_N380), .IN2(P1_N5583), .QN(n4956) );
  NAND2X0 U7028 ( .IN1(n4958), .IN2(n4959), .QN(P1_N4166) );
  NAND2X0 U7029 ( .IN1(P1_N4107), .IN2(n4932), .QN(n4959) );
  NAND2X0 U7030 ( .IN1(P1_N379), .IN2(P1_N5583), .QN(n4958) );
  NAND2X0 U7031 ( .IN1(n4960), .IN2(n4961), .QN(P1_N4165) );
  NAND2X0 U7032 ( .IN1(P1_N4106), .IN2(n4932), .QN(n4961) );
  NAND2X0 U7033 ( .IN1(P1_N378), .IN2(P1_N5583), .QN(n4960) );
  NAND2X0 U7034 ( .IN1(n4962), .IN2(n4963), .QN(P1_N4164) );
  NAND2X0 U6841 ( .IN1(n4847), .IN2(n4848), .QN(n4840) );
  AND2X1 U6842 ( .IN1(n4849), .IN2(n4850), .Q(n4848) );
  NOR2X0 U6843 ( .QN(n4850), .IN1(P1_N411), .IN2(P1_N410) );
  NOR2X0 U6844 ( .QN(n4849), .IN1(P1_N409), .IN2(P1_N408) );
  NOR2X0 U6845 ( .QN(n4847), .IN1(P1_N405), .IN2(n4851) );
  OR2X1 U6846 ( .IN2(P1_N406), .IN1(P1_N407), .Q(n4851) );
  NAND2X0 U6847 ( .IN1(n4852), .IN2(n4853), .QN(P1_N4549) );
  NAND2X0 U6848 ( .IN1(P1_N4490), .IN2(n4818), .QN(n4853) );
  NAND2X0 U6849 ( .IN1(P1_N389), .IN2(P1_N5584), .QN(n4852) );
  NAND2X0 U6850 ( .IN1(n4854), .IN2(n4855), .QN(P1_N4548) );
  NAND2X0 U6851 ( .IN1(P1_N4489), .IN2(n4818), .QN(n4855) );
  NAND2X0 U6852 ( .IN1(P1_N388), .IN2(P1_N5584), .QN(n4854) );
  NAND2X0 U6853 ( .IN1(n4856), .IN2(n4857), .QN(P1_N4547) );
  NAND2X0 U6854 ( .IN1(P1_N4488), .IN2(n4818), .QN(n4857) );
  NAND2X0 U6855 ( .IN1(P1_N387), .IN2(P1_N5584), .QN(n4856) );
  NAND2X0 U6856 ( .IN1(n4858), .IN2(n4859), .QN(P1_N4546) );
  NAND2X0 U6857 ( .IN1(P1_N4487), .IN2(n4818), .QN(n4859) );
  NAND2X0 U6858 ( .IN1(P1_N386), .IN2(P1_N5584), .QN(n4858) );
  NAND2X0 U6859 ( .IN1(n4860), .IN2(n4861), .QN(P1_N4545) );
  NAND2X0 U6860 ( .IN1(P1_N4486), .IN2(n4818), .QN(n4861) );
  NAND2X0 U6861 ( .IN1(P1_N385), .IN2(P1_N5584), .QN(n4860) );
  NAND2X0 U6862 ( .IN1(n4862), .IN2(n4863), .QN(P1_N4544) );
  NAND2X0 U6863 ( .IN1(P1_N4485), .IN2(n4818), .QN(n4863) );
  NAND2X0 U6864 ( .IN1(P1_N384), .IN2(P1_N5584), .QN(n4862) );
  NAND2X0 U6865 ( .IN1(n4864), .IN2(n4865), .QN(P1_N4543) );
  NAND2X0 U6866 ( .IN1(P1_N4484), .IN2(n4818), .QN(n4865) );
  NAND2X0 U6867 ( .IN1(P1_N383), .IN2(P1_N5584), .QN(n4864) );
  NAND2X0 U6868 ( .IN1(n4866), .IN2(n4867), .QN(P1_N4542) );
  NAND2X0 U6869 ( .IN1(P1_N4483), .IN2(n4818), .QN(n4867) );
  NAND2X0 U6870 ( .IN1(P1_N382), .IN2(P1_N5584), .QN(n4866) );
  NAND2X0 U6871 ( .IN1(n4868), .IN2(n4869), .QN(P1_N4541) );
  NAND2X0 U6872 ( .IN1(P1_N4482), .IN2(n4818), .QN(n4869) );
  NAND2X0 U6873 ( .IN1(P1_N381), .IN2(P1_N5584), .QN(n4868) );
  NAND2X0 U6874 ( .IN1(n4870), .IN2(n4871), .QN(P1_N4540) );
  NAND2X0 U6875 ( .IN1(P1_N4481), .IN2(n4818), .QN(n4871) );
  NAND2X0 U6876 ( .IN1(P1_N380), .IN2(P1_N5584), .QN(n4870) );
  NAND2X0 U6877 ( .IN1(n4872), .IN2(n4873), .QN(P1_N4539) );
  NAND2X0 U6878 ( .IN1(P1_N4480), .IN2(n4818), .QN(n4873) );
  NAND2X0 U6879 ( .IN1(P1_N379), .IN2(P1_N5584), .QN(n4872) );
  NAND2X0 U6880 ( .IN1(n4874), .IN2(n4875), .QN(P1_N4538) );
  NAND2X0 U6881 ( .IN1(P1_N4479), .IN2(n4818), .QN(n4875) );
  NAND2X0 U6882 ( .IN1(P1_N378), .IN2(P1_N5584), .QN(n4874) );
  NAND2X0 U6883 ( .IN1(n4876), .IN2(n4877), .QN(P1_N4537) );
  NAND2X0 U6884 ( .IN1(P1_N4478), .IN2(n4818), .QN(n4877) );
  NAND2X0 U6885 ( .IN1(P1_N377), .IN2(P1_N5584), .QN(n4876) );
  NAND2X0 U6886 ( .IN1(n4878), .IN2(n4879), .QN(P1_N4536) );
  NAND2X0 U6887 ( .IN1(P1_N4477), .IN2(n4818), .QN(n4879) );
  NAND2X0 U6888 ( .IN1(P1_N376), .IN2(P1_N5584), .QN(n4878) );
  NAND2X0 U6889 ( .IN1(n4880), .IN2(n4881), .QN(P1_N4535) );
  NAND2X0 U6890 ( .IN1(P1_N4476), .IN2(n4818), .QN(n4881) );
  NAND2X0 U6891 ( .IN1(P1_N375), .IN2(P1_N5584), .QN(n4880) );
  NAND2X0 U6892 ( .IN1(n4882), .IN2(n4883), .QN(P1_N4534) );
  NAND2X0 U6893 ( .IN1(P1_N4475), .IN2(n4818), .QN(n4883) );
  NAND2X0 U6894 ( .IN1(P1_N374), .IN2(P1_N5584), .QN(n4882) );
  NAND2X0 U6895 ( .IN1(n4884), .IN2(n4885), .QN(P1_N4533) );
  NAND2X0 U6896 ( .IN1(P1_N4474), .IN2(n4818), .QN(n4885) );
  NAND2X0 U6897 ( .IN1(P1_N373), .IN2(P1_N5584), .QN(n4884) );
  NAND2X0 U6898 ( .IN1(n4886), .IN2(n4887), .QN(P1_N4532) );
  NAND2X0 U6899 ( .IN1(P1_N4473), .IN2(n4818), .QN(n4887) );
  NAND2X0 U6900 ( .IN1(P1_N372), .IN2(P1_N5584), .QN(n4886) );
  NAND2X0 U6901 ( .IN1(n4888), .IN2(n4889), .QN(P1_N4531) );
  NAND2X0 U6902 ( .IN1(P1_N4472), .IN2(n4818), .QN(n4889) );
  NAND2X0 U6903 ( .IN1(P1_N371), .IN2(P1_N5584), .QN(n4888) );
  NAND2X0 U6904 ( .IN1(n4890), .IN2(n4891), .QN(P1_N4530) );
  NAND2X0 U6905 ( .IN1(P1_N4471), .IN2(n4818), .QN(n4891) );
  NAND2X0 U6906 ( .IN1(P1_N370), .IN2(P1_N5584), .QN(n4890) );
  NAND2X0 U6907 ( .IN1(n4892), .IN2(n4893), .QN(P1_N4529) );
  NAND2X0 U6908 ( .IN1(P1_N4470), .IN2(n4818), .QN(n4893) );
  NAND2X0 U6909 ( .IN1(P1_N369), .IN2(P1_N5584), .QN(n4892) );
  NAND2X0 U6910 ( .IN1(n4894), .IN2(n4895), .QN(P1_N4528) );
  NAND2X0 U6911 ( .IN1(P1_N4469), .IN2(n4818), .QN(n4895) );
  NAND2X0 U6912 ( .IN1(P1_N368), .IN2(P1_N5584), .QN(n4894) );
  NAND2X0 U6913 ( .IN1(n4896), .IN2(n4897), .QN(P1_N4527) );
  NAND2X0 U6914 ( .IN1(P1_N4468), .IN2(n4818), .QN(n4897) );
  NAND2X0 U6915 ( .IN1(n18451), .IN2(P1_N5584), .QN(n4896) );
  NAND2X0 U6916 ( .IN1(n4898), .IN2(n4899), .QN(P1_N4526) );
  NAND2X0 U6917 ( .IN1(P1_N4467), .IN2(n4818), .QN(n4899) );
  NAND2X0 U6918 ( .IN1(n6623), .IN2(P1_N5584), .QN(n4898) );
  NAND2X0 U6919 ( .IN1(n4900), .IN2(n4901), .QN(P1_N4525) );
  NAND2X0 U6920 ( .IN1(P1_N4466), .IN2(n4818), .QN(n4901) );
  NAND2X0 U6921 ( .IN1(n6622), .IN2(P1_N5584), .QN(n4900) );
  NAND2X0 U6922 ( .IN1(n4902), .IN2(n4903), .QN(P1_N4524) );
  NAND2X0 U6923 ( .IN1(P1_N4465), .IN2(n4818), .QN(n4903) );
  NAND2X0 U6926 ( .IN1(n6621), .IN2(P1_N5584), .QN(n4902) );
  NAND2X0 U6931 ( .IN1(n7374), .IN2(n4906), .QN(P1_N4372) );
  NAND2X0 U6932 ( .IN1(n7373), .IN2(n4907), .QN(P1_N4370) );
  NOR2X0 U6933 ( .QN(P1_N4553), .IN1(n4907), .IN2(n4906) );
  INVX0 U6934 ( .ZN(n4906), .INP(n7373) );
  INVX0 U6935 ( .ZN(n4907), .INP(n7374) );
  NOR2X0 U6936 ( .QN(P1_N4252), .IN1(n7328), .IN2(n7023) );
  NOR2X0 U6937 ( .QN(P1_N4251), .IN1(n7326), .IN2(n7023) );
  NOR2X0 U6938 ( .QN(P1_N4250), .IN1(n7324), .IN2(n7021) );
  OR2X1 U6744 ( .IN2(n4772), .IN1(n4771), .Q(P1_N5153) );
  NAND2X0 U6745 ( .IN1(n4773), .IN2(n4774), .QN(n4772) );
  NAND2X0 U6746 ( .IN1(n9749), .IN2(n7344), .QN(n4774) );
  NAND2X0 U6747 ( .IN1(n9821), .IN2(n7345), .QN(n4773) );
  NAND2X0 U6748 ( .IN1(n4775), .IN2(n4776), .QN(n4771) );
  NAND2X0 U6749 ( .IN1(n8990), .IN2(n4480), .QN(n4776) );
  NAND2X0 U6750 ( .IN1(n7347), .IN2(P1_N368), .QN(n4775) );
  NAND2X0 U6752 ( .IN1(n4777), .IN2(n4778), .QN(P1_N4629) );
  NAND2X0 U6753 ( .IN1(P1_N4561), .IN2(n4584), .QN(n4778) );
  NAND2X0 U6754 ( .IN1(P1_N5571), .IN2(n7041), .QN(n4777) );
  OR2X1 U6755 ( .IN2(n4780), .IN1(n4779), .Q(P1_N5152) );
  NAND2X0 U6756 ( .IN1(n4781), .IN2(n4782), .QN(n4780) );
  NAND2X0 U6757 ( .IN1(n9753), .IN2(n7344), .QN(n4782) );
  NAND2X0 U6758 ( .IN1(n9825), .IN2(n7345), .QN(n4781) );
  NAND2X0 U6759 ( .IN1(n4783), .IN2(n4784), .QN(n4779) );
  NAND2X0 U6760 ( .IN1(n8994), .IN2(n4480), .QN(n4784) );
  NAND2X0 U6761 ( .IN1(n7347), .IN2(n18451), .QN(n4783) );
  NAND2X0 U6762 ( .IN1(n4785), .IN2(n4786), .QN(P1_N4628) );
  NAND2X0 U6763 ( .IN1(P1_N4560), .IN2(n4584), .QN(n4786) );
  NAND2X0 U6764 ( .IN1(P1_N5571), .IN2(n7046), .QN(n4785) );
  OR2X1 U6765 ( .IN2(n4788), .IN1(n4787), .Q(P1_N5151) );
  NAND2X0 U6766 ( .IN1(n4789), .IN2(n4790), .QN(n4788) );
  NAND2X0 U6767 ( .IN1(n9757), .IN2(n7344), .QN(n4790) );
  NAND2X0 U6768 ( .IN1(n9829), .IN2(n7345), .QN(n4789) );
  NAND2X0 U6769 ( .IN1(n4791), .IN2(n4792), .QN(n4787) );
  NAND2X0 U6770 ( .IN1(n8998), .IN2(n4480), .QN(n4792) );
  NAND2X0 U6771 ( .IN1(n7347), .IN2(n6623), .QN(n4791) );
  NAND2X0 U6772 ( .IN1(n4793), .IN2(n4794), .QN(P1_N4627) );
  NAND2X0 U6773 ( .IN1(P1_N4559), .IN2(n4584), .QN(n4794) );
  NAND2X0 U6774 ( .IN1(P1_N5571), .IN2(P1_N5150), .QN(n4793) );
  OR2X1 U6775 ( .IN2(n4796), .IN1(n4795), .Q(P1_N5150) );
  NAND2X0 U6776 ( .IN1(n4797), .IN2(n4798), .QN(n4796) );
  NAND2X0 U6777 ( .IN1(n9761), .IN2(n7344), .QN(n4798) );
  NAND2X0 U6778 ( .IN1(n9833), .IN2(n7345), .QN(n4797) );
  NAND2X0 U6779 ( .IN1(n4799), .IN2(n4800), .QN(n4795) );
  NAND2X0 U6780 ( .IN1(n9002), .IN2(n4480), .QN(n4800) );
  NAND2X0 U6781 ( .IN1(n7347), .IN2(n6622), .QN(n4799) );
  NAND2X0 U6782 ( .IN1(n4801), .IN2(n4802), .QN(P1_N4626) );
  NAND2X0 U6783 ( .IN1(P1_N4558), .IN2(n4584), .QN(n4802) );
  NAND2X0 U6784 ( .IN1(P1_N5571), .IN2(n7034), .QN(n4801) );
  AND2X1 U6786 ( .IN1(P1_N4557), .IN2(n4584), .Q(P1_N4625) );
  OR2X1 U6787 ( .IN2(P1_N583), .IN1(n6996), .Q(n4584) );
  NOR2X0 U6789 ( .QN(P1_N4556), .IN1(n4469), .IN2(n4803) );
  NAND2X0 U6791 ( .IN1(n4806), .IN2(n4807), .QN(n4805) );
  NAND2X0 U6792 ( .IN1(n981), .IN2(n7344), .QN(n4807) );
  NAND2X0 U6793 ( .IN1(n920), .IN2(n7345), .QN(n4806) );
  NAND2X0 U6794 ( .IN1(n4808), .IN2(n4809), .QN(n4804) );
  NAND2X0 U6795 ( .IN1(n9006), .IN2(n4480), .QN(n4809) );
  NAND2X0 U6796 ( .IN1(n7347), .IN2(n6621), .QN(n4808) );
  NOR2X0 U6797 ( .QN(n4469), .IN1(n7349), .IN2(n4811) );
  NAND2X0 U6798 ( .IN1(n4812), .IN2(n4813), .QN(n4811) );
  NAND2X0 U6799 ( .IN1(n9010), .IN2(n7344), .QN(n4813) );
  NAND2X0 U6800 ( .IN1(n8886), .IN2(n7345), .QN(n4812) );
  INVX0 U6804 ( .ZN(n4616), .INP(n7335) );
  INVX0 U6805 ( .ZN(n4615), .INP(n7336) );
  NAND2X0 U6809 ( .IN1(n4816), .IN2(n4817), .QN(P1_N4552) );
  NAND2X0 U6810 ( .IN1(P1_N4493), .IN2(n4818), .QN(n4817) );
  NAND2X0 U6811 ( .IN1(P1_N392), .IN2(P1_N5584), .QN(n4816) );
  NAND2X0 U6812 ( .IN1(n4820), .IN2(n4821), .QN(P1_N4551) );
  NAND2X0 U6813 ( .IN1(P1_N4492), .IN2(n4818), .QN(n4821) );
  NAND2X0 U6814 ( .IN1(P1_N391), .IN2(P1_N5584), .QN(n4820) );
  NAND2X0 U6815 ( .IN1(n4822), .IN2(n4823), .QN(P1_N4550) );
  NAND2X0 U6816 ( .IN1(P1_N4491), .IN2(n4818), .QN(n4823) );
  NAND2X0 U6817 ( .IN1(P1_N390), .IN2(P1_N5584), .QN(n4822) );
  AND2X1 U6818 ( .IN1(P1_N395), .IN2(n4824), .Q(P1_N455) );
  NAND2X0 U6819 ( .IN1(n4825), .IN2(n4826), .QN(n4824) );
  NOR2X0 U6820 ( .QN(n4826), .IN1(n4827), .IN2(n4828) );
  NAND2X0 U6821 ( .IN1(n4829), .IN2(n4830), .QN(n4828) );
  AND2X1 U6822 ( .IN1(n4831), .IN2(n4832), .Q(n4830) );
  NOR2X0 U6823 ( .QN(n4832), .IN1(P1_N418), .IN2(P1_N417) );
  NOR2X0 U6824 ( .QN(n4831), .IN1(P1_N416), .IN2(P1_N415) );
  NOR2X0 U6825 ( .QN(n4829), .IN1(P1_N412), .IN2(n4833) );
  OR2X1 U6826 ( .IN2(P1_N413), .IN1(P1_N414), .Q(n4833) );
  OR2X1 U6827 ( .IN2(n4835), .IN1(n4834), .Q(n4827) );
  NAND2X0 U6828 ( .IN1(n4836), .IN2(n4837), .QN(n4835) );
  NOR2X0 U6829 ( .QN(n4837), .IN1(P1_N422), .IN2(P1_N421) );
  NOR2X0 U6830 ( .QN(n4836), .IN1(P1_N420), .IN2(P1_N419) );
  NAND2X0 U6831 ( .IN1(n4838), .IN2(n4839), .QN(n4834) );
  NOR2X0 U6832 ( .QN(n4839), .IN1(P1_N426), .IN2(P1_N425) );
  NOR2X0 U6833 ( .QN(n4838), .IN1(P1_N424), .IN2(P1_N423) );
  NOR2X0 U6834 ( .QN(n4825), .IN1(n4840), .IN2(n4841) );
  NAND2X0 U6835 ( .IN1(n4842), .IN2(n4843), .QN(n4841) );
  AND2X1 U6836 ( .IN1(n4844), .IN2(n4845), .Q(n4843) );
  NOR2X0 U6837 ( .QN(n4845), .IN1(P1_N404), .IN2(P1_N403) );
  NOR2X0 U6838 ( .QN(n4844), .IN1(P1_N402), .IN2(P1_N401) );
  NOR2X0 U6839 ( .QN(n4842), .IN1(P1_N398), .IN2(n4846) );
  OR2X1 U6840 ( .IN2(P1_N399), .IN1(P1_N400), .Q(n4846) );
  NAND2X0 U6651 ( .IN1(n4697), .IN2(n4698), .QN(P1_N4639) );
  NAND2X0 U6652 ( .IN1(P1_N4571), .IN2(n4584), .QN(n4698) );
  NAND2X0 U6653 ( .IN1(P1_N5571), .IN2(n7055), .QN(n4697) );
  OR2X1 U6654 ( .IN2(n4700), .IN1(n4699), .Q(P1_N5162) );
  NAND2X0 U6655 ( .IN1(n4701), .IN2(n4702), .QN(n4700) );
  NAND2X0 U6656 ( .IN1(n9713), .IN2(n7344), .QN(n4702) );
  NAND2X0 U6657 ( .IN1(n9785), .IN2(n7345), .QN(n4701) );
  NAND2X0 U6658 ( .IN1(n4703), .IN2(n4704), .QN(n4699) );
  NAND2X0 U6659 ( .IN1(n8954), .IN2(n4480), .QN(n4704) );
  NAND2X0 U6660 ( .IN1(n7347), .IN2(P1_N377), .QN(n4703) );
  NAND2X0 U6661 ( .IN1(n4705), .IN2(n4706), .QN(P1_N4638) );
  NAND2X0 U6662 ( .IN1(P1_N4570), .IN2(n4584), .QN(n4706) );
  NAND2X0 U6663 ( .IN1(P1_N5571), .IN2(n7059), .QN(n4705) );
  OR2X1 U6664 ( .IN2(n4708), .IN1(n4707), .Q(P1_N5161) );
  NAND2X0 U6665 ( .IN1(n4709), .IN2(n4710), .QN(n4708) );
  NAND2X0 U6666 ( .IN1(n9717), .IN2(n7344), .QN(n4710) );
  NAND2X0 U6667 ( .IN1(n9789), .IN2(n7345), .QN(n4709) );
  NAND2X0 U6668 ( .IN1(n4711), .IN2(n4712), .QN(n4707) );
  NAND2X0 U6669 ( .IN1(n8958), .IN2(n4480), .QN(n4712) );
  NAND2X0 U6670 ( .IN1(n7347), .IN2(P1_N376), .QN(n4711) );
  NAND2X0 U6671 ( .IN1(n4713), .IN2(n4714), .QN(P1_N4637) );
  NAND2X0 U6672 ( .IN1(P1_N4569), .IN2(n4584), .QN(n4714) );
  NAND2X0 U6673 ( .IN1(P1_N5571), .IN2(n7062), .QN(n4713) );
  OR2X1 U6674 ( .IN2(n4716), .IN1(n4715), .Q(P1_N5160) );
  NAND2X0 U6675 ( .IN1(n4717), .IN2(n4718), .QN(n4716) );
  NAND2X0 U6676 ( .IN1(n9721), .IN2(n7344), .QN(n4718) );
  NAND2X0 U6677 ( .IN1(n9793), .IN2(n7345), .QN(n4717) );
  NAND2X0 U6678 ( .IN1(n4719), .IN2(n4720), .QN(n4715) );
  NAND2X0 U6679 ( .IN1(n8962), .IN2(n4480), .QN(n4720) );
  NAND2X0 U6680 ( .IN1(n7347), .IN2(P1_N375), .QN(n4719) );
  NAND2X0 U6681 ( .IN1(n4721), .IN2(n4722), .QN(P1_N4636) );
  NAND2X0 U6682 ( .IN1(P1_N4568), .IN2(n4584), .QN(n4722) );
  NAND2X0 U6683 ( .IN1(P1_N5571), .IN2(n7066), .QN(n4721) );
  OR2X1 U6684 ( .IN2(n4724), .IN1(n4723), .Q(P1_N5159) );
  NAND2X0 U6685 ( .IN1(n4725), .IN2(n4726), .QN(n4724) );
  NAND2X0 U6686 ( .IN1(n9725), .IN2(n7344), .QN(n4726) );
  NAND2X0 U6687 ( .IN1(n9797), .IN2(n7345), .QN(n4725) );
  NAND2X0 U6688 ( .IN1(n4727), .IN2(n4728), .QN(n4723) );
  NAND2X0 U6689 ( .IN1(n8966), .IN2(n4480), .QN(n4728) );
  NAND2X0 U6690 ( .IN1(n7347), .IN2(P1_N374), .QN(n4727) );
  NAND2X0 U6691 ( .IN1(n4729), .IN2(n4730), .QN(P1_N4635) );
  NAND2X0 U6692 ( .IN1(P1_N4567), .IN2(n4584), .QN(n4730) );
  NAND2X0 U6693 ( .IN1(P1_N5571), .IN2(n7070), .QN(n4729) );
  OR2X1 U6694 ( .IN2(n4732), .IN1(n4731), .Q(P1_N5158) );
  NAND2X0 U6695 ( .IN1(n4733), .IN2(n4734), .QN(n4732) );
  NAND2X0 U6696 ( .IN1(n9729), .IN2(n7344), .QN(n4734) );
  NAND2X0 U6697 ( .IN1(n9801), .IN2(n7345), .QN(n4733) );
  NAND2X0 U6698 ( .IN1(n4735), .IN2(n4736), .QN(n4731) );
  NAND2X0 U6699 ( .IN1(n8970), .IN2(n4480), .QN(n4736) );
  NAND2X0 U6700 ( .IN1(n7347), .IN2(P1_N373), .QN(n4735) );
  NAND2X0 U6701 ( .IN1(n4737), .IN2(n4738), .QN(P1_N4634) );
  NAND2X0 U6702 ( .IN1(P1_N4566), .IN2(n4584), .QN(n4738) );
  NAND2X0 U6703 ( .IN1(P1_N5571), .IN2(P1_N5157), .QN(n4737) );
  OR2X1 U6704 ( .IN2(n4740), .IN1(n4739), .Q(P1_N5157) );
  NAND2X0 U6705 ( .IN1(n4741), .IN2(n4742), .QN(n4740) );
  NAND2X0 U6706 ( .IN1(n9733), .IN2(n7344), .QN(n4742) );
  NAND2X0 U6707 ( .IN1(n9805), .IN2(n7345), .QN(n4741) );
  NAND2X0 U6708 ( .IN1(n4743), .IN2(n4744), .QN(n4739) );
  NAND2X0 U6709 ( .IN1(n8974), .IN2(n4480), .QN(n4744) );
  NAND2X0 U6710 ( .IN1(n7347), .IN2(P1_N372), .QN(n4743) );
  NAND2X0 U6711 ( .IN1(n4745), .IN2(n4746), .QN(P1_N4633) );
  NAND2X0 U6712 ( .IN1(P1_N4565), .IN2(n4584), .QN(n4746) );
  NAND2X0 U6713 ( .IN1(P1_N5571), .IN2(P1_N5156), .QN(n4745) );
  OR2X1 U6714 ( .IN2(n4748), .IN1(n4747), .Q(P1_N5156) );
  NAND2X0 U6715 ( .IN1(n4749), .IN2(n4750), .QN(n4748) );
  NAND2X0 U6716 ( .IN1(n9737), .IN2(n7344), .QN(n4750) );
  NAND2X0 U6717 ( .IN1(n9809), .IN2(n7345), .QN(n4749) );
  NAND2X0 U6718 ( .IN1(n4751), .IN2(n4752), .QN(n4747) );
  NAND2X0 U6719 ( .IN1(n8978), .IN2(n4480), .QN(n4752) );
  NAND2X0 U6720 ( .IN1(n7347), .IN2(P1_N371), .QN(n4751) );
  NAND2X0 U6721 ( .IN1(n4753), .IN2(n4754), .QN(P1_N4632) );
  NAND2X0 U6722 ( .IN1(P1_N4564), .IN2(n4584), .QN(n4754) );
  NAND2X0 U6723 ( .IN1(P1_N5571), .IN2(n7080), .QN(n4753) );
  OR2X1 U6724 ( .IN2(n4756), .IN1(n4755), .Q(P1_N5155) );
  NAND2X0 U6725 ( .IN1(n4757), .IN2(n4758), .QN(n4756) );
  NAND2X0 U6726 ( .IN1(n9741), .IN2(n7344), .QN(n4758) );
  NAND2X0 U6727 ( .IN1(n9813), .IN2(n7345), .QN(n4757) );
  NAND2X0 U6728 ( .IN1(n4759), .IN2(n4760), .QN(n4755) );
  NAND2X0 U6729 ( .IN1(n8982), .IN2(n4480), .QN(n4760) );
  NAND2X0 U6730 ( .IN1(n7347), .IN2(P1_N370), .QN(n4759) );
  NAND2X0 U6731 ( .IN1(n4761), .IN2(n4762), .QN(P1_N4631) );
  NAND2X0 U6732 ( .IN1(P1_N4563), .IN2(n4584), .QN(n4762) );
  NAND2X0 U6733 ( .IN1(P1_N5571), .IN2(n7081), .QN(n4761) );
  OR2X1 U6734 ( .IN2(n4764), .IN1(n4763), .Q(P1_N5154) );
  NAND2X0 U6735 ( .IN1(n4765), .IN2(n4766), .QN(n4764) );
  NAND2X0 U6736 ( .IN1(n9745), .IN2(n7344), .QN(n4766) );
  NAND2X0 U6737 ( .IN1(n9817), .IN2(n7345), .QN(n4765) );
  NAND2X0 U6738 ( .IN1(n4767), .IN2(n4768), .QN(n4763) );
  NAND2X0 U6739 ( .IN1(n8986), .IN2(n4480), .QN(n4768) );
  NAND2X0 U6740 ( .IN1(n7347), .IN2(P1_N369), .QN(n4767) );
  NAND2X0 U6741 ( .IN1(n4769), .IN2(n4770), .QN(P1_N4630) );
  NAND2X0 U6742 ( .IN1(P1_N4562), .IN2(n4584), .QN(n4770) );
  NAND2X0 U6743 ( .IN1(P1_N5571), .IN2(P1_N5153), .QN(n4769) );
  NAND2X0 U6558 ( .IN1(n4623), .IN2(n4624), .QN(n4619) );
  NAND2X0 U6559 ( .IN1(n8914), .IN2(n4480), .QN(n4624) );
  NAND2X0 U6560 ( .IN1(n7347), .IN2(P1_N387), .QN(n4623) );
  NAND2X0 U6561 ( .IN1(n4625), .IN2(n4626), .QN(P1_N4648) );
  NAND2X0 U6562 ( .IN1(P1_N4580), .IN2(n4584), .QN(n4626) );
  NAND2X0 U6563 ( .IN1(P1_N5571), .IN2(P1_N5171), .QN(n4625) );
  OR2X1 U6564 ( .IN2(n4628), .IN1(n4627), .Q(P1_N5171) );
  NAND2X0 U6565 ( .IN1(n4629), .IN2(n4630), .QN(n4628) );
  NAND2X0 U6566 ( .IN1(n9046), .IN2(n7344), .QN(n4630) );
  NAND2X0 U6567 ( .IN1(n9086), .IN2(n7345), .QN(n4629) );
  NAND2X0 U6568 ( .IN1(n4631), .IN2(n4632), .QN(n4627) );
  NAND2X0 U6569 ( .IN1(n8918), .IN2(n4480), .QN(n4632) );
  NAND2X0 U6570 ( .IN1(n7347), .IN2(P1_N386), .QN(n4631) );
  NAND2X0 U6571 ( .IN1(n4633), .IN2(n4634), .QN(P1_N4647) );
  NAND2X0 U6572 ( .IN1(P1_N4579), .IN2(n4584), .QN(n4634) );
  NAND2X0 U6573 ( .IN1(P1_N5571), .IN2(n7093), .QN(n4633) );
  OR2X1 U6574 ( .IN2(n4636), .IN1(n4635), .Q(P1_N5170) );
  NAND2X0 U6575 ( .IN1(n4637), .IN2(n4638), .QN(n4636) );
  NAND2X0 U6576 ( .IN1(n9050), .IN2(n7344), .QN(n4638) );
  NAND2X0 U6577 ( .IN1(n9090), .IN2(n7345), .QN(n4637) );
  NAND2X0 U6578 ( .IN1(n4639), .IN2(n4640), .QN(n4635) );
  NAND2X0 U6579 ( .IN1(n8922), .IN2(n4480), .QN(n4640) );
  NAND2X0 U6580 ( .IN1(n7347), .IN2(P1_N385), .QN(n4639) );
  NAND2X0 U6581 ( .IN1(n4641), .IN2(n4642), .QN(P1_N4646) );
  NAND2X0 U6582 ( .IN1(P1_N4578), .IN2(n4584), .QN(n4642) );
  NAND2X0 U6583 ( .IN1(P1_N5571), .IN2(n7096), .QN(n4641) );
  OR2X1 U6584 ( .IN2(n4644), .IN1(n4643), .Q(P1_N5169) );
  NAND2X0 U6585 ( .IN1(n4645), .IN2(n4646), .QN(n4644) );
  NAND2X0 U6586 ( .IN1(n9054), .IN2(n7344), .QN(n4646) );
  NAND2X0 U6587 ( .IN1(n9094), .IN2(n7345), .QN(n4645) );
  NAND2X0 U6588 ( .IN1(n4647), .IN2(n4648), .QN(n4643) );
  NAND2X0 U6589 ( .IN1(n8926), .IN2(n4480), .QN(n4648) );
  NAND2X0 U6590 ( .IN1(n7347), .IN2(P1_N384), .QN(n4647) );
  NAND2X0 U6591 ( .IN1(n4649), .IN2(n4650), .QN(P1_N4645) );
  NAND2X0 U6592 ( .IN1(P1_N4577), .IN2(n4584), .QN(n4650) );
  NAND2X0 U6593 ( .IN1(P1_N5571), .IN2(n7099), .QN(n4649) );
  OR2X1 U6594 ( .IN2(n4652), .IN1(n4651), .Q(P1_N5168) );
  NAND2X0 U6595 ( .IN1(n4653), .IN2(n4654), .QN(n4652) );
  NAND2X0 U6596 ( .IN1(n9493), .IN2(n7344), .QN(n4654) );
  NAND2X0 U6597 ( .IN1(n9497), .IN2(n7345), .QN(n4653) );
  NAND2X0 U6598 ( .IN1(n4655), .IN2(n4656), .QN(n4651) );
  NAND2X0 U6599 ( .IN1(n8930), .IN2(n4480), .QN(n4656) );
  NAND2X0 U6600 ( .IN1(n7347), .IN2(P1_N383), .QN(n4655) );
  NAND2X0 U6601 ( .IN1(n4657), .IN2(n4658), .QN(P1_N4644) );
  NAND2X0 U6602 ( .IN1(P1_N4576), .IN2(n4584), .QN(n4658) );
  NAND2X0 U6603 ( .IN1(P1_N5571), .IN2(n7103), .QN(n4657) );
  OR2X1 U6604 ( .IN2(n4660), .IN1(n4659), .Q(P1_N5167) );
  NAND2X0 U6605 ( .IN1(n4661), .IN2(n4662), .QN(n4660) );
  NAND2X0 U6606 ( .IN1(n9693), .IN2(n7344), .QN(n4662) );
  NAND2X0 U6607 ( .IN1(n9765), .IN2(n7345), .QN(n4661) );
  NAND2X0 U6608 ( .IN1(n4663), .IN2(n4664), .QN(n4659) );
  NAND2X0 U6609 ( .IN1(n8934), .IN2(n4480), .QN(n4664) );
  NAND2X0 U6610 ( .IN1(n7347), .IN2(P1_N382), .QN(n4663) );
  NAND2X0 U6611 ( .IN1(n4665), .IN2(n4666), .QN(P1_N4643) );
  NAND2X0 U6612 ( .IN1(P1_N4575), .IN2(n4584), .QN(n4666) );
  NAND2X0 U6613 ( .IN1(P1_N5571), .IN2(n7106), .QN(n4665) );
  OR2X1 U6614 ( .IN2(n4668), .IN1(n4667), .Q(P1_N5166) );
  NAND2X0 U6615 ( .IN1(n4669), .IN2(n4670), .QN(n4668) );
  NAND2X0 U6616 ( .IN1(n9697), .IN2(n7344), .QN(n4670) );
  NAND2X0 U6617 ( .IN1(n9769), .IN2(n7345), .QN(n4669) );
  NAND2X0 U6618 ( .IN1(n4671), .IN2(n4672), .QN(n4667) );
  NAND2X0 U6619 ( .IN1(n8938), .IN2(n4480), .QN(n4672) );
  NAND2X0 U6620 ( .IN1(n7347), .IN2(P1_N381), .QN(n4671) );
  NAND2X0 U6621 ( .IN1(n4673), .IN2(n4674), .QN(P1_N4642) );
  NAND2X0 U6622 ( .IN1(P1_N4574), .IN2(n4584), .QN(n4674) );
  NAND2X0 U6623 ( .IN1(P1_N5571), .IN2(n7110), .QN(n4673) );
  OR2X1 U6624 ( .IN2(n4676), .IN1(n4675), .Q(P1_N5165) );
  NAND2X0 U6625 ( .IN1(n4677), .IN2(n4678), .QN(n4676) );
  NAND2X0 U6626 ( .IN1(n9701), .IN2(n7344), .QN(n4678) );
  NAND2X0 U6627 ( .IN1(n9773), .IN2(n7345), .QN(n4677) );
  NAND2X0 U6628 ( .IN1(n4679), .IN2(n4680), .QN(n4675) );
  NAND2X0 U6629 ( .IN1(n8942), .IN2(n4480), .QN(n4680) );
  NAND2X0 U6630 ( .IN1(n7347), .IN2(P1_N380), .QN(n4679) );
  NAND2X0 U6631 ( .IN1(n4681), .IN2(n4682), .QN(P1_N4641) );
  NAND2X0 U6632 ( .IN1(P1_N4573), .IN2(n4584), .QN(n4682) );
  NAND2X0 U6633 ( .IN1(P1_N5571), .IN2(n7113), .QN(n4681) );
  OR2X1 U6634 ( .IN2(n4684), .IN1(n4683), .Q(P1_N5164) );
  NAND2X0 U6635 ( .IN1(n4685), .IN2(n4686), .QN(n4684) );
  NAND2X0 U6636 ( .IN1(n9705), .IN2(n7344), .QN(n4686) );
  NAND2X0 U6637 ( .IN1(n9777), .IN2(n7345), .QN(n4685) );
  NAND2X0 U6638 ( .IN1(n4687), .IN2(n4688), .QN(n4683) );
  NAND2X0 U6639 ( .IN1(n8946), .IN2(n4480), .QN(n4688) );
  NAND2X0 U6640 ( .IN1(n7347), .IN2(P1_N379), .QN(n4687) );
  NAND2X0 U6641 ( .IN1(n4689), .IN2(n4690), .QN(P1_N4640) );
  NAND2X0 U6642 ( .IN1(P1_N4572), .IN2(n4584), .QN(n4690) );
  NAND2X0 U6643 ( .IN1(P1_N5571), .IN2(n7116), .QN(n4689) );
  OR2X1 U6644 ( .IN2(n4692), .IN1(n4691), .Q(P1_N5163) );
  NAND2X0 U6645 ( .IN1(n4693), .IN2(n4694), .QN(n4692) );
  NAND2X0 U6646 ( .IN1(n9709), .IN2(n7344), .QN(n4694) );
  NAND2X0 U6647 ( .IN1(n9781), .IN2(n7345), .QN(n4693) );
  NAND2X0 U6648 ( .IN1(n4695), .IN2(n4696), .QN(n4691) );
  NAND2X0 U6649 ( .IN1(n8950), .IN2(n4480), .QN(n4696) );
  NAND2X0 U6650 ( .IN1(n7347), .IN2(P1_N378), .QN(n4695) );
  NAND2X0 U6460 ( .IN1(n4510), .IN2(P1_N4633), .QN(n4551) );
  NAND2X0 U6461 ( .IN1(P1_N372), .IN2(P1_N5574), .QN(n4550) );
  NAND2X0 U6462 ( .IN1(n4552), .IN2(n4553), .QN(P1_N4794) );
  NAND2X0 U6463 ( .IN1(n4510), .IN2(P1_N4632), .QN(n4553) );
  NAND2X0 U6464 ( .IN1(P1_N371), .IN2(P1_N5574), .QN(n4552) );
  NAND2X0 U6465 ( .IN1(n4554), .IN2(n4555), .QN(P1_N4793) );
  NAND2X0 U6466 ( .IN1(n4510), .IN2(P1_N4631), .QN(n4555) );
  NAND2X0 U6467 ( .IN1(P1_N370), .IN2(P1_N5574), .QN(n4554) );
  NAND2X0 U6468 ( .IN1(n4556), .IN2(n4557), .QN(P1_N4792) );
  NAND2X0 U6469 ( .IN1(n4510), .IN2(P1_N4630), .QN(n4557) );
  NAND2X0 U6470 ( .IN1(P1_N369), .IN2(P1_N5574), .QN(n4556) );
  NAND2X0 U6471 ( .IN1(n4558), .IN2(n4559), .QN(P1_N4791) );
  NAND2X0 U6472 ( .IN1(n4510), .IN2(P1_N4629), .QN(n4559) );
  NAND2X0 U6473 ( .IN1(P1_N368), .IN2(P1_N5574), .QN(n4558) );
  NAND2X0 U6474 ( .IN1(n4560), .IN2(n4561), .QN(P1_N4790) );
  NAND2X0 U6475 ( .IN1(n4510), .IN2(P1_N4628), .QN(n4561) );
  NAND2X0 U6476 ( .IN1(n18451), .IN2(P1_N5574), .QN(n4560) );
  NAND2X0 U6477 ( .IN1(n4562), .IN2(n4563), .QN(P1_N4789) );
  NAND2X0 U6478 ( .IN1(n4510), .IN2(P1_N4627), .QN(n4563) );
  NAND2X0 U6479 ( .IN1(n6623), .IN2(P1_N5574), .QN(n4562) );
  NAND2X0 U6480 ( .IN1(n4564), .IN2(n4565), .QN(P1_N4788) );
  NAND2X0 U6481 ( .IN1(n4510), .IN2(P1_N4626), .QN(n4565) );
  NAND2X0 U6482 ( .IN1(n6622), .IN2(P1_N5574), .QN(n4564) );
  NAND2X0 U6483 ( .IN1(n4566), .IN2(n4567), .QN(P1_N4787) );
  NAND2X0 U6484 ( .IN1(P1_N4625), .IN2(n4510), .QN(n4567) );
  NAND2X0 U6487 ( .IN1(n6621), .IN2(P1_N5574), .QN(n4566) );
  NAND2X0 U6492 ( .IN1(n7400), .IN2(n4570), .QN(P1_N4754) );
  NAND2X0 U6493 ( .IN1(n7399), .IN2(n4571), .QN(P1_N4752) );
  NOR2X0 U6494 ( .QN(P1_N4816), .IN1(n4571), .IN2(n4570) );
  INVX0 U6495 ( .ZN(n4570), .INP(n7399) );
  INVX0 U6496 ( .ZN(n4571), .INP(n7400) );
  NAND2X0 U6497 ( .IN1(n4572), .IN2(n4573), .QN(P1_N4654) );
  NAND2X0 U6498 ( .IN1(P1_N4586), .IN2(n4574), .QN(n4573) );
  INVX0 U6499 ( .ZN(n4574), .INP(n4506) );
  NOR2X0 U6500 ( .QN(n4506), .IN1(P1_N583), .IN2(n4575) );
  AND2X1 U6501 ( .IN1(P1_N506), .IN2(n6996), .Q(n4575) );
  NAND2X0 U6502 ( .IN1(P1_N5571), .IN2(P1_N5177), .QN(n4572) );
  OR2X1 U6503 ( .IN2(n4577), .IN1(n4576), .Q(P1_N5177) );
  NAND2X0 U6504 ( .IN1(n4578), .IN2(n4579), .QN(n4577) );
  NAND2X0 U6505 ( .IN1(n9022), .IN2(n7344), .QN(n4579) );
  NAND2X0 U6506 ( .IN1(n9062), .IN2(n7345), .QN(n4578) );
  NAND2X0 U6507 ( .IN1(n4580), .IN2(n4581), .QN(n4576) );
  NAND2X0 U6508 ( .IN1(n8894), .IN2(n4480), .QN(n4581) );
  NAND2X0 U6509 ( .IN1(n7347), .IN2(P1_N392), .QN(n4580) );
  NAND2X0 U6510 ( .IN1(n4582), .IN2(n4583), .QN(P1_N4653) );
  NAND2X0 U6511 ( .IN1(P1_N4585), .IN2(n4584), .QN(n4583) );
  NAND2X0 U6512 ( .IN1(P1_N5571), .IN2(n7122), .QN(n4582) );
  OR2X1 U6513 ( .IN2(n4586), .IN1(n4585), .Q(P1_N5176) );
  NAND2X0 U6514 ( .IN1(n4587), .IN2(n4588), .QN(n4586) );
  NAND2X0 U6515 ( .IN1(n9026), .IN2(n7344), .QN(n4588) );
  NAND2X0 U6516 ( .IN1(n9066), .IN2(n7345), .QN(n4587) );
  NAND2X0 U6517 ( .IN1(n4589), .IN2(n4590), .QN(n4585) );
  NAND2X0 U6518 ( .IN1(n8898), .IN2(n4480), .QN(n4590) );
  NAND2X0 U6519 ( .IN1(n7347), .IN2(P1_N391), .QN(n4589) );
  NAND2X0 U6520 ( .IN1(n4591), .IN2(n4592), .QN(P1_N4652) );
  NAND2X0 U6521 ( .IN1(P1_N4584), .IN2(n4584), .QN(n4592) );
  NAND2X0 U6522 ( .IN1(P1_N5571), .IN2(n7124), .QN(n4591) );
  OR2X1 U6523 ( .IN2(n4594), .IN1(n4593), .Q(P1_N5175) );
  NAND2X0 U6524 ( .IN1(n4595), .IN2(n4596), .QN(n4594) );
  NAND2X0 U6525 ( .IN1(n9030), .IN2(n7344), .QN(n4596) );
  NAND2X0 U6526 ( .IN1(n9070), .IN2(n7345), .QN(n4595) );
  NAND2X0 U6527 ( .IN1(n4597), .IN2(n4598), .QN(n4593) );
  NAND2X0 U6528 ( .IN1(n8902), .IN2(n4480), .QN(n4598) );
  NAND2X0 U6529 ( .IN1(n7347), .IN2(P1_N390), .QN(n4597) );
  NAND2X0 U6530 ( .IN1(n4599), .IN2(n4600), .QN(P1_N4651) );
  NAND2X0 U6531 ( .IN1(P1_N4583), .IN2(n4584), .QN(n4600) );
  NAND2X0 U6532 ( .IN1(P1_N5571), .IN2(P1_N5174), .QN(n4599) );
  OR2X1 U6533 ( .IN2(n4602), .IN1(n4601), .Q(P1_N5174) );
  NAND2X0 U6534 ( .IN1(n4603), .IN2(n4604), .QN(n4602) );
  NAND2X0 U6535 ( .IN1(n9034), .IN2(n7344), .QN(n4604) );
  NAND2X0 U6536 ( .IN1(n9074), .IN2(n7345), .QN(n4603) );
  NAND2X0 U6537 ( .IN1(n4605), .IN2(n4606), .QN(n4601) );
  NAND2X0 U6538 ( .IN1(n8906), .IN2(n4480), .QN(n4606) );
  NAND2X0 U6539 ( .IN1(n7347), .IN2(P1_N389), .QN(n4605) );
  NAND2X0 U6540 ( .IN1(n4607), .IN2(n4608), .QN(P1_N4650) );
  NAND2X0 U6541 ( .IN1(P1_N4582), .IN2(n4584), .QN(n4608) );
  NAND2X0 U6542 ( .IN1(P1_N5571), .IN2(n7138), .QN(n4607) );
  OR2X1 U6543 ( .IN2(n4610), .IN1(n4609), .Q(P1_N5173) );
  NAND2X0 U6544 ( .IN1(n4611), .IN2(n4612), .QN(n4610) );
  NAND2X0 U6545 ( .IN1(n9038), .IN2(n7344), .QN(n4612) );
  NAND2X0 U6546 ( .IN1(n9078), .IN2(n7345), .QN(n4611) );
  NAND2X0 U6547 ( .IN1(n4613), .IN2(n4614), .QN(n4609) );
  NAND2X0 U6548 ( .IN1(n8910), .IN2(n4480), .QN(n4614) );
  NAND2X0 U6549 ( .IN1(n7347), .IN2(P1_N388), .QN(n4613) );
  NAND2X0 U6551 ( .IN1(n4617), .IN2(n4618), .QN(P1_N4649) );
  NAND2X0 U6552 ( .IN1(P1_N4581), .IN2(n4584), .QN(n4618) );
  NAND2X0 U6553 ( .IN1(P1_N5571), .IN2(n7141), .QN(n4617) );
  OR2X1 U6554 ( .IN2(n4620), .IN1(n4619), .Q(P1_N5172) );
  NAND2X0 U6555 ( .IN1(n4621), .IN2(n4622), .QN(n4620) );
  NAND2X0 U6556 ( .IN1(n9042), .IN2(n7344), .QN(n4622) );
  NAND2X0 U6557 ( .IN1(n9082), .IN2(n7345), .QN(n4621) );
  NAND2X0 U6362 ( .IN1(n4483), .IN2(n4484), .QN(n4482) );
  NAND2X0 U6363 ( .IN1(n9018), .IN2(n7344), .QN(n4484) );
  NAND2X0 U6364 ( .IN1(n9058), .IN2(n7345), .QN(n4483) );
  NAND2X0 U6365 ( .IN1(n4485), .IN2(n4486), .QN(n4481) );
  NAND2X0 U6366 ( .IN1(n8890), .IN2(n4480), .QN(n4486) );
  NAND2X0 U6367 ( .IN1(P1_N393), .IN2(n7347), .QN(n4485) );
  NAND2X0 U6374 ( .IN1(P1_N815), .IN2(P1_N543), .QN(n4491) );
  NOR2X0 U6375 ( .QN(n4490), .IN1(n4492), .IN2(n4493) );
  NOR2X0 U6376 ( .QN(n4493), .IN1(n4084), .IN2(n4494) );
  INVX0 U6377 ( .ZN(n4084), .INP(n4175) );
  NAND2X0 U6378 ( .IN1(n4495), .IN2(n4496), .QN(n4175) );
  NAND2X0 U6379 ( .IN1(N38), .IN2(N5), .QN(n4496) );
  NAND2X0 U6380 ( .IN1(n9341), .IN2(n6739), .QN(n4495) );
  AND2X1 U6381 ( .IN1(n4497), .IN2(P1_N4588), .Q(n4492) );
  NAND2X0 U6383 ( .IN1(P1_N814), .IN2(P1_N543), .QN(n4499) );
  AND2X1 U6384 ( .IN1(P1_N542), .IN2(P1_N541), .Q(P1_N543) );
  NOR2X0 U6385 ( .QN(n4498), .IN1(n4500), .IN2(n4501) );
  NOR2X0 U6386 ( .QN(n4501), .IN1(n4086), .IN2(n4494) );
  AND2X1 U6387 ( .IN1(n4502), .IN2(n4503), .Q(n4494) );
  NAND2X0 U6388 ( .IN1(n7416), .IN2(n7019), .QN(n4503) );
  NAND2X0 U6389 ( .IN1(n7417), .IN2(n7019), .QN(n4502) );
  INVX0 U6390 ( .ZN(n4086), .INP(n4178) );
  NAND2X0 U6391 ( .IN1(n4504), .IN2(n4505), .QN(n4178) );
  NAND2X0 U6392 ( .IN1(N37), .IN2(N5), .QN(n4505) );
  NAND2X0 U6393 ( .IN1(n10107), .IN2(n6739), .QN(n4504) );
  AND2X1 U6394 ( .IN1(n4497), .IN2(P1_N4587), .Q(n4500) );
  NOR2X0 U6395 ( .QN(n4497), .IN1(n4506), .IN2(n7419) );
  NAND2X0 U6399 ( .IN1(n4508), .IN2(n4509), .QN(P1_N4815) );
  NAND2X0 U6400 ( .IN1(n4510), .IN2(P1_N4653), .QN(n4509) );
  NAND2X0 U6401 ( .IN1(P1_N392), .IN2(P1_N5574), .QN(n4508) );
  NAND2X0 U6402 ( .IN1(n4512), .IN2(n4513), .QN(P1_N4814) );
  NAND2X0 U6403 ( .IN1(n4510), .IN2(P1_N4652), .QN(n4513) );
  NAND2X0 U6404 ( .IN1(P1_N391), .IN2(P1_N5574), .QN(n4512) );
  NAND2X0 U6405 ( .IN1(n4514), .IN2(n4515), .QN(P1_N4813) );
  NAND2X0 U6406 ( .IN1(n4510), .IN2(P1_N4651), .QN(n4515) );
  NAND2X0 U6407 ( .IN1(P1_N390), .IN2(P1_N5574), .QN(n4514) );
  NAND2X0 U6408 ( .IN1(n4516), .IN2(n4517), .QN(P1_N4812) );
  NAND2X0 U6409 ( .IN1(n4510), .IN2(P1_N4650), .QN(n4517) );
  NAND2X0 U6410 ( .IN1(P1_N389), .IN2(P1_N5574), .QN(n4516) );
  NAND2X0 U6411 ( .IN1(n4518), .IN2(n4519), .QN(P1_N4811) );
  NAND2X0 U6412 ( .IN1(n4510), .IN2(P1_N4649), .QN(n4519) );
  NAND2X0 U6413 ( .IN1(P1_N388), .IN2(P1_N5574), .QN(n4518) );
  NAND2X0 U6414 ( .IN1(n4520), .IN2(n4521), .QN(P1_N4810) );
  NAND2X0 U6415 ( .IN1(n4510), .IN2(P1_N4648), .QN(n4521) );
  NAND2X0 U6416 ( .IN1(P1_N387), .IN2(P1_N5574), .QN(n4520) );
  NAND2X0 U6417 ( .IN1(n4522), .IN2(n4523), .QN(P1_N4809) );
  NAND2X0 U6418 ( .IN1(n4510), .IN2(P1_N4647), .QN(n4523) );
  NAND2X0 U6419 ( .IN1(P1_N386), .IN2(P1_N5574), .QN(n4522) );
  NAND2X0 U6420 ( .IN1(n4524), .IN2(n4525), .QN(P1_N4808) );
  NAND2X0 U6421 ( .IN1(n4510), .IN2(P1_N4646), .QN(n4525) );
  NAND2X0 U6422 ( .IN1(P1_N385), .IN2(P1_N5574), .QN(n4524) );
  NAND2X0 U6423 ( .IN1(n4526), .IN2(n4527), .QN(P1_N4807) );
  NAND2X0 U6424 ( .IN1(n4510), .IN2(P1_N4645), .QN(n4527) );
  NAND2X0 U6425 ( .IN1(P1_N384), .IN2(P1_N5574), .QN(n4526) );
  NAND2X0 U6426 ( .IN1(n4528), .IN2(n4529), .QN(P1_N4806) );
  NAND2X0 U6427 ( .IN1(n4510), .IN2(P1_N4644), .QN(n4529) );
  NAND2X0 U6428 ( .IN1(P1_N383), .IN2(P1_N5574), .QN(n4528) );
  NAND2X0 U6429 ( .IN1(n4530), .IN2(n4531), .QN(P1_N4805) );
  NAND2X0 U6430 ( .IN1(n4510), .IN2(P1_N4643), .QN(n4531) );
  NAND2X0 U6431 ( .IN1(P1_N382), .IN2(P1_N5574), .QN(n4530) );
  NAND2X0 U6432 ( .IN1(n4532), .IN2(n4533), .QN(P1_N4804) );
  NAND2X0 U6433 ( .IN1(n4510), .IN2(P1_N4642), .QN(n4533) );
  NAND2X0 U6434 ( .IN1(P1_N381), .IN2(P1_N5574), .QN(n4532) );
  NAND2X0 U6435 ( .IN1(n4534), .IN2(n4535), .QN(P1_N4803) );
  NAND2X0 U6436 ( .IN1(n4510), .IN2(P1_N4641), .QN(n4535) );
  NAND2X0 U6437 ( .IN1(P1_N380), .IN2(P1_N5574), .QN(n4534) );
  NAND2X0 U6438 ( .IN1(n4536), .IN2(n4537), .QN(P1_N4802) );
  NAND2X0 U6439 ( .IN1(n4510), .IN2(P1_N4640), .QN(n4537) );
  NAND2X0 U6440 ( .IN1(P1_N379), .IN2(P1_N5574), .QN(n4536) );
  NAND2X0 U6441 ( .IN1(n4538), .IN2(n4539), .QN(P1_N4801) );
  NAND2X0 U6442 ( .IN1(n4510), .IN2(P1_N4639), .QN(n4539) );
  NAND2X0 U6443 ( .IN1(P1_N378), .IN2(P1_N5574), .QN(n4538) );
  NAND2X0 U6444 ( .IN1(n4540), .IN2(n4541), .QN(P1_N4800) );
  NAND2X0 U6445 ( .IN1(n4510), .IN2(P1_N4638), .QN(n4541) );
  NAND2X0 U6446 ( .IN1(P1_N377), .IN2(P1_N5574), .QN(n4540) );
  NAND2X0 U6447 ( .IN1(n4542), .IN2(n4543), .QN(P1_N4799) );
  NAND2X0 U6448 ( .IN1(n4510), .IN2(P1_N4637), .QN(n4543) );
  NAND2X0 U6449 ( .IN1(P1_N376), .IN2(P1_N5574), .QN(n4542) );
  NAND2X0 U6450 ( .IN1(n4544), .IN2(n4545), .QN(P1_N4798) );
  NAND2X0 U6451 ( .IN1(n4510), .IN2(P1_N4636), .QN(n4545) );
  NAND2X0 U6452 ( .IN1(P1_N375), .IN2(P1_N5574), .QN(n4544) );
  NAND2X0 U6453 ( .IN1(n4546), .IN2(n4547), .QN(P1_N4797) );
  NAND2X0 U6454 ( .IN1(n4510), .IN2(P1_N4635), .QN(n4547) );
  NAND2X0 U6455 ( .IN1(P1_N374), .IN2(P1_N5574), .QN(n4546) );
  NAND2X0 U6456 ( .IN1(n4548), .IN2(n4549), .QN(P1_N4796) );
  NAND2X0 U6457 ( .IN1(n4510), .IN2(P1_N4634), .QN(n4549) );
  NAND2X0 U6458 ( .IN1(P1_N373), .IN2(P1_N5574), .QN(n4548) );
  NAND2X0 U6459 ( .IN1(n4550), .IN2(n4551), .QN(P1_N4795) );
  NAND2X0 U6267 ( .IN1(P1_N5158), .IN2(P1_N5147), .QN(n4429) );
  NAND2X0 U6268 ( .IN1(n4431), .IN2(n4432), .QN(P1_N5407) );
  NAND2X0 U6269 ( .IN1(n7072), .IN2(n7281), .QN(n4432) );
  NAND2X0 U6270 ( .IN1(n7072), .IN2(P1_N5147), .QN(n4431) );
  NAND2X0 U6271 ( .IN1(n4433), .IN2(n4434), .QN(P1_N5406) );
  NAND2X0 U6272 ( .IN1(n7075), .IN2(n7281), .QN(n4434) );
  NAND2X0 U6273 ( .IN1(n7075), .IN2(P1_N5147), .QN(n4433) );
  NAND2X0 U6274 ( .IN1(n4435), .IN2(n4436), .QN(P1_N5405) );
  NAND2X0 U6275 ( .IN1(P1_N5155), .IN2(n7281), .QN(n4436) );
  NAND2X0 U6276 ( .IN1(P1_N5155), .IN2(P1_N5147), .QN(n4435) );
  NAND2X0 U6277 ( .IN1(n4437), .IN2(n4438), .QN(P1_N5404) );
  NAND2X0 U6278 ( .IN1(P1_N5154), .IN2(n7281), .QN(n4438) );
  NAND2X0 U6279 ( .IN1(P1_N5154), .IN2(P1_N5147), .QN(n4437) );
  NAND2X0 U6280 ( .IN1(n4439), .IN2(n4440), .QN(P1_N5403) );
  NAND2X0 U6281 ( .IN1(n7036), .IN2(n7281), .QN(n4440) );
  NAND2X0 U6282 ( .IN1(n7036), .IN2(P1_N5147), .QN(n4439) );
  NAND2X0 U6283 ( .IN1(n4441), .IN2(n4442), .QN(P1_N5402) );
  NAND2X0 U6284 ( .IN1(P1_N5152), .IN2(n7281), .QN(n4442) );
  NAND2X0 U6285 ( .IN1(P1_N5152), .IN2(P1_N5147), .QN(n4441) );
  NAND2X0 U6286 ( .IN1(n4443), .IN2(n4444), .QN(P1_N5401) );
  NAND2X0 U6287 ( .IN1(P1_N5151), .IN2(n7281), .QN(n4444) );
  NAND2X0 U6288 ( .IN1(P1_N5151), .IN2(P1_N5147), .QN(n4443) );
  NAND2X0 U6289 ( .IN1(n4445), .IN2(n4446), .QN(P1_N5400) );
  NAND2X0 U6290 ( .IN1(P1_N5150), .IN2(n7281), .QN(n4446) );
  NAND2X0 U6291 ( .IN1(P1_N5150), .IN2(P1_N5147), .QN(n4445) );
  NAND2X0 U6292 ( .IN1(n4447), .IN2(n4448), .QN(P1_N5399) );
  NAND2X0 U6293 ( .IN1(n7034), .IN2(n7281), .QN(n4448) );
  NAND2X0 U6295 ( .IN1(n7034), .IN2(P1_N5147), .QN(n4447) );
  NOR2X0 U6296 ( .QN(P1_N5115), .IN1(n4084), .IN2(n7027) );
  NOR2X0 U6297 ( .QN(P1_N5114), .IN1(n4086), .IN2(n7027) );
  NOR2X0 U6298 ( .QN(P1_N5113), .IN1(n7328), .IN2(n7029) );
  NOR2X0 U6299 ( .QN(P1_N5112), .IN1(n7326), .IN2(n7029) );
  NOR2X0 U6300 ( .QN(P1_N5111), .IN1(n7324), .IN2(n7029) );
  NOR2X0 U6301 ( .QN(P1_N5110), .IN1(n7322), .IN2(n7029) );
  NOR2X0 U6302 ( .QN(P1_N5109), .IN1(n7320), .IN2(n7027) );
  NOR2X0 U6303 ( .QN(P1_N5108), .IN1(n7318), .IN2(n7027) );
  NOR2X0 U6304 ( .QN(P1_N5107), .IN1(n7316), .IN2(n7027) );
  NOR2X0 U6305 ( .QN(P1_N5106), .IN1(n7314), .IN2(n7027) );
  NOR2X0 U6306 ( .QN(P1_N5105), .IN1(n7312), .IN2(n7027) );
  NOR2X0 U6307 ( .QN(P1_N5104), .IN1(n7310), .IN2(n7023) );
  NAND2X0 U6309 ( .IN1(n4097), .IN2(n4449), .QN(P1_N5103) );
  NAND2X0 U6310 ( .IN1(n7019), .IN2(n4099), .QN(n4449) );
  NAND2X0 U6311 ( .IN1(n4100), .IN2(n4450), .QN(P1_N5102) );
  NAND2X0 U6312 ( .IN1(n7028), .IN2(n4102), .QN(n4450) );
  NAND2X0 U6313 ( .IN1(n4103), .IN2(n4451), .QN(P1_N5101) );
  NAND2X0 U6314 ( .IN1(n7028), .IN2(n4105), .QN(n4451) );
  NAND2X0 U6315 ( .IN1(n4106), .IN2(n4452), .QN(P1_N5100) );
  NAND2X0 U6316 ( .IN1(n7028), .IN2(n4108), .QN(n4452) );
  NAND2X0 U6317 ( .IN1(n4109), .IN2(n4453), .QN(P1_N5099) );
  NAND2X0 U6318 ( .IN1(n7028), .IN2(n4111), .QN(n4453) );
  NAND2X0 U6319 ( .IN1(n4112), .IN2(n4454), .QN(P1_N5098) );
  NAND2X0 U6320 ( .IN1(n7024), .IN2(n4114), .QN(n4454) );
  NAND2X0 U6321 ( .IN1(n4115), .IN2(n4455), .QN(P1_N5097) );
  NAND2X0 U6322 ( .IN1(n7024), .IN2(n4117), .QN(n4455) );
  NAND2X0 U6323 ( .IN1(n4118), .IN2(n4456), .QN(P1_N5096) );
  NAND2X0 U6324 ( .IN1(n7024), .IN2(n4120), .QN(n4456) );
  NAND2X0 U6325 ( .IN1(n4121), .IN2(n4457), .QN(P1_N5095) );
  NAND2X0 U6326 ( .IN1(n7024), .IN2(n4123), .QN(n4457) );
  NAND2X0 U6327 ( .IN1(n4124), .IN2(n4458), .QN(P1_N5094) );
  NAND2X0 U6328 ( .IN1(n7024), .IN2(n4126), .QN(n4458) );
  NAND2X0 U6329 ( .IN1(n4127), .IN2(n4459), .QN(P1_N5093) );
  NAND2X0 U6330 ( .IN1(n7463), .IN2(n4129), .QN(n4459) );
  NAND2X0 U6331 ( .IN1(n4130), .IN2(n4460), .QN(P1_N5092) );
  NAND2X0 U6332 ( .IN1(n7463), .IN2(n4132), .QN(n4460) );
  NAND2X0 U6333 ( .IN1(n4133), .IN2(n4461), .QN(P1_N5091) );
  NAND2X0 U6334 ( .IN1(n7463), .IN2(n4135), .QN(n4461) );
  NAND2X0 U6335 ( .IN1(n4136), .IN2(n4462), .QN(P1_N5090) );
  NAND2X0 U6336 ( .IN1(n7463), .IN2(n4138), .QN(n4462) );
  NAND2X0 U6337 ( .IN1(n4139), .IN2(n4463), .QN(P1_N5089) );
  NAND2X0 U6338 ( .IN1(n7026), .IN2(n4141), .QN(n4463) );
  NAND2X0 U6339 ( .IN1(n4142), .IN2(n4464), .QN(P1_N5088) );
  NAND2X0 U6340 ( .IN1(n7026), .IN2(n4144), .QN(n4464) );
  NAND2X0 U6341 ( .IN1(n4145), .IN2(n4465), .QN(P1_N5087) );
  NAND2X0 U6342 ( .IN1(n7026), .IN2(n4147), .QN(n4465) );
  NAND2X0 U6343 ( .IN1(n4148), .IN2(n4466), .QN(P1_N5086) );
  NAND2X0 U6344 ( .IN1(n7022), .IN2(n4150), .QN(n4466) );
  NAND2X0 U6345 ( .IN1(n4151), .IN2(n4467), .QN(P1_N5085) );
  NAND2X0 U6346 ( .IN1(n7022), .IN2(n4153), .QN(n4467) );
  NAND2X0 U6347 ( .IN1(n4154), .IN2(n4468), .QN(P1_N5084) );
  NAND2X0 U6348 ( .IN1(n7022), .IN2(n4156), .QN(n4468) );
  NAND2X0 U6350 ( .IN1(n4470), .IN2(n4471), .QN(P1_N4977) );
  NAND2X0 U6351 ( .IN1(P1_N4971), .IN2(n7340), .QN(n4471) );
  AND2X1 U6352 ( .IN1(n4472), .IN2(n4473), .Q(n4470) );
  NAND2X0 U6353 ( .IN1(P1_N5570), .IN2(P1_N363), .QN(n4473) );
  NAND2X0 U6354 ( .IN1(P1_N4970), .IN2(n7337), .QN(n4472) );
  OR2X1 U6355 ( .IN2(n4475), .IN1(n7348), .Q(P1_N497) );
  NAND2X0 U6356 ( .IN1(n4476), .IN2(n4477), .QN(n4475) );
  NAND2X0 U6357 ( .IN1(n9014), .IN2(n7344), .QN(n4477) );
  NAND2X0 U6358 ( .IN1(n8882), .IN2(n7345), .QN(n4476) );
  OR2X1 U6361 ( .IN2(n4482), .IN1(n4481), .Q(P1_N5178) );
  AND2X1 U6170 ( .IN1(P1_N4818), .IN2(n4366), .Q(n4363) );
  NAND2X0 U6171 ( .IN1(n4359), .IN2(P1_N4969), .QN(n4360) );
  NOR2X0 U6172 ( .QN(n4359), .IN1(n7414), .IN2(n4367) );
  INVX0 U6181 ( .ZN(n4367), .INP(P1_N499) );
  NAND2X0 U6182 ( .IN1(n4370), .IN2(n4371), .QN(P1_N531) );
  NAND2X0 U6183 ( .IN1(n4370), .IN2(n4372), .QN(P1_N530) );
  NAND2X0 U6184 ( .IN1(P1_N517), .IN2(n4371), .QN(n4372) );
  INVX0 U6185 ( .ZN(n4371), .INP(P1_N514) );
  AND2X1 U6186 ( .IN1(n4373), .IN2(n4374), .Q(n4370) );
  NOR2X0 U6187 ( .QN(n4373), .IN1(P1_N511), .IN2(P1_N508) );
  NAND2X0 U6189 ( .IN1(n4377), .IN2(n4374), .QN(n4376) );
  INVX0 U6190 ( .ZN(n4374), .INP(P1_N504) );
  NAND2X0 U6191 ( .IN1(n4378), .IN2(n4379), .QN(n4377) );
  NAND2X0 U6192 ( .IN1(n4380), .IN2(n4381), .QN(n4379) );
  NAND2X0 U6193 ( .IN1(n4382), .IN2(n4383), .QN(n4380) );
  NOR2X0 U6194 ( .QN(n4383), .IN1(P1_N519), .IN2(P1_N517) );
  NOR2X0 U6195 ( .QN(n4382), .IN1(P1_N514), .IN2(P1_N511) );
  OR2X1 U6196 ( .IN2(P1_N506), .IN1(n4381), .Q(n4378) );
  INVX0 U6197 ( .ZN(n4381), .INP(P1_N508) );
  NAND2X0 U6198 ( .IN1(P1_N506), .IN2(P1_N504), .QN(n4375) );
  NAND2X0 U6199 ( .IN1(n4384), .IN2(n4385), .QN(P1_N5430) );
  NAND2X0 U6200 ( .IN1(n7052), .IN2(n7281), .QN(n4385) );
  NAND2X0 U6201 ( .IN1(P1_N5180), .IN2(P1_N5147), .QN(n4384) );
  NAND2X0 U6202 ( .IN1(n4387), .IN2(n4388), .QN(P1_N5429) );
  NAND2X0 U6203 ( .IN1(P1_N497), .IN2(n7281), .QN(n4388) );
  NAND2X0 U6204 ( .IN1(n7145), .IN2(P1_N5147), .QN(n4387) );
  NAND2X0 U6205 ( .IN1(n4389), .IN2(n4390), .QN(P1_N5428) );
  NAND2X0 U6206 ( .IN1(P1_N5178), .IN2(n7281), .QN(n4390) );
  NAND2X0 U6207 ( .IN1(P1_N5178), .IN2(P1_N5147), .QN(n4389) );
  NAND2X0 U6208 ( .IN1(n4391), .IN2(n4392), .QN(P1_N5427) );
  NAND2X0 U6209 ( .IN1(P1_N5177), .IN2(n7281), .QN(n4392) );
  NAND2X0 U6210 ( .IN1(P1_N5177), .IN2(P1_N5147), .QN(n4391) );
  NAND2X0 U6211 ( .IN1(n4393), .IN2(n4394), .QN(P1_N5426) );
  NAND2X0 U6212 ( .IN1(P1_N5176), .IN2(n7281), .QN(n4394) );
  NAND2X0 U6213 ( .IN1(P1_N5176), .IN2(P1_N5147), .QN(n4393) );
  NAND2X0 U6214 ( .IN1(n4395), .IN2(n4396), .QN(P1_N5425) );
  NAND2X0 U6215 ( .IN1(P1_N5175), .IN2(n7281), .QN(n4396) );
  NAND2X0 U6216 ( .IN1(P1_N5175), .IN2(P1_N5147), .QN(n4395) );
  NAND2X0 U6217 ( .IN1(n4397), .IN2(n4398), .QN(P1_N5424) );
  NAND2X0 U6218 ( .IN1(P1_N5174), .IN2(n7281), .QN(n4398) );
  NAND2X0 U6219 ( .IN1(P1_N5174), .IN2(P1_N5147), .QN(n4397) );
  NAND2X0 U6220 ( .IN1(n4399), .IN2(n4400), .QN(P1_N5423) );
  NAND2X0 U6221 ( .IN1(P1_N5173), .IN2(n7281), .QN(n4400) );
  NAND2X0 U6222 ( .IN1(P1_N5173), .IN2(P1_N5147), .QN(n4399) );
  NAND2X0 U6223 ( .IN1(n4401), .IN2(n4402), .QN(P1_N5422) );
  NAND2X0 U6224 ( .IN1(n7141), .IN2(n7281), .QN(n4402) );
  NAND2X0 U6225 ( .IN1(n7141), .IN2(P1_N5147), .QN(n4401) );
  NAND2X0 U6226 ( .IN1(n4403), .IN2(n4404), .QN(P1_N5421) );
  NAND2X0 U6227 ( .IN1(P1_N5171), .IN2(n7281), .QN(n4404) );
  NAND2X0 U6228 ( .IN1(n7089), .IN2(P1_N5147), .QN(n4403) );
  NAND2X0 U6229 ( .IN1(n4405), .IN2(n4406), .QN(P1_N5420) );
  NAND2X0 U6230 ( .IN1(P1_N5170), .IN2(n7281), .QN(n4406) );
  NAND2X0 U6231 ( .IN1(P1_N5170), .IN2(P1_N5147), .QN(n4405) );
  NAND2X0 U6232 ( .IN1(n4407), .IN2(n4408), .QN(P1_N5419) );
  NAND2X0 U6233 ( .IN1(P1_N5169), .IN2(n7281), .QN(n4408) );
  NAND2X0 U6234 ( .IN1(P1_N5169), .IN2(P1_N5147), .QN(n4407) );
  NAND2X0 U6235 ( .IN1(n4409), .IN2(n4410), .QN(P1_N5418) );
  NAND2X0 U6236 ( .IN1(n7099), .IN2(n7281), .QN(n4410) );
  NAND2X0 U6237 ( .IN1(n7099), .IN2(P1_N5147), .QN(n4409) );
  NAND2X0 U6238 ( .IN1(n4411), .IN2(n4412), .QN(P1_N5417) );
  NAND2X0 U6239 ( .IN1(P1_N5167), .IN2(n7281), .QN(n4412) );
  NAND2X0 U6240 ( .IN1(P1_N5167), .IN2(P1_N5147), .QN(n4411) );
  NAND2X0 U6241 ( .IN1(n4413), .IN2(n4414), .QN(P1_N5416) );
  NAND2X0 U6242 ( .IN1(P1_N5166), .IN2(n7281), .QN(n4414) );
  NAND2X0 U6243 ( .IN1(n7106), .IN2(P1_N5147), .QN(n4413) );
  NAND2X0 U6244 ( .IN1(n4415), .IN2(n4416), .QN(P1_N5415) );
  NAND2X0 U6245 ( .IN1(P1_N5165), .IN2(n7281), .QN(n4416) );
  NAND2X0 U6246 ( .IN1(n7110), .IN2(P1_N5147), .QN(n4415) );
  NAND2X0 U6247 ( .IN1(n4417), .IN2(n4418), .QN(P1_N5414) );
  NAND2X0 U6248 ( .IN1(P1_N5164), .IN2(n7281), .QN(n4418) );
  NAND2X0 U6249 ( .IN1(P1_N5164), .IN2(P1_N5147), .QN(n4417) );
  NAND2X0 U6250 ( .IN1(n4419), .IN2(n4420), .QN(P1_N5413) );
  NAND2X0 U6251 ( .IN1(P1_N5163), .IN2(n7281), .QN(n4420) );
  NAND2X0 U6252 ( .IN1(P1_N5163), .IN2(P1_N5147), .QN(n4419) );
  NAND2X0 U6253 ( .IN1(n4421), .IN2(n4422), .QN(P1_N5412) );
  NAND2X0 U6254 ( .IN1(P1_N5162), .IN2(n7281), .QN(n4422) );
  NAND2X0 U6255 ( .IN1(P1_N5162), .IN2(P1_N5147), .QN(n4421) );
  NAND2X0 U6256 ( .IN1(n4423), .IN2(n4424), .QN(P1_N5411) );
  NAND2X0 U6257 ( .IN1(P1_N5161), .IN2(n7281), .QN(n4424) );
  NAND2X0 U6258 ( .IN1(P1_N5161), .IN2(P1_N5147), .QN(n4423) );
  NAND2X0 U6259 ( .IN1(n4425), .IN2(n4426), .QN(P1_N5410) );
  NAND2X0 U6260 ( .IN1(P1_N5160), .IN2(n7281), .QN(n4426) );
  NAND2X0 U6261 ( .IN1(P1_N5160), .IN2(P1_N5147), .QN(n4425) );
  NAND2X0 U6262 ( .IN1(n4427), .IN2(n4428), .QN(P1_N5409) );
  NAND2X0 U6263 ( .IN1(P1_N5159), .IN2(n7281), .QN(n4428) );
  NAND2X0 U6264 ( .IN1(P1_N5159), .IN2(P1_N5147), .QN(n4427) );
  NAND2X0 U6265 ( .IN1(n4429), .IN2(n4430), .QN(P1_N5408) );
  NAND2X0 U6266 ( .IN1(P1_N5158), .IN2(n7281), .QN(n4430) );
  OR2X1 U6058 ( .IN2(n4272), .IN1(n7428), .Q(P1_N5513) );
  NAND2X0 U6059 ( .IN1(n4273), .IN2(n4274), .QN(n4272) );
  NAND2X0 U6060 ( .IN1(P1_N4834), .IN2(n4164), .QN(n4274) );
  NAND2X0 U6061 ( .IN1(n9669), .IN2(n6583), .QN(n4273) );
  OR2X1 U6064 ( .IN2(n4277), .IN1(n7429), .Q(P1_N5512) );
  NAND2X0 U6065 ( .IN1(n4278), .IN2(n4279), .QN(n4277) );
  NAND2X0 U6066 ( .IN1(P1_N4833), .IN2(n4164), .QN(n4279) );
  NAND2X0 U6067 ( .IN1(n9859), .IN2(n6583), .QN(n4278) );
  OR2X1 U6070 ( .IN2(n4282), .IN1(n7430), .Q(P1_N5511) );
  NAND2X0 U6071 ( .IN1(n4283), .IN2(n4284), .QN(n4282) );
  NAND2X0 U6072 ( .IN1(P1_N4832), .IN2(n4164), .QN(n4284) );
  NAND2X0 U6073 ( .IN1(n9673), .IN2(n6583), .QN(n4283) );
  OR2X1 U6076 ( .IN2(n4287), .IN1(n7431), .Q(P1_N5510) );
  NAND2X0 U6077 ( .IN1(n4288), .IN2(n4289), .QN(n4287) );
  NAND2X0 U6078 ( .IN1(P1_N4831), .IN2(n4164), .QN(n4289) );
  NAND2X0 U6079 ( .IN1(n9863), .IN2(n6583), .QN(n4288) );
  OR2X1 U6082 ( .IN2(n4292), .IN1(n7432), .Q(P1_N5509) );
  NAND2X0 U6083 ( .IN1(n4293), .IN2(n4294), .QN(n4292) );
  NAND2X0 U6084 ( .IN1(P1_N4830), .IN2(n4164), .QN(n4294) );
  NAND2X0 U6085 ( .IN1(n9677), .IN2(n6583), .QN(n4293) );
  OR2X1 U6088 ( .IN2(n4297), .IN1(n7433), .Q(P1_N5508) );
  NAND2X0 U6089 ( .IN1(n4298), .IN2(n4299), .QN(n4297) );
  NAND2X0 U6090 ( .IN1(P1_N4829), .IN2(n4164), .QN(n4299) );
  NAND2X0 U6091 ( .IN1(n9867), .IN2(n6583), .QN(n4298) );
  OR2X1 U6094 ( .IN2(n4302), .IN1(n7434), .Q(P1_N5507) );
  NAND2X0 U6095 ( .IN1(n4303), .IN2(n4304), .QN(n4302) );
  NAND2X0 U6096 ( .IN1(P1_N4828), .IN2(n4164), .QN(n4304) );
  NAND2X0 U6097 ( .IN1(n9681), .IN2(n6583), .QN(n4303) );
  OR2X1 U6100 ( .IN2(n4307), .IN1(n7435), .Q(P1_N5506) );
  NAND2X0 U6101 ( .IN1(n4308), .IN2(n4309), .QN(n4307) );
  NAND2X0 U6102 ( .IN1(P1_N4827), .IN2(n4164), .QN(n4309) );
  NAND2X0 U6103 ( .IN1(n10011), .IN2(n6583), .QN(n4308) );
  OR2X1 U6106 ( .IN2(n4312), .IN1(n7436), .Q(P1_N5505) );
  NAND2X0 U6107 ( .IN1(n4313), .IN2(n4314), .QN(n4312) );
  NAND2X0 U6108 ( .IN1(P1_N4826), .IN2(n4164), .QN(n4314) );
  NAND2X0 U6109 ( .IN1(n9685), .IN2(n6583), .QN(n4313) );
  OR2X1 U6113 ( .IN2(n4317), .IN1(n7437), .Q(P1_N5504) );
  NAND2X0 U6114 ( .IN1(n4318), .IN2(n4319), .QN(n4317) );
  NAND2X0 U6115 ( .IN1(P1_N4825), .IN2(n4164), .QN(n4319) );
  NAND2X0 U6116 ( .IN1(n10015), .IN2(n6580), .QN(n4318) );
  OR2X1 U6120 ( .IN2(n4323), .IN1(n7438), .Q(P1_N5503) );
  NAND2X0 U6121 ( .IN1(n4324), .IN2(n4325), .QN(n4323) );
  NAND2X0 U6122 ( .IN1(P1_N4824), .IN2(n4164), .QN(n4325) );
  NAND2X0 U6123 ( .IN1(n9689), .IN2(n6580), .QN(n4324) );
  OR2X1 U6127 ( .IN2(n4329), .IN1(n4328), .Q(P1_N5502) );
  NAND2X0 U6128 ( .IN1(n4330), .IN2(n4331), .QN(n4329) );
  NAND2X0 U6129 ( .IN1(P1_N4823), .IN2(n4164), .QN(n4331) );
  NAND2X0 U6130 ( .IN1(n9657), .IN2(n6580), .QN(n4330) );
  NAND2X0 U6131 ( .IN1(n4332), .IN2(n4333), .QN(n4328) );
  NAND2X0 U6132 ( .IN1(P1_N4977), .IN2(n4172), .QN(n4333) );
  NAND2X0 U6133 ( .IN1(n4171), .IN2(P1_N667), .QN(n4332) );
  OR2X1 U6134 ( .IN2(n4335), .IN1(n7439), .Q(P1_N5501) );
  NAND2X0 U6135 ( .IN1(n4336), .IN2(n4337), .QN(n4335) );
  NAND2X0 U6136 ( .IN1(P1_N4822), .IN2(n4164), .QN(n4337) );
  NAND2X0 U6137 ( .IN1(n6594), .IN2(n6580), .QN(n4336) );
  OR2X1 U6141 ( .IN2(n4341), .IN1(n4340), .Q(P1_N5500) );
  NAND2X0 U6142 ( .IN1(n4342), .IN2(n4343), .QN(n4341) );
  NAND2X0 U6143 ( .IN1(P1_N4821), .IN2(n4164), .QN(n4343) );
  NAND2X0 U6144 ( .IN1(n6623), .IN2(n6580), .QN(n4342) );
  NAND2X0 U6145 ( .IN1(n4344), .IN2(n4345), .QN(n4340) );
  NAND2X0 U6146 ( .IN1(P1_N4977), .IN2(n4172), .QN(n4345) );
  NAND2X0 U6147 ( .IN1(n4171), .IN2(P1_N665), .QN(n4344) );
  OR2X1 U6148 ( .IN2(n4347), .IN1(n7440), .Q(P1_N5499) );
  NAND2X0 U6149 ( .IN1(n4348), .IN2(n4349), .QN(n4347) );
  NAND2X0 U6150 ( .IN1(P1_N4820), .IN2(n4164), .QN(n4349) );
  NAND2X0 U6151 ( .IN1(n6622), .IN2(n6580), .QN(n4348) );
  OR2X1 U6155 ( .IN2(n4353), .IN1(n7441), .Q(P1_N5498) );
  NAND2X0 U6156 ( .IN1(n4354), .IN2(n4355), .QN(n4353) );
  NAND2X0 U6157 ( .IN1(P1_N4819), .IN2(n4164), .QN(n4355) );
  NAND2X0 U6159 ( .IN1(n6621), .IN2(n6580), .QN(n4354) );
  AND2X1 U6162 ( .IN1(n4359), .IN2(n6584), .Q(n4172) );
  NAND2X0 U6165 ( .IN1(n4360), .IN2(n4361), .QN(P1_N5497) );
  INVX0 U6166 ( .ZN(n4361), .INP(P1_N5518) );
  NAND2X0 U6167 ( .IN1(n4362), .IN2(n6584), .QN(P1_N5518) );
  NOR2X0 U6168 ( .QN(n4362), .IN1(n4363), .IN2(n4364) );
  NOR2X0 U6169 ( .QN(n4364), .IN1(P1_N499), .IN2(n7023) );
  NAND2X0 U5960 ( .IN1(n4199), .IN2(n6580), .QN(n4198) );
  NAND2X0 U5961 ( .IN1(P1_N125), .IN2(n6584), .QN(n4197) );
  NAND2X0 U5962 ( .IN1(n4200), .IN2(n4201), .QN(P1_N5543) );
  NAND2X0 U5963 ( .IN1(n4202), .IN2(n6580), .QN(n4201) );
  NAND2X0 U5964 ( .IN1(P1_N124), .IN2(n6584), .QN(n4200) );
  NAND2X0 U5965 ( .IN1(n4203), .IN2(n4204), .QN(P1_N5542) );
  NAND2X0 U5966 ( .IN1(n4205), .IN2(n6583), .QN(n4204) );
  NAND2X0 U5967 ( .IN1(P1_N123), .IN2(n6582), .QN(n4203) );
  NAND2X0 U5968 ( .IN1(n4206), .IN2(n4207), .QN(P1_N5541) );
  NAND2X0 U5969 ( .IN1(n4208), .IN2(n6583), .QN(n4207) );
  NAND2X0 U5970 ( .IN1(P1_N122), .IN2(n6582), .QN(n4206) );
  NAND2X0 U5971 ( .IN1(n4209), .IN2(n4210), .QN(P1_N5540) );
  NAND2X0 U5972 ( .IN1(n4099), .IN2(n4169), .QN(n4210) );
  NAND2X0 U5973 ( .IN1(P1_N121), .IN2(n6582), .QN(n4209) );
  NAND2X0 U5974 ( .IN1(n4211), .IN2(n4212), .QN(P1_N5539) );
  NAND2X0 U5975 ( .IN1(n4102), .IN2(n4169), .QN(n4212) );
  NAND2X0 U5976 ( .IN1(P1_N120), .IN2(n6582), .QN(n4211) );
  NAND2X0 U5977 ( .IN1(n4213), .IN2(n4214), .QN(P1_N5538) );
  NAND2X0 U5978 ( .IN1(n4105), .IN2(n4169), .QN(n4214) );
  NAND2X0 U5979 ( .IN1(P1_N119), .IN2(n6582), .QN(n4213) );
  NAND2X0 U5980 ( .IN1(n4215), .IN2(n4216), .QN(P1_N5537) );
  NAND2X0 U5981 ( .IN1(n4108), .IN2(n4169), .QN(n4216) );
  NAND2X0 U5982 ( .IN1(P1_N118), .IN2(n6582), .QN(n4215) );
  NAND2X0 U5983 ( .IN1(n4217), .IN2(n4218), .QN(P1_N5536) );
  NAND2X0 U5984 ( .IN1(n4111), .IN2(n4169), .QN(n4218) );
  NAND2X0 U5985 ( .IN1(P1_N117), .IN2(n6582), .QN(n4217) );
  NAND2X0 U5986 ( .IN1(n4219), .IN2(n4220), .QN(P1_N5535) );
  NAND2X0 U5987 ( .IN1(n4114), .IN2(n4169), .QN(n4220) );
  NAND2X0 U5988 ( .IN1(P1_N116), .IN2(n6582), .QN(n4219) );
  NAND2X0 U5989 ( .IN1(n4221), .IN2(n4222), .QN(P1_N5534) );
  NAND2X0 U5990 ( .IN1(n4117), .IN2(n4169), .QN(n4222) );
  NAND2X0 U5991 ( .IN1(P1_N115), .IN2(n6582), .QN(n4221) );
  NAND2X0 U5992 ( .IN1(n4223), .IN2(n4224), .QN(P1_N5532) );
  NAND2X0 U5993 ( .IN1(n4120), .IN2(n4169), .QN(n4224) );
  NAND2X0 U5994 ( .IN1(P1_N114), .IN2(n6582), .QN(n4223) );
  NAND2X0 U5995 ( .IN1(n4225), .IN2(n4226), .QN(P1_N5531) );
  NAND2X0 U5996 ( .IN1(n4123), .IN2(n4169), .QN(n4226) );
  NAND2X0 U5997 ( .IN1(P1_N113), .IN2(n6582), .QN(n4225) );
  NAND2X0 U5998 ( .IN1(n4227), .IN2(n4228), .QN(P1_N5530) );
  NAND2X0 U5999 ( .IN1(n4126), .IN2(n4169), .QN(n4228) );
  NAND2X0 U6000 ( .IN1(P1_N112), .IN2(n6582), .QN(n4227) );
  NAND2X0 U6001 ( .IN1(n4229), .IN2(n4230), .QN(P1_N5529) );
  NAND2X0 U6002 ( .IN1(n4129), .IN2(n4169), .QN(n4230) );
  NAND2X0 U6003 ( .IN1(P1_N111), .IN2(n6582), .QN(n4229) );
  NAND2X0 U6004 ( .IN1(n4231), .IN2(n4232), .QN(P1_N5528) );
  NAND2X0 U6005 ( .IN1(n4132), .IN2(n4169), .QN(n4232) );
  NAND2X0 U6006 ( .IN1(P1_N110), .IN2(n6582), .QN(n4231) );
  NAND2X0 U6007 ( .IN1(n4233), .IN2(n4234), .QN(P1_N5527) );
  NAND2X0 U6008 ( .IN1(n4135), .IN2(n4169), .QN(n4234) );
  NAND2X0 U6009 ( .IN1(P1_N109), .IN2(n6582), .QN(n4233) );
  NAND2X0 U6010 ( .IN1(n4235), .IN2(n4236), .QN(P1_N5526) );
  NAND2X0 U6011 ( .IN1(n4138), .IN2(n4169), .QN(n4236) );
  NAND2X0 U6012 ( .IN1(P1_N108), .IN2(n6582), .QN(n4235) );
  NAND2X0 U6013 ( .IN1(n4237), .IN2(n4238), .QN(P1_N5525) );
  NAND2X0 U6014 ( .IN1(n4141), .IN2(n4169), .QN(n4238) );
  NAND2X0 U6015 ( .IN1(P1_N107), .IN2(n6582), .QN(n4237) );
  NAND2X0 U6016 ( .IN1(n4239), .IN2(n4240), .QN(P1_N5524) );
  NAND2X0 U6017 ( .IN1(n4144), .IN2(n4169), .QN(n4240) );
  NAND2X0 U6018 ( .IN1(P1_N106), .IN2(n6582), .QN(n4239) );
  NAND2X0 U6019 ( .IN1(n4241), .IN2(n4242), .QN(P1_N5523) );
  NAND2X0 U6020 ( .IN1(n4147), .IN2(n4169), .QN(n4242) );
  NAND2X0 U6021 ( .IN1(P1_N105), .IN2(n6582), .QN(n4241) );
  NAND2X0 U6022 ( .IN1(n4243), .IN2(n4244), .QN(P1_N5522) );
  NAND2X0 U6023 ( .IN1(n4150), .IN2(n4169), .QN(n4244) );
  NAND2X0 U6024 ( .IN1(P1_N104), .IN2(n6582), .QN(n4243) );
  NAND2X0 U6025 ( .IN1(n4245), .IN2(n4246), .QN(P1_N5521) );
  NAND2X0 U6026 ( .IN1(n4153), .IN2(n4169), .QN(n4246) );
  NAND2X0 U6027 ( .IN1(P1_N103), .IN2(n6582), .QN(n4245) );
  NAND2X0 U6028 ( .IN1(n4247), .IN2(n4248), .QN(P1_N5520) );
  NAND2X0 U6029 ( .IN1(n4156), .IN2(n6583), .QN(n4248) );
  NAND2X0 U6030 ( .IN1(n6624), .IN2(n6582), .QN(n4247) );
  NAND2X0 U6033 ( .IN1(n6713), .IN2(n6582), .QN(P1_N5548) );
  OR2X1 U6034 ( .IN2(n4251), .IN1(n7424), .Q(P1_N5517) );
  NAND2X0 U6035 ( .IN1(n4252), .IN2(n4253), .QN(n4251) );
  NAND2X0 U6036 ( .IN1(P1_N4838), .IN2(n4164), .QN(n4253) );
  NAND2X0 U6037 ( .IN1(n9661), .IN2(n6583), .QN(n4252) );
  OR2X1 U6040 ( .IN2(n4257), .IN1(n7425), .Q(P1_N5516) );
  NAND2X0 U6041 ( .IN1(n4258), .IN2(n4259), .QN(n4257) );
  NAND2X0 U6042 ( .IN1(P1_N4837), .IN2(n4164), .QN(n4259) );
  NAND2X0 U6043 ( .IN1(n9851), .IN2(n6583), .QN(n4258) );
  OR2X1 U6046 ( .IN2(n4262), .IN1(n7426), .Q(P1_N5515) );
  NAND2X0 U6047 ( .IN1(n4263), .IN2(n4264), .QN(n4262) );
  NAND2X0 U6048 ( .IN1(P1_N4836), .IN2(n4164), .QN(n4264) );
  NAND2X0 U6049 ( .IN1(n9665), .IN2(n6583), .QN(n4263) );
  OR2X1 U6052 ( .IN2(n4267), .IN1(n7427), .Q(P1_N5514) );
  NAND2X0 U6053 ( .IN1(n4268), .IN2(n4269), .QN(n4267) );
  NAND2X0 U6054 ( .IN1(P1_N4835), .IN2(n4164), .QN(n4269) );
  NAND2X0 U6055 ( .IN1(n9855), .IN2(n6583), .QN(n4268) );
  NOR2X0 U5866 ( .QN(P1_N661), .IN1(n4084), .IN2(n7027) );
  NOR2X0 U5867 ( .QN(P1_N660), .IN1(n4086), .IN2(n7027) );
  NOR2X0 U5868 ( .QN(P1_N659), .IN1(n7328), .IN2(n7029) );
  NOR2X0 U5869 ( .QN(P1_N658), .IN1(n7326), .IN2(n7029) );
  NOR2X0 U5870 ( .QN(P1_N657), .IN1(n7324), .IN2(n7029) );
  NOR2X0 U5871 ( .QN(P1_N656), .IN1(n7322), .IN2(n7029) );
  NOR2X0 U5872 ( .QN(P1_N655), .IN1(n7320), .IN2(n7029) );
  NOR2X0 U5873 ( .QN(P1_N654), .IN1(n7318), .IN2(n7029) );
  NOR2X0 U5874 ( .QN(P1_N653), .IN1(n7316), .IN2(n7029) );
  NOR2X0 U5875 ( .QN(P1_N652), .IN1(n7314), .IN2(n7027) );
  NOR2X0 U5876 ( .QN(P1_N651), .IN1(n7312), .IN2(n7027) );
  NOR2X0 U5877 ( .QN(P1_N650), .IN1(n7310), .IN2(n7023) );
  NAND2X0 U5879 ( .IN1(n4097), .IN2(n4098), .QN(P1_N649) );
  NAND2X0 U5880 ( .IN1(n7019), .IN2(n4099), .QN(n4098) );
  NAND2X0 U5881 ( .IN1(n4100), .IN2(n4101), .QN(P1_N648) );
  NAND2X0 U5882 ( .IN1(n7028), .IN2(n4102), .QN(n4101) );
  NAND2X0 U5883 ( .IN1(n4103), .IN2(n4104), .QN(P1_N647) );
  NAND2X0 U5884 ( .IN1(n7028), .IN2(n4105), .QN(n4104) );
  NAND2X0 U5885 ( .IN1(n4106), .IN2(n4107), .QN(P1_N646) );
  NAND2X0 U5886 ( .IN1(n7028), .IN2(n4108), .QN(n4107) );
  NAND2X0 U5887 ( .IN1(n4109), .IN2(n4110), .QN(P1_N645) );
  NAND2X0 U5888 ( .IN1(n7028), .IN2(n4111), .QN(n4110) );
  NAND2X0 U5889 ( .IN1(n4112), .IN2(n4113), .QN(P1_N644) );
  NAND2X0 U5890 ( .IN1(n7028), .IN2(n4114), .QN(n4113) );
  NAND2X0 U5891 ( .IN1(n4115), .IN2(n4116), .QN(P1_N643) );
  NAND2X0 U5892 ( .IN1(n7028), .IN2(n4117), .QN(n4116) );
  NAND2X0 U5893 ( .IN1(n4118), .IN2(n4119), .QN(P1_N642) );
  NAND2X0 U5894 ( .IN1(n7024), .IN2(n4120), .QN(n4119) );
  NAND2X0 U5895 ( .IN1(n4121), .IN2(n4122), .QN(P1_N641) );
  NAND2X0 U5896 ( .IN1(n7024), .IN2(n4123), .QN(n4122) );
  NAND2X0 U5897 ( .IN1(n4124), .IN2(n4125), .QN(P1_N640) );
  NAND2X0 U5898 ( .IN1(n7463), .IN2(n4126), .QN(n4125) );
  NAND2X0 U5899 ( .IN1(n4127), .IN2(n4128), .QN(P1_N639) );
  NAND2X0 U5900 ( .IN1(n7463), .IN2(n4129), .QN(n4128) );
  NAND2X0 U5901 ( .IN1(n4130), .IN2(n4131), .QN(P1_N638) );
  NAND2X0 U5902 ( .IN1(n7463), .IN2(n4132), .QN(n4131) );
  NAND2X0 U5903 ( .IN1(n4133), .IN2(n4134), .QN(P1_N637) );
  NAND2X0 U5904 ( .IN1(n7463), .IN2(n4135), .QN(n4134) );
  NAND2X0 U5905 ( .IN1(n4136), .IN2(n4137), .QN(P1_N636) );
  NAND2X0 U5906 ( .IN1(n7463), .IN2(n4138), .QN(n4137) );
  NAND2X0 U5907 ( .IN1(n4139), .IN2(n4140), .QN(P1_N635) );
  NAND2X0 U5908 ( .IN1(n7026), .IN2(n4141), .QN(n4140) );
  NAND2X0 U5909 ( .IN1(n4142), .IN2(n4143), .QN(P1_N634) );
  NAND2X0 U5910 ( .IN1(n7026), .IN2(n4144), .QN(n4143) );
  NAND2X0 U5911 ( .IN1(n4145), .IN2(n4146), .QN(P1_N633) );
  NAND2X0 U5912 ( .IN1(n7026), .IN2(n4147), .QN(n4146) );
  NAND2X0 U5913 ( .IN1(n4148), .IN2(n4149), .QN(P1_N632) );
  NAND2X0 U5914 ( .IN1(n7026), .IN2(n4150), .QN(n4149) );
  NAND2X0 U5915 ( .IN1(n4151), .IN2(n4152), .QN(P1_N631) );
  NAND2X0 U5916 ( .IN1(n7026), .IN2(n4153), .QN(n4152) );
  NAND2X0 U5917 ( .IN1(n4154), .IN2(n4155), .QN(P1_N630) );
  NAND2X0 U5918 ( .IN1(n7026), .IN2(n4156), .QN(n4155) );
  NAND2X0 U5921 ( .IN1(n7330), .IN2(n4157), .QN(P1_N584) );
  AND2X1 U5924 ( .IN1(P1_N4905), .IN2(n4164), .Q(P1_N5564) );
  AND2X1 U5925 ( .IN1(P1_N4872), .IN2(n4164), .Q(P1_N5563) );
  AND2X1 U5926 ( .IN1(P1_N4839), .IN2(n4164), .Q(P1_N5562) );
  NAND2X0 U5927 ( .IN1(n6927), .IN2(n4166), .QN(P1_N5561) );
  NAND2X0 U5928 ( .IN1(n4167), .IN2(n4168), .QN(n4166) );
  AND2X1 U5929 ( .IN1(n7340), .IN2(n7414), .Q(n4168) );
  NOR2X0 U5930 ( .QN(n4167), .IN1(n6580), .IN2(n7419) );
  AND2X1 U5933 ( .IN1(n4164), .IN2(P1_N536), .Q(P1_N5560) );
  AND2X1 U5934 ( .IN1(n4172), .IN2(P1_N4969), .Q(P1_N5554) );
  NAND2X0 U5935 ( .IN1(n4173), .IN2(n4174), .QN(P1_N5553) );
  NAND2X0 U5936 ( .IN1(n4175), .IN2(n6583), .QN(n4174) );
  NAND2X0 U5937 ( .IN1(P1_N133), .IN2(n6584), .QN(n4173) );
  NAND2X0 U5938 ( .IN1(n4176), .IN2(n4177), .QN(P1_N5552) );
  NAND2X0 U5939 ( .IN1(n4178), .IN2(n6580), .QN(n4177) );
  NAND2X0 U5940 ( .IN1(P1_N132), .IN2(n6584), .QN(n4176) );
  NAND2X0 U5941 ( .IN1(n4179), .IN2(n4180), .QN(P1_N5551) );
  NAND2X0 U5942 ( .IN1(n4181), .IN2(n6580), .QN(n4180) );
  NAND2X0 U5943 ( .IN1(P1_N131), .IN2(n6584), .QN(n4179) );
  NAND2X0 U5944 ( .IN1(n4182), .IN2(n4183), .QN(P1_N5550) );
  NAND2X0 U5945 ( .IN1(n4184), .IN2(n6580), .QN(n4183) );
  NAND2X0 U5946 ( .IN1(P1_N130), .IN2(n6584), .QN(n4182) );
  NAND2X0 U5947 ( .IN1(n4185), .IN2(n4186), .QN(P1_N5549) );
  NAND2X0 U5948 ( .IN1(n4187), .IN2(n6580), .QN(n4186) );
  NAND2X0 U5949 ( .IN1(P1_N129), .IN2(n6584), .QN(n4185) );
  NAND2X0 U5950 ( .IN1(n4188), .IN2(n4189), .QN(P1_N5547) );
  NAND2X0 U5951 ( .IN1(n4190), .IN2(n6580), .QN(n4189) );
  NAND2X0 U5952 ( .IN1(P1_N128), .IN2(n6584), .QN(n4188) );
  NAND2X0 U5953 ( .IN1(n4191), .IN2(n4192), .QN(P1_N5546) );
  NAND2X0 U5954 ( .IN1(n4193), .IN2(n6580), .QN(n4192) );
  NAND2X0 U5955 ( .IN1(P1_N127), .IN2(n6584), .QN(n4191) );
  NAND2X0 U5956 ( .IN1(n4194), .IN2(n4195), .QN(P1_N5545) );
  NAND2X0 U5957 ( .IN1(n4196), .IN2(n6580), .QN(n4195) );
  NAND2X0 U5958 ( .IN1(P1_N126), .IN2(n6584), .QN(n4194) );
  NAND2X0 U5959 ( .IN1(n4197), .IN2(n4198), .QN(P1_N5544) );
  NAND2X0 U5768 ( .IN1(n4020), .IN2(n4021), .QN(P1_N967) );
  NAND2X0 U5769 ( .IN1(P1_N908), .IN2(n4022), .QN(n4021) );
  NAND2X0 U5770 ( .IN1(P1_N392), .IN2(P1_N5576), .QN(n4020) );
  NAND2X0 U5771 ( .IN1(n4024), .IN2(n4025), .QN(P1_N966) );
  NAND2X0 U5772 ( .IN1(P1_N907), .IN2(n4022), .QN(n4025) );
  NAND2X0 U5773 ( .IN1(P1_N391), .IN2(P1_N5576), .QN(n4024) );
  NAND2X0 U5774 ( .IN1(n4026), .IN2(n4027), .QN(P1_N965) );
  NAND2X0 U5775 ( .IN1(P1_N906), .IN2(n4022), .QN(n4027) );
  NAND2X0 U5776 ( .IN1(P1_N390), .IN2(P1_N5576), .QN(n4026) );
  NAND2X0 U5777 ( .IN1(n4028), .IN2(n4029), .QN(P1_N964) );
  NAND2X0 U5778 ( .IN1(P1_N905), .IN2(n4022), .QN(n4029) );
  NAND2X0 U5779 ( .IN1(P1_N389), .IN2(P1_N5576), .QN(n4028) );
  NAND2X0 U5780 ( .IN1(n4030), .IN2(n4031), .QN(P1_N963) );
  NAND2X0 U5781 ( .IN1(P1_N904), .IN2(n4022), .QN(n4031) );
  NAND2X0 U5782 ( .IN1(P1_N388), .IN2(P1_N5576), .QN(n4030) );
  NAND2X0 U5783 ( .IN1(n4032), .IN2(n4033), .QN(P1_N962) );
  NAND2X0 U5784 ( .IN1(P1_N903), .IN2(n4022), .QN(n4033) );
  NAND2X0 U5785 ( .IN1(P1_N387), .IN2(P1_N5576), .QN(n4032) );
  NAND2X0 U5786 ( .IN1(n4034), .IN2(n4035), .QN(P1_N961) );
  NAND2X0 U5787 ( .IN1(P1_N902), .IN2(n4022), .QN(n4035) );
  NAND2X0 U5788 ( .IN1(P1_N386), .IN2(P1_N5576), .QN(n4034) );
  NAND2X0 U5789 ( .IN1(n4036), .IN2(n4037), .QN(P1_N960) );
  NAND2X0 U5790 ( .IN1(P1_N901), .IN2(n4022), .QN(n4037) );
  NAND2X0 U5791 ( .IN1(P1_N385), .IN2(P1_N5576), .QN(n4036) );
  NAND2X0 U5792 ( .IN1(n4038), .IN2(n4039), .QN(P1_N959) );
  NAND2X0 U5793 ( .IN1(P1_N900), .IN2(n4022), .QN(n4039) );
  NAND2X0 U5794 ( .IN1(P1_N384), .IN2(P1_N5576), .QN(n4038) );
  NAND2X0 U5795 ( .IN1(n4040), .IN2(n4041), .QN(P1_N958) );
  NAND2X0 U5796 ( .IN1(P1_N899), .IN2(n4022), .QN(n4041) );
  NAND2X0 U5797 ( .IN1(P1_N383), .IN2(P1_N5576), .QN(n4040) );
  NAND2X0 U5798 ( .IN1(n4042), .IN2(n4043), .QN(P1_N957) );
  NAND2X0 U5799 ( .IN1(P1_N898), .IN2(n4022), .QN(n4043) );
  NAND2X0 U5800 ( .IN1(P1_N382), .IN2(P1_N5576), .QN(n4042) );
  NAND2X0 U5801 ( .IN1(n4044), .IN2(n4045), .QN(P1_N956) );
  NAND2X0 U5802 ( .IN1(P1_N897), .IN2(n4022), .QN(n4045) );
  NAND2X0 U5803 ( .IN1(P1_N381), .IN2(P1_N5576), .QN(n4044) );
  NAND2X0 U5804 ( .IN1(n4046), .IN2(n4047), .QN(P1_N955) );
  NAND2X0 U5805 ( .IN1(P1_N896), .IN2(n4022), .QN(n4047) );
  NAND2X0 U5806 ( .IN1(P1_N380), .IN2(P1_N5576), .QN(n4046) );
  NAND2X0 U5807 ( .IN1(n4048), .IN2(n4049), .QN(P1_N954) );
  NAND2X0 U5808 ( .IN1(P1_N895), .IN2(n4022), .QN(n4049) );
  NAND2X0 U5809 ( .IN1(P1_N379), .IN2(P1_N5576), .QN(n4048) );
  NAND2X0 U5810 ( .IN1(n4050), .IN2(n4051), .QN(P1_N953) );
  NAND2X0 U5811 ( .IN1(P1_N894), .IN2(n4022), .QN(n4051) );
  NAND2X0 U5812 ( .IN1(P1_N378), .IN2(P1_N5576), .QN(n4050) );
  NAND2X0 U5813 ( .IN1(n4052), .IN2(n4053), .QN(P1_N952) );
  NAND2X0 U5814 ( .IN1(P1_N893), .IN2(n4022), .QN(n4053) );
  NAND2X0 U5815 ( .IN1(P1_N377), .IN2(P1_N5576), .QN(n4052) );
  NAND2X0 U5816 ( .IN1(n4054), .IN2(n4055), .QN(P1_N951) );
  NAND2X0 U5817 ( .IN1(P1_N892), .IN2(n4022), .QN(n4055) );
  NAND2X0 U5818 ( .IN1(P1_N376), .IN2(P1_N5576), .QN(n4054) );
  NAND2X0 U5819 ( .IN1(n4056), .IN2(n4057), .QN(P1_N950) );
  NAND2X0 U5820 ( .IN1(P1_N891), .IN2(n4022), .QN(n4057) );
  NAND2X0 U5821 ( .IN1(P1_N375), .IN2(P1_N5576), .QN(n4056) );
  NAND2X0 U5822 ( .IN1(n4058), .IN2(n4059), .QN(P1_N949) );
  NAND2X0 U5823 ( .IN1(P1_N890), .IN2(n4022), .QN(n4059) );
  NAND2X0 U5824 ( .IN1(P1_N374), .IN2(P1_N5576), .QN(n4058) );
  NAND2X0 U5825 ( .IN1(n4060), .IN2(n4061), .QN(P1_N948) );
  NAND2X0 U5826 ( .IN1(P1_N889), .IN2(n4022), .QN(n4061) );
  NAND2X0 U5827 ( .IN1(P1_N373), .IN2(P1_N5576), .QN(n4060) );
  NAND2X0 U5828 ( .IN1(n4062), .IN2(n4063), .QN(P1_N947) );
  NAND2X0 U5829 ( .IN1(P1_N888), .IN2(n4022), .QN(n4063) );
  NAND2X0 U5830 ( .IN1(P1_N372), .IN2(P1_N5576), .QN(n4062) );
  NAND2X0 U5831 ( .IN1(n4064), .IN2(n4065), .QN(P1_N946) );
  NAND2X0 U5832 ( .IN1(P1_N887), .IN2(n4022), .QN(n4065) );
  NAND2X0 U5833 ( .IN1(P1_N371), .IN2(P1_N5576), .QN(n4064) );
  NAND2X0 U5834 ( .IN1(n4066), .IN2(n4067), .QN(P1_N945) );
  NAND2X0 U5835 ( .IN1(P1_N886), .IN2(n4022), .QN(n4067) );
  NAND2X0 U5836 ( .IN1(P1_N370), .IN2(P1_N5576), .QN(n4066) );
  NAND2X0 U5837 ( .IN1(n4068), .IN2(n4069), .QN(P1_N944) );
  NAND2X0 U5838 ( .IN1(P1_N885), .IN2(n4022), .QN(n4069) );
  NAND2X0 U5839 ( .IN1(P1_N369), .IN2(P1_N5576), .QN(n4068) );
  NAND2X0 U5840 ( .IN1(n4070), .IN2(n4071), .QN(P1_N943) );
  NAND2X0 U5841 ( .IN1(P1_N884), .IN2(n4022), .QN(n4071) );
  NAND2X0 U5842 ( .IN1(P1_N368), .IN2(P1_N5576), .QN(n4070) );
  NAND2X0 U5843 ( .IN1(n4072), .IN2(n4073), .QN(P1_N942) );
  NAND2X0 U5844 ( .IN1(P1_N883), .IN2(n4022), .QN(n4073) );
  NAND2X0 U5845 ( .IN1(n18451), .IN2(P1_N5576), .QN(n4072) );
  NAND2X0 U5846 ( .IN1(n4074), .IN2(n4075), .QN(P1_N941) );
  NAND2X0 U5847 ( .IN1(P1_N882), .IN2(n4022), .QN(n4075) );
  NAND2X0 U5848 ( .IN1(n6623), .IN2(P1_N5576), .QN(n4074) );
  NAND2X0 U5849 ( .IN1(n4076), .IN2(n4077), .QN(P1_N940) );
  NAND2X0 U5850 ( .IN1(P1_N881), .IN2(n4022), .QN(n4077) );
  NAND2X0 U5851 ( .IN1(n6622), .IN2(P1_N5576), .QN(n4076) );
  NAND2X0 U5852 ( .IN1(n4078), .IN2(n4079), .QN(P1_N939) );
  NAND2X0 U5853 ( .IN1(P1_N630), .IN2(n4022), .QN(n4079) );
  NAND2X0 U5856 ( .IN1(n6621), .IN2(P1_N5576), .QN(n4078) );
  NAND2X0 U5861 ( .IN1(n7376), .IN2(n4082), .QN(P1_N781) );
  NAND2X0 U5862 ( .IN1(n7375), .IN2(n4083), .QN(P1_N779) );
  NOR2X0 U5863 ( .QN(P1_N968), .IN1(n4083), .IN2(n4082) );
  INVX0 U5864 ( .ZN(n4082), .INP(n7375) );
  INVX0 U5865 ( .ZN(n4083), .INP(n7376) );
  AND2X1 U5672 ( .IN1(n3957), .IN2(n3958), .Q(n3955) );
  NAND2X0 U5673 ( .IN1(n6999), .IN2(P2_N351), .QN(n3958) );
  NAND2X0 U5674 ( .IN1(n123), .IN2(n7334), .QN(n3957) );
  NAND2X0 U5675 ( .IN1(n3959), .IN2(n3960), .QN(P2_N926) );
  NAND2X0 U5676 ( .IN1(n103), .IN2(n7341), .QN(n3960) );
  AND2X1 U5677 ( .IN1(n3961), .IN2(n3962), .Q(n3959) );
  NAND2X0 U5678 ( .IN1(n6999), .IN2(P2_N352), .QN(n3962) );
  NAND2X0 U5679 ( .IN1(n124), .IN2(n7334), .QN(n3961) );
  NAND2X0 U5681 ( .IN1(n104), .IN2(n7341), .QN(n3964) );
  AND2X1 U5682 ( .IN1(n3965), .IN2(n3966), .Q(n3963) );
  NAND2X0 U5683 ( .IN1(n6999), .IN2(P2_N353), .QN(n3966) );
  NAND2X0 U5684 ( .IN1(n125), .IN2(n7334), .QN(n3965) );
  NAND2X0 U5685 ( .IN1(n3967), .IN2(n3968), .QN(P2_N924) );
  NAND2X0 U5686 ( .IN1(n105), .IN2(n7341), .QN(n3968) );
  AND2X1 U5687 ( .IN1(n3969), .IN2(n3970), .Q(n3967) );
  NAND2X0 U5688 ( .IN1(n6999), .IN2(P2_N354), .QN(n3970) );
  NAND2X0 U5689 ( .IN1(n126), .IN2(n7334), .QN(n3969) );
  NAND2X0 U5690 ( .IN1(n3971), .IN2(n3972), .QN(P2_N923) );
  NAND2X0 U5691 ( .IN1(n106), .IN2(n7341), .QN(n3972) );
  AND2X1 U5692 ( .IN1(n3973), .IN2(n3974), .Q(n3971) );
  NAND2X0 U5693 ( .IN1(n6999), .IN2(P2_N355), .QN(n3974) );
  NAND2X0 U5694 ( .IN1(n127), .IN2(n7334), .QN(n3973) );
  NAND2X0 U5695 ( .IN1(n3975), .IN2(n3976), .QN(P2_N922) );
  NAND2X0 U5696 ( .IN1(n107), .IN2(n7341), .QN(n3976) );
  AND2X1 U5697 ( .IN1(n3977), .IN2(n3978), .Q(n3975) );
  NAND2X0 U5698 ( .IN1(n6999), .IN2(P2_N356), .QN(n3978) );
  NAND2X0 U5699 ( .IN1(n128), .IN2(n7334), .QN(n3977) );
  NAND2X0 U5700 ( .IN1(n3979), .IN2(n3980), .QN(P2_N921) );
  NAND2X0 U5701 ( .IN1(n108), .IN2(n7341), .QN(n3980) );
  AND2X1 U5702 ( .IN1(n3981), .IN2(n3982), .Q(n3979) );
  NAND2X0 U5703 ( .IN1(n6999), .IN2(P2_N357), .QN(n3982) );
  NAND2X0 U5704 ( .IN1(n129), .IN2(n7334), .QN(n3981) );
  NAND2X0 U5705 ( .IN1(n3983), .IN2(n3984), .QN(P2_N920) );
  NAND2X0 U5706 ( .IN1(n109), .IN2(n7341), .QN(n3984) );
  AND2X1 U5707 ( .IN1(n3985), .IN2(n3986), .Q(n3983) );
  NAND2X0 U5708 ( .IN1(n6999), .IN2(P2_N358), .QN(n3986) );
  NAND2X0 U5709 ( .IN1(n130), .IN2(n7334), .QN(n3985) );
  NAND2X0 U5710 ( .IN1(n3987), .IN2(n3988), .QN(P2_N919) );
  NAND2X0 U5711 ( .IN1(n110), .IN2(n7341), .QN(n3988) );
  AND2X1 U5712 ( .IN1(n3989), .IN2(n3990), .Q(n3987) );
  NAND2X0 U5713 ( .IN1(n6999), .IN2(P2_N359), .QN(n3990) );
  NAND2X0 U5714 ( .IN1(n131), .IN2(n7334), .QN(n3989) );
  NAND2X0 U5715 ( .IN1(n3991), .IN2(n3992), .QN(P2_N918) );
  NAND2X0 U5716 ( .IN1(n111), .IN2(n7341), .QN(n3992) );
  AND2X1 U5717 ( .IN1(n3993), .IN2(n3994), .Q(n3991) );
  NAND2X0 U5718 ( .IN1(n6999), .IN2(P2_N360), .QN(n3994) );
  NAND2X0 U5719 ( .IN1(n132), .IN2(n7334), .QN(n3993) );
  NAND2X0 U5720 ( .IN1(n3995), .IN2(n3996), .QN(P2_N917) );
  NAND2X0 U5721 ( .IN1(n112), .IN2(n7341), .QN(n3996) );
  AND2X1 U5722 ( .IN1(n3997), .IN2(n3998), .Q(n3995) );
  NAND2X0 U5723 ( .IN1(n6999), .IN2(P2_N361), .QN(n3998) );
  NAND2X0 U5724 ( .IN1(n133), .IN2(n7334), .QN(n3997) );
  NAND2X0 U5725 ( .IN1(n3999), .IN2(n4000), .QN(P2_N916) );
  NAND2X0 U5726 ( .IN1(n113), .IN2(n7341), .QN(n4000) );
  AND2X1 U5727 ( .IN1(n4001), .IN2(n4002), .Q(n3999) );
  NAND2X0 U5728 ( .IN1(n6999), .IN2(P2_N362), .QN(n4002) );
  NAND2X0 U5729 ( .IN1(n134), .IN2(n7334), .QN(n4001) );
  NAND2X0 U5730 ( .IN1(n4003), .IN2(n4004), .QN(P2_N915) );
  NAND2X0 U5731 ( .IN1(n114), .IN2(n7341), .QN(n4004) );
  AND2X1 U5732 ( .IN1(n4005), .IN2(n4006), .Q(n4003) );
  NAND2X0 U5733 ( .IN1(n6999), .IN2(P2_N363), .QN(n4006) );
  NAND2X0 U5734 ( .IN1(n135), .IN2(n7334), .QN(n4005) );
  NOR2X0 U5735 ( .QN(P2_N1005), .IN1(n7329), .IN2(n7007) );
  NAND2X0 U5737 ( .IN1(n4007), .IN2(n4008), .QN(n2178) );
  NAND2X0 U5738 ( .IN1(N68), .IN2(n6739), .QN(n4008) );
  NAND2X0 U5739 ( .IN1(n10095), .IN2(N5), .QN(n4007) );
  NOR2X0 U5740 ( .QN(P2_N1004), .IN1(n7013), .IN2(n7327) );
  NAND2X0 U5742 ( .IN1(n4009), .IN2(n4010), .QN(n2181) );
  NAND2X0 U5743 ( .IN1(N67), .IN2(n6739), .QN(n4010) );
  NAND2X0 U5744 ( .IN1(n9935), .IN2(N5), .QN(n4009) );
  NOR2X0 U5745 ( .QN(P2_N1003), .IN1(n7015), .IN2(n7325) );
  NAND2X0 U5747 ( .IN1(n4011), .IN2(n4012), .QN(n2184) );
  NAND2X0 U5748 ( .IN1(N66), .IN2(n6739), .QN(n4012) );
  NAND2X0 U5749 ( .IN1(n9939), .IN2(N5), .QN(n4011) );
  NOR2X0 U5750 ( .QN(P2_N1002), .IN1(n7015), .IN2(n7323) );
  NAND2X0 U5752 ( .IN1(n4013), .IN2(n4014), .QN(n2187) );
  NAND2X0 U5753 ( .IN1(N65), .IN2(n6739), .QN(n4014) );
  NAND2X0 U5754 ( .IN1(n9943), .IN2(N5), .QN(n4013) );
  NOR2X0 U5755 ( .QN(P2_N1001), .IN1(n7015), .IN2(n7321) );
  NAND2X0 U5757 ( .IN1(n4015), .IN2(n4016), .QN(n2190) );
  NAND2X0 U5758 ( .IN1(N64), .IN2(n6739), .QN(n4016) );
  NAND2X0 U5759 ( .IN1(n9947), .IN2(N5), .QN(n4015) );
  NOR2X0 U5760 ( .QN(P2_N1000), .IN1(n7015), .IN2(n7319) );
  NAND2X0 U5762 ( .IN1(n4017), .IN2(n4018), .QN(n2193) );
  NAND2X0 U5763 ( .IN1(N63), .IN2(n6739), .QN(n4018) );
  NAND2X0 U5764 ( .IN1(n9951), .IN2(N5), .QN(n4017) );
  NAND2X0 U5574 ( .IN1(P2_N358), .IN2(n2693), .QN(n2048) );
  NAND2X0 U5575 ( .IN1(P2_N369), .IN2(P2_N5495), .QN(n3893) );
  NAND2X0 U5576 ( .IN1(n3898), .IN2(n3899), .QN(P2_N1163) );
  NAND2X0 U5577 ( .IN1(n3796), .IN2(P2_N980), .QN(n3899) );
  NAND2X0 U5578 ( .IN1(n2051), .IN2(n3900), .QN(P2_N980) );
  NAND2X0 U5579 ( .IN1(n7462), .IN2(n2053), .QN(n3900) );
  NAND2X0 U5580 ( .IN1(n3901), .IN2(n3902), .QN(n2053) );
  NAND2X0 U5581 ( .IN1(N43), .IN2(n6737), .QN(n3902) );
  NAND2X0 U5582 ( .IN1(n9891), .IN2(n6736), .QN(n3901) );
  NAND2X0 U5583 ( .IN1(P2_N359), .IN2(n2693), .QN(n2051) );
  NAND2X0 U5584 ( .IN1(P2_N368), .IN2(P2_N5495), .QN(n3898) );
  NAND2X0 U5585 ( .IN1(n3903), .IN2(n3904), .QN(P2_N1162) );
  NAND2X0 U5586 ( .IN1(n3796), .IN2(P2_N979), .QN(n3904) );
  NAND2X0 U5587 ( .IN1(n2054), .IN2(n3905), .QN(P2_N979) );
  NAND2X0 U5588 ( .IN1(n7462), .IN2(n2056), .QN(n3905) );
  NAND2X0 U5589 ( .IN1(n3906), .IN2(n3907), .QN(n2056) );
  NAND2X0 U5590 ( .IN1(N42), .IN2(n6737), .QN(n3907) );
  NAND2X0 U5591 ( .IN1(n9895), .IN2(n6736), .QN(n3906) );
  NAND2X0 U5592 ( .IN1(P2_N360), .IN2(n2693), .QN(n2054) );
  NAND2X0 U5593 ( .IN1(n18813), .IN2(P2_N5495), .QN(n3903) );
  NAND2X0 U5594 ( .IN1(n3908), .IN2(n3909), .QN(P2_N1161) );
  NAND2X0 U5595 ( .IN1(n3796), .IN2(P2_N978), .QN(n3909) );
  NAND2X0 U5596 ( .IN1(n2057), .IN2(n3910), .QN(P2_N978) );
  NAND2X0 U5597 ( .IN1(n7462), .IN2(n2059), .QN(n3910) );
  NAND2X0 U5598 ( .IN1(n3911), .IN2(n3912), .QN(n2059) );
  NAND2X0 U5599 ( .IN1(N41), .IN2(n6737), .QN(n3912) );
  NAND2X0 U5600 ( .IN1(n9899), .IN2(n6736), .QN(n3911) );
  NAND2X0 U5601 ( .IN1(P2_N361), .IN2(n2693), .QN(n2057) );
  NAND2X0 U5602 ( .IN1(n6683), .IN2(P2_N5495), .QN(n3908) );
  NAND2X0 U5603 ( .IN1(n3913), .IN2(n3914), .QN(P2_N1160) );
  NAND2X0 U5604 ( .IN1(n3796), .IN2(P2_N977), .QN(n3914) );
  NAND2X0 U5605 ( .IN1(n2060), .IN2(n3915), .QN(P2_N977) );
  NAND2X0 U5606 ( .IN1(n7462), .IN2(n2062), .QN(n3915) );
  NAND2X0 U5607 ( .IN1(n3916), .IN2(n3917), .QN(n2062) );
  NAND2X0 U5608 ( .IN1(N40), .IN2(n6737), .QN(n3917) );
  NAND2X0 U5609 ( .IN1(n9333), .IN2(n6736), .QN(n3916) );
  NAND2X0 U5610 ( .IN1(P2_N362), .IN2(n2693), .QN(n2060) );
  NAND2X0 U5611 ( .IN1(n6682), .IN2(P2_N5495), .QN(n3913) );
  NAND2X0 U5612 ( .IN1(n3918), .IN2(n3919), .QN(P2_N1159) );
  NAND2X0 U5613 ( .IN1(n3796), .IN2(P2_N976), .QN(n3919) );
  NAND2X0 U5614 ( .IN1(n2063), .IN2(n3920), .QN(P2_N976) );
  NAND2X0 U5615 ( .IN1(n7462), .IN2(n2065), .QN(n3920) );
  NAND2X0 U5616 ( .IN1(n3921), .IN2(n3922), .QN(n2065) );
  NAND2X0 U5617 ( .IN1(N39), .IN2(n6737), .QN(n3922) );
  NAND2X0 U5618 ( .IN1(n9385), .IN2(n6736), .QN(n3921) );
  NAND2X0 U5619 ( .IN1(P2_N363), .IN2(n2693), .QN(n2063) );
  INVX0 U5621 ( .ZN(n2154), .INP(n7332) );
  INVX0 U5622 ( .ZN(n2153), .INP(n7333) );
  NAND2X0 U5625 ( .IN1(n6681), .IN2(P2_N5495), .QN(n3918) );
  NAND2X0 U5630 ( .IN1(n7378), .IN2(n3925), .QN(P2_N1126) );
  NAND2X0 U5631 ( .IN1(n7377), .IN2(n3926), .QN(P2_N1124) );
  NOR2X0 U5632 ( .QN(P2_N1188), .IN1(n3926), .IN2(n3925) );
  INVX0 U5633 ( .ZN(n3925), .INP(n7377) );
  INVX0 U5634 ( .ZN(n3926), .INP(n7378) );
  NAND2X0 U5635 ( .IN1(n3927), .IN2(n3928), .QN(P2_N934) );
  NAND2X0 U5636 ( .IN1(n95), .IN2(n7341), .QN(n3928) );
  AND2X1 U5637 ( .IN1(n3929), .IN2(n3930), .Q(n3927) );
  NAND2X0 U5638 ( .IN1(n6999), .IN2(P2_N344), .QN(n3930) );
  NAND2X0 U5639 ( .IN1(n116), .IN2(n7334), .QN(n3929) );
  NAND2X0 U5640 ( .IN1(n3931), .IN2(n3932), .QN(P2_N933) );
  NAND2X0 U5641 ( .IN1(n96), .IN2(n7341), .QN(n3932) );
  AND2X1 U5642 ( .IN1(n3933), .IN2(n3934), .Q(n3931) );
  NAND2X0 U5643 ( .IN1(n6999), .IN2(P2_N345), .QN(n3934) );
  NAND2X0 U5644 ( .IN1(n117), .IN2(n7334), .QN(n3933) );
  NAND2X0 U5645 ( .IN1(n3935), .IN2(n3936), .QN(P2_N932) );
  NAND2X0 U5646 ( .IN1(n97), .IN2(n7341), .QN(n3936) );
  AND2X1 U5647 ( .IN1(n3937), .IN2(n3938), .Q(n3935) );
  NAND2X0 U5648 ( .IN1(n6999), .IN2(P2_N346), .QN(n3938) );
  NAND2X0 U5649 ( .IN1(n118), .IN2(n7334), .QN(n3937) );
  NAND2X0 U5650 ( .IN1(n3939), .IN2(n3940), .QN(P2_N931) );
  NAND2X0 U5651 ( .IN1(n98), .IN2(n7341), .QN(n3940) );
  AND2X1 U5652 ( .IN1(n3941), .IN2(n3942), .Q(n3939) );
  NAND2X0 U5653 ( .IN1(n6999), .IN2(P2_N347), .QN(n3942) );
  NAND2X0 U5654 ( .IN1(n119), .IN2(n7334), .QN(n3941) );
  NAND2X0 U5655 ( .IN1(n3943), .IN2(n3944), .QN(P2_N930) );
  NAND2X0 U5656 ( .IN1(n99), .IN2(n7341), .QN(n3944) );
  AND2X1 U5657 ( .IN1(n3945), .IN2(n3946), .Q(n3943) );
  NAND2X0 U5658 ( .IN1(n6999), .IN2(P2_N348), .QN(n3946) );
  NAND2X0 U5659 ( .IN1(n120), .IN2(n7334), .QN(n3945) );
  NAND2X0 U5661 ( .IN1(n100), .IN2(n7341), .QN(n3948) );
  AND2X1 U5662 ( .IN1(n3949), .IN2(n3950), .Q(n3947) );
  NAND2X0 U5663 ( .IN1(n6999), .IN2(P2_N349), .QN(n3950) );
  NAND2X0 U5664 ( .IN1(n121), .IN2(n7334), .QN(n3949) );
  NAND2X0 U5666 ( .IN1(n101), .IN2(n7341), .QN(n3952) );
  AND2X1 U5667 ( .IN1(n3953), .IN2(n3954), .Q(n3951) );
  NAND2X0 U5668 ( .IN1(n6999), .IN2(P2_N350), .QN(n3954) );
  NAND2X0 U5669 ( .IN1(n122), .IN2(n7334), .QN(n3953) );
  NAND2X0 U5670 ( .IN1(n3955), .IN2(n3956), .QN(P2_N927) );
  NAND2X0 U5671 ( .IN1(n102), .IN2(n7341), .QN(n3956) );
  NAND2X0 U5482 ( .IN1(N54), .IN2(n6737), .QN(n3847) );
  NAND2X0 U5483 ( .IN1(n9987), .IN2(n6736), .QN(n3846) );
  NAND2X0 U5484 ( .IN1(P2_N348), .IN2(n2693), .QN(n2018) );
  NAND2X0 U5485 ( .IN1(P2_N379), .IN2(P2_N5495), .QN(n3843) );
  NAND2X0 U5486 ( .IN1(n3848), .IN2(n3849), .QN(P2_N1173) );
  NAND2X0 U5487 ( .IN1(n3796), .IN2(P2_N990), .QN(n3849) );
  NAND2X0 U5488 ( .IN1(n2021), .IN2(n3850), .QN(P2_N990) );
  NAND2X0 U5489 ( .IN1(n7009), .IN2(n2023), .QN(n3850) );
  NAND2X0 U5491 ( .IN1(N53), .IN2(n6737), .QN(n3852) );
  NAND2X0 U5492 ( .IN1(n9991), .IN2(n6736), .QN(n3851) );
  NAND2X0 U5493 ( .IN1(P2_N349), .IN2(n2693), .QN(n2021) );
  NAND2X0 U5494 ( .IN1(P2_N378), .IN2(P2_N5495), .QN(n3848) );
  NAND2X0 U5495 ( .IN1(n3853), .IN2(n3854), .QN(P2_N1172) );
  NAND2X0 U5496 ( .IN1(n3796), .IN2(P2_N989), .QN(n3854) );
  NAND2X0 U5497 ( .IN1(n2024), .IN2(n3855), .QN(P2_N989) );
  NAND2X0 U5498 ( .IN1(n7009), .IN2(n2026), .QN(n3855) );
  NAND2X0 U5500 ( .IN1(N52), .IN2(n6737), .QN(n3857) );
  NAND2X0 U5501 ( .IN1(n9995), .IN2(n6736), .QN(n3856) );
  NAND2X0 U5503 ( .IN1(P2_N377), .IN2(P2_N5495), .QN(n3853) );
  NAND2X0 U5504 ( .IN1(n3858), .IN2(n3859), .QN(P2_N1171) );
  NAND2X0 U5505 ( .IN1(n3796), .IN2(P2_N988), .QN(n3859) );
  NAND2X0 U5506 ( .IN1(n2027), .IN2(n3860), .QN(P2_N988) );
  NAND2X0 U5507 ( .IN1(n7010), .IN2(n2029), .QN(n3860) );
  NAND2X0 U5509 ( .IN1(N51), .IN2(n6737), .QN(n3862) );
  NAND2X0 U5510 ( .IN1(n9999), .IN2(n6736), .QN(n3861) );
  NAND2X0 U5512 ( .IN1(P2_N376), .IN2(P2_N5495), .QN(n3858) );
  NAND2X0 U5513 ( .IN1(n3863), .IN2(n3864), .QN(P2_N1170) );
  NAND2X0 U5514 ( .IN1(n3796), .IN2(P2_N987), .QN(n3864) );
  NAND2X0 U5515 ( .IN1(n2030), .IN2(n3865), .QN(P2_N987) );
  NAND2X0 U5516 ( .IN1(n7010), .IN2(n2032), .QN(n3865) );
  NAND2X0 U5517 ( .IN1(n3866), .IN2(n3867), .QN(n2032) );
  NAND2X0 U5518 ( .IN1(N50), .IN2(n6737), .QN(n3867) );
  NAND2X0 U5519 ( .IN1(n10003), .IN2(n6736), .QN(n3866) );
  NAND2X0 U5521 ( .IN1(P2_N375), .IN2(P2_N5495), .QN(n3863) );
  NAND2X0 U5522 ( .IN1(n3868), .IN2(n3869), .QN(P2_N1169) );
  NAND2X0 U5523 ( .IN1(n3796), .IN2(P2_N986), .QN(n3869) );
  NAND2X0 U5524 ( .IN1(n2033), .IN2(n3870), .QN(P2_N986) );
  NAND2X0 U5525 ( .IN1(n7010), .IN2(n2035), .QN(n3870) );
  NAND2X0 U5526 ( .IN1(n3871), .IN2(n3872), .QN(n2035) );
  NAND2X0 U5527 ( .IN1(N49), .IN2(n6737), .QN(n3872) );
  NAND2X0 U5528 ( .IN1(n10007), .IN2(n6736), .QN(n3871) );
  NAND2X0 U5529 ( .IN1(P2_N353), .IN2(n2693), .QN(n2033) );
  NAND2X0 U5530 ( .IN1(P2_N374), .IN2(P2_N5495), .QN(n3868) );
  NAND2X0 U5531 ( .IN1(n3873), .IN2(n3874), .QN(P2_N1168) );
  NAND2X0 U5532 ( .IN1(n3796), .IN2(P2_N985), .QN(n3874) );
  NAND2X0 U5533 ( .IN1(n2036), .IN2(n3875), .QN(P2_N985) );
  NAND2X0 U5534 ( .IN1(n7010), .IN2(n2038), .QN(n3875) );
  NAND2X0 U5535 ( .IN1(n3876), .IN2(n3877), .QN(n2038) );
  NAND2X0 U5536 ( .IN1(N48), .IN2(n6737), .QN(n3877) );
  NAND2X0 U5537 ( .IN1(n9871), .IN2(n6736), .QN(n3876) );
  NAND2X0 U5538 ( .IN1(P2_N354), .IN2(n2693), .QN(n2036) );
  NAND2X0 U5539 ( .IN1(P2_N373), .IN2(P2_N5495), .QN(n3873) );
  NAND2X0 U5540 ( .IN1(n3878), .IN2(n3879), .QN(P2_N1167) );
  NAND2X0 U5541 ( .IN1(n3796), .IN2(P2_N984), .QN(n3879) );
  NAND2X0 U5542 ( .IN1(n2039), .IN2(n3880), .QN(P2_N984) );
  NAND2X0 U5543 ( .IN1(n7010), .IN2(n2041), .QN(n3880) );
  NAND2X0 U5545 ( .IN1(N47), .IN2(n6737), .QN(n3882) );
  NAND2X0 U5546 ( .IN1(n9875), .IN2(n6736), .QN(n3881) );
  NAND2X0 U5547 ( .IN1(P2_N355), .IN2(n2693), .QN(n2039) );
  NAND2X0 U5548 ( .IN1(P2_N372), .IN2(P2_N5495), .QN(n3878) );
  NAND2X0 U5549 ( .IN1(n3883), .IN2(n3884), .QN(P2_N1166) );
  NAND2X0 U5550 ( .IN1(n3796), .IN2(P2_N983), .QN(n3884) );
  NAND2X0 U5551 ( .IN1(n2042), .IN2(n3885), .QN(P2_N983) );
  NAND2X0 U5552 ( .IN1(n7010), .IN2(n2044), .QN(n3885) );
  NAND2X0 U5554 ( .IN1(N46), .IN2(n6737), .QN(n3887) );
  NAND2X0 U5555 ( .IN1(n9879), .IN2(n6736), .QN(n3886) );
  NAND2X0 U5556 ( .IN1(P2_N356), .IN2(n2693), .QN(n2042) );
  NAND2X0 U5557 ( .IN1(P2_N371), .IN2(P2_N5495), .QN(n3883) );
  NAND2X0 U5558 ( .IN1(n3888), .IN2(n3889), .QN(P2_N1165) );
  NAND2X0 U5559 ( .IN1(n3796), .IN2(P2_N982), .QN(n3889) );
  NAND2X0 U5560 ( .IN1(n2045), .IN2(n3890), .QN(P2_N982) );
  NAND2X0 U5561 ( .IN1(n7006), .IN2(n2047), .QN(n3890) );
  NAND2X0 U5562 ( .IN1(n3891), .IN2(n3892), .QN(n2047) );
  NAND2X0 U5563 ( .IN1(N45), .IN2(n6737), .QN(n3892) );
  NAND2X0 U5564 ( .IN1(n9883), .IN2(n6736), .QN(n3891) );
  NAND2X0 U5565 ( .IN1(P2_N357), .IN2(n2693), .QN(n2045) );
  NAND2X0 U5566 ( .IN1(P2_N370), .IN2(P2_N5495), .QN(n3888) );
  NAND2X0 U5567 ( .IN1(n3893), .IN2(n3894), .QN(P2_N1164) );
  NAND2X0 U5568 ( .IN1(n3796), .IN2(P2_N981), .QN(n3894) );
  NAND2X0 U5569 ( .IN1(n2048), .IN2(n3895), .QN(P2_N981) );
  NAND2X0 U5570 ( .IN1(n7006), .IN2(n2050), .QN(n3895) );
  NAND2X0 U5571 ( .IN1(n3896), .IN2(n3897), .QN(n2050) );
  NAND2X0 U5572 ( .IN1(N44), .IN2(n6737), .QN(n3897) );
  NAND2X0 U5573 ( .IN1(n9887), .IN2(n6736), .QN(n3896) );
  NAND2X0 U5386 ( .IN1(n2057), .IN2(n3790), .QN(P2_N1233) );
  NAND2X0 U5387 ( .IN1(n7462), .IN2(n2059), .QN(n3790) );
  NAND2X0 U5388 ( .IN1(n2060), .IN2(n3791), .QN(P2_N1232) );
  NAND2X0 U5389 ( .IN1(n7462), .IN2(n2062), .QN(n3791) );
  NAND2X0 U5390 ( .IN1(n2063), .IN2(n3792), .QN(P2_N1231) );
  NAND2X0 U5391 ( .IN1(n7462), .IN2(n2065), .QN(n3792) );
  NAND2X0 U5394 ( .IN1(n3794), .IN2(n3795), .QN(P2_N1187) );
  NAND2X0 U5395 ( .IN1(P2_N1004), .IN2(n3796), .QN(n3795) );
  NAND2X0 U5396 ( .IN1(P2_N392), .IN2(P2_N5495), .QN(n3794) );
  NAND2X0 U5397 ( .IN1(n3798), .IN2(n3799), .QN(P2_N1186) );
  NAND2X0 U5398 ( .IN1(P2_N1003), .IN2(n3796), .QN(n3799) );
  NAND2X0 U5399 ( .IN1(P2_N391), .IN2(P2_N5495), .QN(n3798) );
  NAND2X0 U5400 ( .IN1(n3800), .IN2(n3801), .QN(P2_N1185) );
  NAND2X0 U5401 ( .IN1(P2_N1002), .IN2(n3796), .QN(n3801) );
  NAND2X0 U5402 ( .IN1(P2_N390), .IN2(P2_N5495), .QN(n3800) );
  NAND2X0 U5403 ( .IN1(n3802), .IN2(n3803), .QN(P2_N1184) );
  NAND2X0 U5404 ( .IN1(P2_N1001), .IN2(n3796), .QN(n3803) );
  NAND2X0 U5405 ( .IN1(P2_N389), .IN2(P2_N5495), .QN(n3802) );
  NAND2X0 U5406 ( .IN1(n3804), .IN2(n3805), .QN(P2_N1183) );
  NAND2X0 U5407 ( .IN1(P2_N1000), .IN2(n3796), .QN(n3805) );
  NAND2X0 U5408 ( .IN1(P2_N388), .IN2(P2_N5495), .QN(n3804) );
  NAND2X0 U5409 ( .IN1(n3806), .IN2(n3807), .QN(P2_N1182) );
  NAND2X0 U5410 ( .IN1(P2_N999), .IN2(n3796), .QN(n3807) );
  NOR2X0 U5411 ( .QN(P2_N999), .IN1(n7015), .IN2(n7317) );
  NAND2X0 U5413 ( .IN1(n3809), .IN2(n3810), .QN(n2196) );
  NAND2X0 U5414 ( .IN1(N62), .IN2(n6739), .QN(n3810) );
  NAND2X0 U5415 ( .IN1(n9955), .IN2(N5), .QN(n3809) );
  NAND2X0 U5416 ( .IN1(P2_N387), .IN2(P2_N5495), .QN(n3806) );
  NAND2X0 U5417 ( .IN1(n3811), .IN2(n3812), .QN(P2_N1181) );
  NAND2X0 U5418 ( .IN1(P2_N998), .IN2(n3796), .QN(n3812) );
  NOR2X0 U5419 ( .QN(P2_N998), .IN1(n7015), .IN2(n7315) );
  NAND2X0 U5421 ( .IN1(n3813), .IN2(n3814), .QN(n2199) );
  NAND2X0 U5422 ( .IN1(N61), .IN2(n6739), .QN(n3814) );
  NAND2X0 U5423 ( .IN1(n9959), .IN2(N5), .QN(n3813) );
  NAND2X0 U5424 ( .IN1(P2_N386), .IN2(P2_N5495), .QN(n3811) );
  NAND2X0 U5425 ( .IN1(n3815), .IN2(n3816), .QN(P2_N1180) );
  NAND2X0 U5426 ( .IN1(P2_N997), .IN2(n3796), .QN(n3816) );
  NOR2X0 U5427 ( .QN(P2_N997), .IN1(n7013), .IN2(n7313) );
  NAND2X0 U5429 ( .IN1(n3817), .IN2(n3818), .QN(n2202) );
  NAND2X0 U5430 ( .IN1(N60), .IN2(n6739), .QN(n3818) );
  NAND2X0 U5431 ( .IN1(n9963), .IN2(N5), .QN(n3817) );
  NAND2X0 U5432 ( .IN1(P2_N385), .IN2(P2_N5495), .QN(n3815) );
  NAND2X0 U5433 ( .IN1(n3819), .IN2(n3820), .QN(P2_N1179) );
  NAND2X0 U5434 ( .IN1(P2_N996), .IN2(n3796), .QN(n3820) );
  NOR2X0 U5435 ( .QN(P2_N996), .IN1(n7013), .IN2(n7311) );
  NAND2X0 U5437 ( .IN1(n3821), .IN2(n3822), .QN(n2205) );
  NAND2X0 U5438 ( .IN1(N59), .IN2(n6739), .QN(n3822) );
  NAND2X0 U5439 ( .IN1(n9967), .IN2(N5), .QN(n3821) );
  NAND2X0 U5440 ( .IN1(P2_N384), .IN2(P2_N5495), .QN(n3819) );
  NAND2X0 U5441 ( .IN1(n3823), .IN2(n3824), .QN(P2_N1178) );
  NAND2X0 U5442 ( .IN1(n3796), .IN2(P2_N995), .QN(n3824) );
  NAND2X0 U5443 ( .IN1(n2006), .IN2(n3825), .QN(P2_N995) );
  NAND2X0 U5444 ( .IN1(P2_N914), .IN2(n2008), .QN(n3825) );
  NAND2X0 U5446 ( .IN1(N58), .IN2(n6737), .QN(n3827) );
  NAND2X0 U5447 ( .IN1(n9971), .IN2(n6736), .QN(n3826) );
  NAND2X0 U5448 ( .IN1(P2_N344), .IN2(n2693), .QN(n2006) );
  NAND2X0 U5449 ( .IN1(P2_N383), .IN2(P2_N5495), .QN(n3823) );
  NAND2X0 U5450 ( .IN1(n3828), .IN2(n3829), .QN(P2_N1177) );
  NAND2X0 U5451 ( .IN1(n3796), .IN2(P2_N994), .QN(n3829) );
  NAND2X0 U5452 ( .IN1(n2009), .IN2(n3830), .QN(P2_N994) );
  NAND2X0 U5453 ( .IN1(P2_N914), .IN2(n2011), .QN(n3830) );
  NAND2X0 U5455 ( .IN1(N57), .IN2(n6737), .QN(n3832) );
  NAND2X0 U5456 ( .IN1(n9975), .IN2(n6736), .QN(n3831) );
  NAND2X0 U5457 ( .IN1(P2_N345), .IN2(n2693), .QN(n2009) );
  NAND2X0 U5458 ( .IN1(P2_N382), .IN2(P2_N5495), .QN(n3828) );
  NAND2X0 U5459 ( .IN1(n3833), .IN2(n3834), .QN(P2_N1176) );
  NAND2X0 U5460 ( .IN1(n3796), .IN2(P2_N993), .QN(n3834) );
  NAND2X0 U5461 ( .IN1(n2012), .IN2(n3835), .QN(P2_N993) );
  NAND2X0 U5462 ( .IN1(P2_N914), .IN2(n2014), .QN(n3835) );
  NAND2X0 U5464 ( .IN1(N56), .IN2(n6737), .QN(n3837) );
  NAND2X0 U5465 ( .IN1(n9979), .IN2(n6736), .QN(n3836) );
  NAND2X0 U5466 ( .IN1(P2_N346), .IN2(n2693), .QN(n2012) );
  NAND2X0 U5467 ( .IN1(P2_N381), .IN2(P2_N5495), .QN(n3833) );
  NAND2X0 U5468 ( .IN1(n3838), .IN2(n3839), .QN(P2_N1175) );
  NAND2X0 U5469 ( .IN1(n3796), .IN2(P2_N992), .QN(n3839) );
  NAND2X0 U5470 ( .IN1(n2015), .IN2(n3840), .QN(P2_N992) );
  NAND2X0 U5471 ( .IN1(P2_N914), .IN2(n2017), .QN(n3840) );
  NAND2X0 U5473 ( .IN1(N55), .IN2(n6737), .QN(n3842) );
  NAND2X0 U5474 ( .IN1(n9983), .IN2(n6736), .QN(n3841) );
  NAND2X0 U5475 ( .IN1(P2_N347), .IN2(n2693), .QN(n2015) );
  NAND2X0 U5476 ( .IN1(P2_N380), .IN2(P2_N5495), .QN(n3838) );
  NAND2X0 U5477 ( .IN1(n3843), .IN2(n3844), .QN(P2_N1174) );
  NAND2X0 U5478 ( .IN1(n3796), .IN2(P2_N991), .QN(n3844) );
  NAND2X0 U5479 ( .IN1(n2018), .IN2(n3845), .QN(P2_N991) );
  NAND2X0 U5480 ( .IN1(n7009), .IN2(n2020), .QN(n3845) );
  NAND2X0 U5287 ( .IN1(P2_N378), .IN2(P2_N5496), .QN(n3738) );
  NAND2X0 U5288 ( .IN1(n3740), .IN2(n3741), .QN(P2_N1427) );
  NAND2X0 U5289 ( .IN1(n3710), .IN2(P2_N1244), .QN(n3741) );
  NAND2X0 U5290 ( .IN1(P2_N377), .IN2(P2_N5496), .QN(n3740) );
  NAND2X0 U5291 ( .IN1(n3742), .IN2(n3743), .QN(P2_N1426) );
  NAND2X0 U5292 ( .IN1(n3710), .IN2(P2_N1243), .QN(n3743) );
  NAND2X0 U5293 ( .IN1(P2_N376), .IN2(P2_N5496), .QN(n3742) );
  NAND2X0 U5294 ( .IN1(n3744), .IN2(n3745), .QN(P2_N1425) );
  NAND2X0 U5295 ( .IN1(n3710), .IN2(P2_N1242), .QN(n3745) );
  NAND2X0 U5296 ( .IN1(P2_N375), .IN2(P2_N5496), .QN(n3744) );
  NAND2X0 U5297 ( .IN1(n3746), .IN2(n3747), .QN(P2_N1424) );
  NAND2X0 U5298 ( .IN1(n3710), .IN2(P2_N1241), .QN(n3747) );
  NAND2X0 U5299 ( .IN1(P2_N374), .IN2(P2_N5496), .QN(n3746) );
  NAND2X0 U5300 ( .IN1(n3748), .IN2(n3749), .QN(P2_N1423) );
  NAND2X0 U5301 ( .IN1(n3710), .IN2(P2_N1240), .QN(n3749) );
  NAND2X0 U5302 ( .IN1(P2_N373), .IN2(P2_N5496), .QN(n3748) );
  NAND2X0 U5303 ( .IN1(n3750), .IN2(n3751), .QN(P2_N1422) );
  NAND2X0 U5304 ( .IN1(n3710), .IN2(P2_N1239), .QN(n3751) );
  NAND2X0 U5305 ( .IN1(P2_N372), .IN2(P2_N5496), .QN(n3750) );
  NAND2X0 U5306 ( .IN1(n3752), .IN2(n3753), .QN(P2_N1421) );
  NAND2X0 U5307 ( .IN1(n3710), .IN2(P2_N1238), .QN(n3753) );
  NAND2X0 U5308 ( .IN1(P2_N371), .IN2(P2_N5496), .QN(n3752) );
  NAND2X0 U5309 ( .IN1(n3754), .IN2(n3755), .QN(P2_N1420) );
  NAND2X0 U5310 ( .IN1(n3710), .IN2(P2_N1237), .QN(n3755) );
  NAND2X0 U5311 ( .IN1(P2_N370), .IN2(P2_N5496), .QN(n3754) );
  NAND2X0 U5312 ( .IN1(n3756), .IN2(n3757), .QN(P2_N1419) );
  NAND2X0 U5313 ( .IN1(n3710), .IN2(P2_N1236), .QN(n3757) );
  NAND2X0 U5314 ( .IN1(P2_N369), .IN2(P2_N5496), .QN(n3756) );
  NAND2X0 U5315 ( .IN1(n3758), .IN2(n3759), .QN(P2_N1418) );
  NAND2X0 U5316 ( .IN1(n3710), .IN2(P2_N1235), .QN(n3759) );
  NAND2X0 U5317 ( .IN1(P2_N368), .IN2(P2_N5496), .QN(n3758) );
  NAND2X0 U5318 ( .IN1(n3760), .IN2(n3761), .QN(P2_N1417) );
  NAND2X0 U5319 ( .IN1(n3710), .IN2(P2_N1234), .QN(n3761) );
  NAND2X0 U5320 ( .IN1(n18813), .IN2(P2_N5496), .QN(n3760) );
  NAND2X0 U5321 ( .IN1(n3762), .IN2(n3763), .QN(P2_N1416) );
  NAND2X0 U5322 ( .IN1(n3710), .IN2(P2_N1233), .QN(n3763) );
  NAND2X0 U5323 ( .IN1(n6683), .IN2(P2_N5496), .QN(n3762) );
  NAND2X0 U5324 ( .IN1(n3764), .IN2(n3765), .QN(P2_N1415) );
  NAND2X0 U5325 ( .IN1(n3710), .IN2(P2_N1232), .QN(n3765) );
  NAND2X0 U5326 ( .IN1(n6682), .IN2(P2_N5496), .QN(n3764) );
  NAND2X0 U5327 ( .IN1(n3766), .IN2(n3767), .QN(P2_N1414) );
  NAND2X0 U5328 ( .IN1(n3710), .IN2(P2_N1231), .QN(n3767) );
  NAND2X0 U5331 ( .IN1(n6681), .IN2(P2_N5496), .QN(n3766) );
  NAND2X0 U5336 ( .IN1(n7380), .IN2(n3770), .QN(P2_N1381) );
  NAND2X0 U5337 ( .IN1(n7379), .IN2(n3771), .QN(P2_N1379) );
  NOR2X0 U5338 ( .QN(P2_N1443), .IN1(n3771), .IN2(n3770) );
  INVX0 U5339 ( .ZN(n3770), .INP(n7379) );
  INVX0 U5340 ( .ZN(n3771), .INP(n7380) );
  NOR2X0 U5341 ( .QN(P2_N1260), .IN1(n7329), .IN2(n7007) );
  NOR2X0 U5342 ( .QN(P2_N1259), .IN1(n7013), .IN2(n7327) );
  NOR2X0 U5343 ( .QN(P2_N1258), .IN1(n7015), .IN2(n7325) );
  NOR2X0 U5344 ( .QN(P2_N1257), .IN1(n7015), .IN2(n7323) );
  NOR2X0 U5345 ( .QN(P2_N1256), .IN1(n7015), .IN2(n7321) );
  NOR2X0 U5346 ( .QN(P2_N1255), .IN1(n7015), .IN2(n7319) );
  NOR2X0 U5347 ( .QN(P2_N1254), .IN1(n7015), .IN2(n7317) );
  NOR2X0 U5348 ( .QN(P2_N1253), .IN1(n7015), .IN2(n7315) );
  NOR2X0 U5349 ( .QN(P2_N1252), .IN1(n7013), .IN2(n7313) );
  NOR2X0 U5350 ( .QN(P2_N1251), .IN1(n7013), .IN2(n7311) );
  NAND2X0 U5352 ( .IN1(n2006), .IN2(n3773), .QN(P2_N1250) );
  NAND2X0 U5353 ( .IN1(P2_N914), .IN2(n2008), .QN(n3773) );
  NAND2X0 U5354 ( .IN1(n2009), .IN2(n3774), .QN(P2_N1249) );
  NAND2X0 U5355 ( .IN1(P2_N914), .IN2(n2011), .QN(n3774) );
  NAND2X0 U5356 ( .IN1(n2012), .IN2(n3775), .QN(P2_N1248) );
  NAND2X0 U5357 ( .IN1(P2_N914), .IN2(n2014), .QN(n3775) );
  NAND2X0 U5358 ( .IN1(n2015), .IN2(n3776), .QN(P2_N1247) );
  NAND2X0 U5359 ( .IN1(P2_N914), .IN2(n2017), .QN(n3776) );
  NAND2X0 U5360 ( .IN1(n2018), .IN2(n3777), .QN(P2_N1246) );
  NAND2X0 U5361 ( .IN1(n7009), .IN2(n2020), .QN(n3777) );
  NAND2X0 U5362 ( .IN1(n2021), .IN2(n3778), .QN(P2_N1245) );
  NAND2X0 U5363 ( .IN1(n7009), .IN2(n2023), .QN(n3778) );
  NAND2X0 U5364 ( .IN1(n2024), .IN2(n3779), .QN(P2_N1244) );
  NAND2X0 U5365 ( .IN1(n7009), .IN2(n2026), .QN(n3779) );
  NAND2X0 U5366 ( .IN1(n2027), .IN2(n3780), .QN(P2_N1243) );
  NAND2X0 U5367 ( .IN1(n7010), .IN2(n2029), .QN(n3780) );
  NAND2X0 U5368 ( .IN1(n2030), .IN2(n3781), .QN(P2_N1242) );
  NAND2X0 U5369 ( .IN1(n7010), .IN2(n2032), .QN(n3781) );
  NAND2X0 U5370 ( .IN1(n2033), .IN2(n3782), .QN(P2_N1241) );
  NAND2X0 U5371 ( .IN1(n7010), .IN2(n2035), .QN(n3782) );
  NAND2X0 U5372 ( .IN1(n2036), .IN2(n3783), .QN(P2_N1240) );
  NAND2X0 U5373 ( .IN1(n7010), .IN2(n2038), .QN(n3783) );
  NAND2X0 U5374 ( .IN1(n2039), .IN2(n3784), .QN(P2_N1239) );
  NAND2X0 U5375 ( .IN1(n7010), .IN2(n2041), .QN(n3784) );
  NAND2X0 U5376 ( .IN1(n2042), .IN2(n3785), .QN(P2_N1238) );
  NAND2X0 U5377 ( .IN1(n7010), .IN2(n2044), .QN(n3785) );
  NAND2X0 U5378 ( .IN1(n2045), .IN2(n3786), .QN(P2_N1237) );
  NAND2X0 U5379 ( .IN1(n7006), .IN2(n2047), .QN(n3786) );
  NAND2X0 U5380 ( .IN1(n2048), .IN2(n3787), .QN(P2_N1236) );
  NAND2X0 U5381 ( .IN1(n7006), .IN2(n2050), .QN(n3787) );
  NAND2X0 U5382 ( .IN1(n2051), .IN2(n3788), .QN(P2_N1235) );
  NAND2X0 U5383 ( .IN1(n7006), .IN2(n2053), .QN(n3788) );
  NAND2X0 U5384 ( .IN1(n2054), .IN2(n3789), .QN(P2_N1234) );
  NAND2X0 U5385 ( .IN1(n7462), .IN2(n2056), .QN(n3789) );
  NOR2X0 U5191 ( .QN(P2_N1514), .IN1(n7327), .IN2(n7007) );
  NOR2X0 U5192 ( .QN(P2_N1513), .IN1(n7325), .IN2(n7007) );
  NOR2X0 U5193 ( .QN(P2_N1512), .IN1(n7323), .IN2(n7011) );
  NOR2X0 U5194 ( .QN(P2_N1511), .IN1(n7321), .IN2(n7011) );
  NOR2X0 U5195 ( .QN(P2_N1510), .IN1(n7319), .IN2(n7011) );
  NOR2X0 U5196 ( .QN(P2_N1509), .IN1(n7317), .IN2(n7011) );
  NOR2X0 U5197 ( .QN(P2_N1508), .IN1(n7315), .IN2(n7015) );
  NOR2X0 U5198 ( .QN(P2_N1507), .IN1(n7313), .IN2(n7015) );
  NOR2X0 U5199 ( .QN(P2_N1506), .IN1(n7311), .IN2(n7015) );
  NAND2X0 U5201 ( .IN1(n2006), .IN2(n3687), .QN(P2_N1505) );
  NAND2X0 U5202 ( .IN1(P2_N914), .IN2(n2008), .QN(n3687) );
  NAND2X0 U5203 ( .IN1(n2009), .IN2(n3688), .QN(P2_N1504) );
  NAND2X0 U5204 ( .IN1(P2_N914), .IN2(n2011), .QN(n3688) );
  NAND2X0 U5205 ( .IN1(n2012), .IN2(n3689), .QN(P2_N1503) );
  NAND2X0 U5206 ( .IN1(n7012), .IN2(n2014), .QN(n3689) );
  NAND2X0 U5207 ( .IN1(n2015), .IN2(n3690), .QN(P2_N1502) );
  NAND2X0 U5208 ( .IN1(P2_N914), .IN2(n2017), .QN(n3690) );
  NAND2X0 U5209 ( .IN1(n2018), .IN2(n3691), .QN(P2_N1501) );
  NAND2X0 U5210 ( .IN1(n7009), .IN2(n2020), .QN(n3691) );
  NAND2X0 U5211 ( .IN1(n2021), .IN2(n3692), .QN(P2_N1500) );
  NAND2X0 U5212 ( .IN1(n7009), .IN2(n2023), .QN(n3692) );
  NAND2X0 U5213 ( .IN1(n2024), .IN2(n3693), .QN(P2_N1499) );
  NAND2X0 U5214 ( .IN1(n7009), .IN2(n2026), .QN(n3693) );
  NAND2X0 U5215 ( .IN1(n2027), .IN2(n3694), .QN(P2_N1498) );
  NAND2X0 U5216 ( .IN1(n7009), .IN2(n2029), .QN(n3694) );
  NAND2X0 U5217 ( .IN1(n2030), .IN2(n3695), .QN(P2_N1497) );
  NAND2X0 U5218 ( .IN1(n7010), .IN2(n2032), .QN(n3695) );
  NAND2X0 U5219 ( .IN1(n2033), .IN2(n3696), .QN(P2_N1496) );
  NAND2X0 U5220 ( .IN1(n7010), .IN2(n2035), .QN(n3696) );
  NAND2X0 U5221 ( .IN1(n2036), .IN2(n3697), .QN(P2_N1495) );
  NAND2X0 U5222 ( .IN1(n7016), .IN2(n2038), .QN(n3697) );
  NAND2X0 U5223 ( .IN1(n2039), .IN2(n3698), .QN(P2_N1494) );
  NAND2X0 U5224 ( .IN1(n7016), .IN2(n2041), .QN(n3698) );
  NAND2X0 U5225 ( .IN1(n2042), .IN2(n3699), .QN(P2_N1493) );
  NAND2X0 U5226 ( .IN1(n7016), .IN2(n2044), .QN(n3699) );
  NAND2X0 U5227 ( .IN1(n2045), .IN2(n3700), .QN(P2_N1492) );
  NAND2X0 U5228 ( .IN1(n7016), .IN2(n2047), .QN(n3700) );
  NAND2X0 U5229 ( .IN1(n2048), .IN2(n3701), .QN(P2_N1491) );
  NAND2X0 U5230 ( .IN1(n7016), .IN2(n2050), .QN(n3701) );
  NAND2X0 U5231 ( .IN1(n2051), .IN2(n3702), .QN(P2_N1490) );
  NAND2X0 U5232 ( .IN1(n7006), .IN2(n2053), .QN(n3702) );
  NAND2X0 U5233 ( .IN1(n2054), .IN2(n3703), .QN(P2_N1489) );
  NAND2X0 U5234 ( .IN1(n7006), .IN2(n2056), .QN(n3703) );
  NAND2X0 U5235 ( .IN1(n2057), .IN2(n3704), .QN(P2_N1488) );
  NAND2X0 U5236 ( .IN1(n7006), .IN2(n2059), .QN(n3704) );
  NAND2X0 U5237 ( .IN1(n2060), .IN2(n3705), .QN(P2_N1487) );
  NAND2X0 U5238 ( .IN1(n7006), .IN2(n2062), .QN(n3705) );
  NAND2X0 U5239 ( .IN1(n2063), .IN2(n3706), .QN(P2_N1486) );
  NAND2X0 U5240 ( .IN1(n7006), .IN2(n2065), .QN(n3706) );
  NAND2X0 U5243 ( .IN1(n3708), .IN2(n3709), .QN(P2_N1442) );
  NAND2X0 U5244 ( .IN1(P2_N1259), .IN2(n3710), .QN(n3709) );
  NAND2X0 U5245 ( .IN1(P2_N392), .IN2(P2_N5496), .QN(n3708) );
  NAND2X0 U5246 ( .IN1(n3712), .IN2(n3713), .QN(P2_N1441) );
  NAND2X0 U5247 ( .IN1(P2_N1258), .IN2(n3710), .QN(n3713) );
  NAND2X0 U5248 ( .IN1(P2_N391), .IN2(P2_N5496), .QN(n3712) );
  NAND2X0 U5249 ( .IN1(n3714), .IN2(n3715), .QN(P2_N1440) );
  NAND2X0 U5250 ( .IN1(P2_N1257), .IN2(n3710), .QN(n3715) );
  NAND2X0 U5251 ( .IN1(P2_N390), .IN2(P2_N5496), .QN(n3714) );
  NAND2X0 U5252 ( .IN1(n3716), .IN2(n3717), .QN(P2_N1439) );
  NAND2X0 U5253 ( .IN1(P2_N1256), .IN2(n3710), .QN(n3717) );
  NAND2X0 U5254 ( .IN1(P2_N389), .IN2(P2_N5496), .QN(n3716) );
  NAND2X0 U5255 ( .IN1(n3718), .IN2(n3719), .QN(P2_N1438) );
  NAND2X0 U5256 ( .IN1(P2_N1255), .IN2(n3710), .QN(n3719) );
  NAND2X0 U5257 ( .IN1(P2_N388), .IN2(P2_N5496), .QN(n3718) );
  NAND2X0 U5258 ( .IN1(n3720), .IN2(n3721), .QN(P2_N1437) );
  NAND2X0 U5259 ( .IN1(P2_N1254), .IN2(n3710), .QN(n3721) );
  NAND2X0 U5260 ( .IN1(P2_N387), .IN2(P2_N5496), .QN(n3720) );
  NAND2X0 U5261 ( .IN1(n3722), .IN2(n3723), .QN(P2_N1436) );
  NAND2X0 U5262 ( .IN1(P2_N1253), .IN2(n3710), .QN(n3723) );
  NAND2X0 U5263 ( .IN1(P2_N386), .IN2(P2_N5496), .QN(n3722) );
  NAND2X0 U5264 ( .IN1(n3724), .IN2(n3725), .QN(P2_N1435) );
  NAND2X0 U5265 ( .IN1(P2_N1252), .IN2(n3710), .QN(n3725) );
  NAND2X0 U5266 ( .IN1(P2_N385), .IN2(P2_N5496), .QN(n3724) );
  NAND2X0 U5267 ( .IN1(n3726), .IN2(n3727), .QN(P2_N1434) );
  NAND2X0 U5268 ( .IN1(P2_N1251), .IN2(n3710), .QN(n3727) );
  NAND2X0 U5269 ( .IN1(P2_N384), .IN2(P2_N5496), .QN(n3726) );
  NAND2X0 U5270 ( .IN1(n3728), .IN2(n3729), .QN(P2_N1433) );
  NAND2X0 U5271 ( .IN1(n3710), .IN2(P2_N1250), .QN(n3729) );
  NAND2X0 U5272 ( .IN1(P2_N383), .IN2(P2_N5496), .QN(n3728) );
  NAND2X0 U5273 ( .IN1(n3730), .IN2(n3731), .QN(P2_N1432) );
  NAND2X0 U5274 ( .IN1(n3710), .IN2(P2_N1249), .QN(n3731) );
  NAND2X0 U5275 ( .IN1(P2_N382), .IN2(P2_N5496), .QN(n3730) );
  NAND2X0 U5276 ( .IN1(n3732), .IN2(n3733), .QN(P2_N1431) );
  NAND2X0 U5277 ( .IN1(n3710), .IN2(P2_N1248), .QN(n3733) );
  NAND2X0 U5278 ( .IN1(P2_N381), .IN2(P2_N5496), .QN(n3732) );
  NAND2X0 U5279 ( .IN1(n3734), .IN2(n3735), .QN(P2_N1430) );
  NAND2X0 U5280 ( .IN1(n3710), .IN2(P2_N1247), .QN(n3735) );
  NAND2X0 U5281 ( .IN1(P2_N380), .IN2(P2_N5496), .QN(n3734) );
  NAND2X0 U5282 ( .IN1(n3736), .IN2(n3737), .QN(P2_N1429) );
  NAND2X0 U5283 ( .IN1(n3710), .IN2(P2_N1246), .QN(n3737) );
  NAND2X0 U5284 ( .IN1(P2_N379), .IN2(P2_N5496), .QN(n3736) );
  NAND2X0 U5285 ( .IN1(n3738), .IN2(n3739), .QN(P2_N1428) );
  NAND2X0 U5286 ( .IN1(n3710), .IN2(P2_N1245), .QN(n3739) );
  NAND2X0 U5093 ( .IN1(P2_N1756), .IN2(n3624), .QN(n3623) );
  NAND2X0 U5094 ( .IN1(P2_N392), .IN2(P2_N5502), .QN(n3622) );
  NAND2X0 U5095 ( .IN1(n3626), .IN2(n3627), .QN(P2_N1814) );
  NAND2X0 U5096 ( .IN1(P2_N1755), .IN2(n3624), .QN(n3627) );
  NAND2X0 U5097 ( .IN1(P2_N391), .IN2(P2_N5502), .QN(n3626) );
  NAND2X0 U5098 ( .IN1(n3628), .IN2(n3629), .QN(P2_N1813) );
  NAND2X0 U5099 ( .IN1(P2_N1754), .IN2(n3624), .QN(n3629) );
  NAND2X0 U5100 ( .IN1(P2_N390), .IN2(P2_N5502), .QN(n3628) );
  NAND2X0 U5101 ( .IN1(n3630), .IN2(n3631), .QN(P2_N1812) );
  NAND2X0 U5102 ( .IN1(P2_N1753), .IN2(n3624), .QN(n3631) );
  NAND2X0 U5103 ( .IN1(P2_N389), .IN2(P2_N5502), .QN(n3630) );
  NAND2X0 U5104 ( .IN1(n3632), .IN2(n3633), .QN(P2_N1811) );
  NAND2X0 U5105 ( .IN1(P2_N1752), .IN2(n3624), .QN(n3633) );
  NAND2X0 U5106 ( .IN1(P2_N388), .IN2(P2_N5502), .QN(n3632) );
  NAND2X0 U5107 ( .IN1(n3634), .IN2(n3635), .QN(P2_N1810) );
  NAND2X0 U5108 ( .IN1(P2_N1751), .IN2(n3624), .QN(n3635) );
  NAND2X0 U5109 ( .IN1(P2_N387), .IN2(P2_N5502), .QN(n3634) );
  NAND2X0 U5110 ( .IN1(n3636), .IN2(n3637), .QN(P2_N1809) );
  NAND2X0 U5111 ( .IN1(P2_N1750), .IN2(n3624), .QN(n3637) );
  NAND2X0 U5112 ( .IN1(P2_N386), .IN2(P2_N5502), .QN(n3636) );
  NAND2X0 U5113 ( .IN1(n3638), .IN2(n3639), .QN(P2_N1808) );
  NAND2X0 U5114 ( .IN1(P2_N1749), .IN2(n3624), .QN(n3639) );
  NAND2X0 U5115 ( .IN1(P2_N385), .IN2(P2_N5502), .QN(n3638) );
  NAND2X0 U5116 ( .IN1(n3640), .IN2(n3641), .QN(P2_N1807) );
  NAND2X0 U5117 ( .IN1(P2_N1748), .IN2(n3624), .QN(n3641) );
  NAND2X0 U5118 ( .IN1(P2_N384), .IN2(P2_N5502), .QN(n3640) );
  NAND2X0 U5119 ( .IN1(n3642), .IN2(n3643), .QN(P2_N1806) );
  NAND2X0 U5120 ( .IN1(P2_N1747), .IN2(n3624), .QN(n3643) );
  NAND2X0 U5121 ( .IN1(P2_N383), .IN2(P2_N5502), .QN(n3642) );
  NAND2X0 U5122 ( .IN1(n3644), .IN2(n3645), .QN(P2_N1805) );
  NAND2X0 U5123 ( .IN1(P2_N1746), .IN2(n3624), .QN(n3645) );
  NAND2X0 U5124 ( .IN1(P2_N382), .IN2(P2_N5502), .QN(n3644) );
  NAND2X0 U5125 ( .IN1(n3646), .IN2(n3647), .QN(P2_N1804) );
  NAND2X0 U5126 ( .IN1(P2_N1745), .IN2(n3624), .QN(n3647) );
  NAND2X0 U5127 ( .IN1(P2_N381), .IN2(P2_N5502), .QN(n3646) );
  NAND2X0 U5128 ( .IN1(n3648), .IN2(n3649), .QN(P2_N1803) );
  NAND2X0 U5129 ( .IN1(P2_N1744), .IN2(n3624), .QN(n3649) );
  NAND2X0 U5130 ( .IN1(P2_N380), .IN2(P2_N5502), .QN(n3648) );
  NAND2X0 U5131 ( .IN1(n3650), .IN2(n3651), .QN(P2_N1802) );
  NAND2X0 U5132 ( .IN1(P2_N1743), .IN2(n3624), .QN(n3651) );
  NAND2X0 U5133 ( .IN1(P2_N379), .IN2(P2_N5502), .QN(n3650) );
  NAND2X0 U5134 ( .IN1(n3652), .IN2(n3653), .QN(P2_N1801) );
  NAND2X0 U5135 ( .IN1(P2_N1742), .IN2(n3624), .QN(n3653) );
  NAND2X0 U5136 ( .IN1(P2_N378), .IN2(P2_N5502), .QN(n3652) );
  NAND2X0 U5137 ( .IN1(n3654), .IN2(n3655), .QN(P2_N1800) );
  NAND2X0 U5138 ( .IN1(P2_N1741), .IN2(n3624), .QN(n3655) );
  NAND2X0 U5139 ( .IN1(P2_N377), .IN2(P2_N5502), .QN(n3654) );
  NAND2X0 U5140 ( .IN1(n3656), .IN2(n3657), .QN(P2_N1799) );
  NAND2X0 U5141 ( .IN1(P2_N1740), .IN2(n3624), .QN(n3657) );
  NAND2X0 U5142 ( .IN1(P2_N376), .IN2(P2_N5502), .QN(n3656) );
  NAND2X0 U5143 ( .IN1(n3658), .IN2(n3659), .QN(P2_N1798) );
  NAND2X0 U5144 ( .IN1(P2_N1739), .IN2(n3624), .QN(n3659) );
  NAND2X0 U5145 ( .IN1(P2_N375), .IN2(P2_N5502), .QN(n3658) );
  NAND2X0 U5146 ( .IN1(n3660), .IN2(n3661), .QN(P2_N1797) );
  NAND2X0 U5147 ( .IN1(P2_N1738), .IN2(n3624), .QN(n3661) );
  NAND2X0 U5148 ( .IN1(P2_N374), .IN2(P2_N5502), .QN(n3660) );
  NAND2X0 U5149 ( .IN1(n3662), .IN2(n3663), .QN(P2_N1796) );
  NAND2X0 U5150 ( .IN1(P2_N1737), .IN2(n3624), .QN(n3663) );
  NAND2X0 U5151 ( .IN1(P2_N373), .IN2(P2_N5502), .QN(n3662) );
  NAND2X0 U5152 ( .IN1(n3664), .IN2(n3665), .QN(P2_N1795) );
  NAND2X0 U5153 ( .IN1(P2_N1736), .IN2(n3624), .QN(n3665) );
  NAND2X0 U5154 ( .IN1(P2_N372), .IN2(P2_N5502), .QN(n3664) );
  NAND2X0 U5155 ( .IN1(n3666), .IN2(n3667), .QN(P2_N1794) );
  NAND2X0 U5156 ( .IN1(P2_N1735), .IN2(n3624), .QN(n3667) );
  NAND2X0 U5157 ( .IN1(P2_N371), .IN2(P2_N5502), .QN(n3666) );
  NAND2X0 U5158 ( .IN1(n3668), .IN2(n3669), .QN(P2_N1793) );
  NAND2X0 U5159 ( .IN1(P2_N1734), .IN2(n3624), .QN(n3669) );
  NAND2X0 U5160 ( .IN1(P2_N370), .IN2(P2_N5502), .QN(n3668) );
  NAND2X0 U5161 ( .IN1(n3670), .IN2(n3671), .QN(P2_N1792) );
  NAND2X0 U5162 ( .IN1(P2_N1733), .IN2(n3624), .QN(n3671) );
  NAND2X0 U5163 ( .IN1(P2_N369), .IN2(P2_N5502), .QN(n3670) );
  NAND2X0 U5164 ( .IN1(n3672), .IN2(n3673), .QN(P2_N1791) );
  NAND2X0 U5165 ( .IN1(P2_N1732), .IN2(n3624), .QN(n3673) );
  NAND2X0 U5166 ( .IN1(P2_N368), .IN2(P2_N5502), .QN(n3672) );
  NAND2X0 U5167 ( .IN1(n3674), .IN2(n3675), .QN(P2_N1790) );
  NAND2X0 U5168 ( .IN1(P2_N1731), .IN2(n3624), .QN(n3675) );
  NAND2X0 U5169 ( .IN1(n18813), .IN2(P2_N5502), .QN(n3674) );
  NAND2X0 U5170 ( .IN1(n3676), .IN2(n3677), .QN(P2_N1789) );
  NAND2X0 U5171 ( .IN1(P2_N1730), .IN2(n3624), .QN(n3677) );
  NAND2X0 U5172 ( .IN1(n6683), .IN2(P2_N5502), .QN(n3676) );
  NAND2X0 U5173 ( .IN1(n3678), .IN2(n3679), .QN(P2_N1788) );
  NAND2X0 U5174 ( .IN1(P2_N1729), .IN2(n3624), .QN(n3679) );
  NAND2X0 U5175 ( .IN1(n6682), .IN2(P2_N5502), .QN(n3678) );
  NAND2X0 U5176 ( .IN1(n3680), .IN2(n3681), .QN(P2_N1787) );
  NAND2X0 U5177 ( .IN1(P2_N1728), .IN2(n3624), .QN(n3681) );
  NAND2X0 U5180 ( .IN1(n6681), .IN2(P2_N5502), .QN(n3680) );
  NAND2X0 U5185 ( .IN1(n7382), .IN2(n3684), .QN(P2_N1635) );
  NAND2X0 U5186 ( .IN1(n7381), .IN2(n3685), .QN(P2_N1633) );
  NOR2X0 U5187 ( .QN(P2_N1816), .IN1(n3685), .IN2(n3684) );
  INVX0 U5188 ( .ZN(n3684), .INP(n7381) );
  INVX0 U5189 ( .ZN(n3685), .INP(n7382) );
  NOR2X0 U5190 ( .QN(P2_N1515), .IN1(n7329), .IN2(n7007) );
  NAND2X0 U4992 ( .IN1(n3564), .IN2(n3565), .QN(P2_N2162) );
  NAND2X0 U4993 ( .IN1(P2_N2103), .IN2(n3512), .QN(n3565) );
  NAND2X0 U4994 ( .IN1(n6683), .IN2(P2_N5503), .QN(n3564) );
  NAND2X0 U4995 ( .IN1(n3566), .IN2(n3567), .QN(P2_N2161) );
  NAND2X0 U4996 ( .IN1(P2_N2102), .IN2(n3512), .QN(n3567) );
  NAND2X0 U4997 ( .IN1(n6682), .IN2(P2_N5503), .QN(n3566) );
  NAND2X0 U4998 ( .IN1(n3568), .IN2(n3569), .QN(P2_N2160) );
  NAND2X0 U4999 ( .IN1(P2_N2101), .IN2(n3512), .QN(n3569) );
  NAND2X0 U5002 ( .IN1(n6681), .IN2(P2_N5503), .QN(n3568) );
  NAND2X0 U5007 ( .IN1(n7384), .IN2(n3572), .QN(P2_N2008) );
  NAND2X0 U5008 ( .IN1(n7383), .IN2(n3573), .QN(P2_N2006) );
  NOR2X0 U5009 ( .QN(P2_N2189), .IN1(n3573), .IN2(n3572) );
  INVX0 U5010 ( .ZN(n3572), .INP(n7383) );
  INVX0 U5011 ( .ZN(n3573), .INP(n7384) );
  AND2X1 U5012 ( .IN1(P2_N134), .IN2(n3574), .Q(P2_N190) );
  NAND2X0 U5013 ( .IN1(n3575), .IN2(n3576), .QN(n3574) );
  NOR2X0 U5014 ( .QN(n3576), .IN1(n3577), .IN2(n3578) );
  NAND2X0 U5015 ( .IN1(n3579), .IN2(n3580), .QN(n3578) );
  AND2X1 U5016 ( .IN1(n3581), .IN2(n3582), .Q(n3580) );
  NOR2X0 U5017 ( .QN(n3582), .IN1(P2_N156), .IN2(P2_N155) );
  NOR2X0 U5018 ( .QN(n3581), .IN1(P2_N154), .IN2(P2_N153) );
  NOR2X0 U5019 ( .QN(n3579), .IN1(P2_N150), .IN2(n3583) );
  OR2X1 U5020 ( .IN2(P2_N151), .IN1(P2_N152), .Q(n3583) );
  NAND2X0 U5021 ( .IN1(n3584), .IN2(n3585), .QN(n3577) );
  AND2X1 U5022 ( .IN1(n3586), .IN2(n3587), .Q(n3585) );
  NOR2X0 U5023 ( .QN(n3587), .IN1(P2_N163), .IN2(P2_N162) );
  NOR2X0 U5024 ( .QN(n3586), .IN1(P2_N161), .IN2(P2_N160) );
  NOR2X0 U5025 ( .QN(n3584), .IN1(P2_N157), .IN2(n3588) );
  OR2X1 U5026 ( .IN2(P2_N158), .IN1(P2_N159), .Q(n3588) );
  NOR2X0 U5027 ( .QN(n3575), .IN1(n3589), .IN2(n3590) );
  NAND2X0 U5028 ( .IN1(n3591), .IN2(n3592), .QN(n3590) );
  NOR2X0 U5029 ( .QN(n3592), .IN1(P2_N140), .IN2(n3593) );
  OR2X1 U5030 ( .IN2(P2_N141), .IN1(P2_N142), .Q(n3593) );
  NOR2X0 U5031 ( .QN(n3591), .IN1(P2_N137), .IN2(n3594) );
  OR2X1 U5032 ( .IN2(P2_N138), .IN1(P2_N139), .Q(n3594) );
  NAND2X0 U5033 ( .IN1(n3595), .IN2(n3596), .QN(n3589) );
  AND2X1 U5034 ( .IN1(n3597), .IN2(n3598), .Q(n3596) );
  NOR2X0 U5035 ( .QN(n3598), .IN1(P2_N149), .IN2(P2_N148) );
  NOR2X0 U5036 ( .QN(n3597), .IN1(P2_N147), .IN2(P2_N146) );
  NOR2X0 U5037 ( .QN(n3595), .IN1(P2_N143), .IN2(n3599) );
  OR2X1 U5038 ( .IN2(P2_N144), .IN1(P2_N145), .Q(n3599) );
  NOR2X0 U5039 ( .QN(P2_N1888), .IN1(n7329), .IN2(n7007) );
  NOR2X0 U5040 ( .QN(P2_N1887), .IN1(n7327), .IN2(n7007) );
  NOR2X0 U5041 ( .QN(P2_N1886), .IN1(n7325), .IN2(n7007) );
  NOR2X0 U5042 ( .QN(P2_N1885), .IN1(n7323), .IN2(n7011) );
  NOR2X0 U5043 ( .QN(P2_N1884), .IN1(n7321), .IN2(n7011) );
  NOR2X0 U5044 ( .QN(P2_N1883), .IN1(n7319), .IN2(n7011) );
  NOR2X0 U5045 ( .QN(P2_N1882), .IN1(n7317), .IN2(n7011) );
  NOR2X0 U5046 ( .QN(P2_N1881), .IN1(n7315), .IN2(n7015) );
  NOR2X0 U5047 ( .QN(P2_N1880), .IN1(n7313), .IN2(n7015) );
  NOR2X0 U5048 ( .QN(P2_N1879), .IN1(n7311), .IN2(n7011) );
  NAND2X0 U5050 ( .IN1(n2006), .IN2(n3601), .QN(P2_N1878) );
  NAND2X0 U5051 ( .IN1(n7012), .IN2(n2008), .QN(n3601) );
  NAND2X0 U5052 ( .IN1(n2009), .IN2(n3602), .QN(P2_N1877) );
  NAND2X0 U5053 ( .IN1(n7012), .IN2(n2011), .QN(n3602) );
  NAND2X0 U5054 ( .IN1(n2012), .IN2(n3603), .QN(P2_N1876) );
  NAND2X0 U5055 ( .IN1(P2_N914), .IN2(n2014), .QN(n3603) );
  NAND2X0 U5056 ( .IN1(n2015), .IN2(n3604), .QN(P2_N1875) );
  NAND2X0 U5057 ( .IN1(P2_N914), .IN2(n2017), .QN(n3604) );
  NAND2X0 U5058 ( .IN1(n2018), .IN2(n3605), .QN(P2_N1874) );
  NAND2X0 U5059 ( .IN1(n7009), .IN2(n2020), .QN(n3605) );
  NAND2X0 U5060 ( .IN1(n2021), .IN2(n3606), .QN(P2_N1873) );
  NAND2X0 U5061 ( .IN1(n7009), .IN2(n2023), .QN(n3606) );
  NAND2X0 U5062 ( .IN1(n2024), .IN2(n3607), .QN(P2_N1872) );
  NAND2X0 U5063 ( .IN1(n7009), .IN2(n2026), .QN(n3607) );
  NAND2X0 U5064 ( .IN1(n2027), .IN2(n3608), .QN(P2_N1871) );
  NAND2X0 U5065 ( .IN1(n7009), .IN2(n2029), .QN(n3608) );
  NAND2X0 U5066 ( .IN1(n2030), .IN2(n3609), .QN(P2_N1870) );
  NAND2X0 U5067 ( .IN1(n7010), .IN2(n2032), .QN(n3609) );
  NAND2X0 U5068 ( .IN1(n2033), .IN2(n3610), .QN(P2_N1869) );
  NAND2X0 U5069 ( .IN1(n7010), .IN2(n2035), .QN(n3610) );
  NAND2X0 U5070 ( .IN1(n2036), .IN2(n3611), .QN(P2_N1868) );
  NAND2X0 U5071 ( .IN1(n7016), .IN2(n2038), .QN(n3611) );
  NAND2X0 U5072 ( .IN1(n2039), .IN2(n3612), .QN(P2_N1867) );
  NAND2X0 U5073 ( .IN1(n7016), .IN2(n2041), .QN(n3612) );
  NAND2X0 U5074 ( .IN1(n2042), .IN2(n3613), .QN(P2_N1866) );
  NAND2X0 U5075 ( .IN1(n7016), .IN2(n2044), .QN(n3613) );
  NAND2X0 U5076 ( .IN1(n2045), .IN2(n3614), .QN(P2_N1865) );
  NAND2X0 U5077 ( .IN1(n7016), .IN2(n2047), .QN(n3614) );
  NAND2X0 U5078 ( .IN1(n2048), .IN2(n3615), .QN(P2_N1864) );
  NAND2X0 U5079 ( .IN1(n7006), .IN2(n2050), .QN(n3615) );
  NAND2X0 U5080 ( .IN1(n2051), .IN2(n3616), .QN(P2_N1863) );
  NAND2X0 U5081 ( .IN1(n7006), .IN2(n2053), .QN(n3616) );
  NAND2X0 U5082 ( .IN1(n2054), .IN2(n3617), .QN(P2_N1862) );
  NAND2X0 U5083 ( .IN1(n7006), .IN2(n2056), .QN(n3617) );
  NAND2X0 U5084 ( .IN1(n2057), .IN2(n3618), .QN(P2_N1861) );
  NAND2X0 U5085 ( .IN1(n7462), .IN2(n2059), .QN(n3618) );
  NAND2X0 U5086 ( .IN1(n2060), .IN2(n3619), .QN(P2_N1860) );
  NAND2X0 U5087 ( .IN1(n7462), .IN2(n2062), .QN(n3619) );
  NAND2X0 U5088 ( .IN1(n2063), .IN2(n3620), .QN(P2_N1859) );
  NAND2X0 U5089 ( .IN1(n7462), .IN2(n2065), .QN(n3620) );
  NAND2X0 U5092 ( .IN1(n3622), .IN2(n3623), .QN(P2_N1815) );
  NAND2X0 U4897 ( .IN1(n7016), .IN2(n2044), .QN(n3501) );
  NAND2X0 U4898 ( .IN1(n2045), .IN2(n3502), .QN(P2_N2238) );
  NAND2X0 U4899 ( .IN1(n7016), .IN2(n2047), .QN(n3502) );
  NAND2X0 U4900 ( .IN1(n2048), .IN2(n3503), .QN(P2_N2237) );
  NAND2X0 U4901 ( .IN1(n7016), .IN2(n2050), .QN(n3503) );
  NAND2X0 U4902 ( .IN1(n2051), .IN2(n3504), .QN(P2_N2236) );
  NAND2X0 U4903 ( .IN1(n7006), .IN2(n2053), .QN(n3504) );
  NAND2X0 U4904 ( .IN1(n2054), .IN2(n3505), .QN(P2_N2235) );
  NAND2X0 U4905 ( .IN1(n7006), .IN2(n2056), .QN(n3505) );
  NAND2X0 U4906 ( .IN1(n2057), .IN2(n3506), .QN(P2_N2234) );
  NAND2X0 U4907 ( .IN1(n7006), .IN2(n2059), .QN(n3506) );
  NAND2X0 U4908 ( .IN1(n2060), .IN2(n3507), .QN(P2_N2233) );
  NAND2X0 U4909 ( .IN1(n7006), .IN2(n2062), .QN(n3507) );
  NAND2X0 U4910 ( .IN1(n2063), .IN2(n3508), .QN(P2_N2232) );
  NAND2X0 U4911 ( .IN1(n7006), .IN2(n2065), .QN(n3508) );
  NAND2X0 U4914 ( .IN1(n3510), .IN2(n3511), .QN(P2_N2188) );
  NAND2X0 U4915 ( .IN1(P2_N2129), .IN2(n3512), .QN(n3511) );
  NAND2X0 U4916 ( .IN1(P2_N392), .IN2(P2_N5503), .QN(n3510) );
  NAND2X0 U4917 ( .IN1(n3514), .IN2(n3515), .QN(P2_N2187) );
  NAND2X0 U4918 ( .IN1(P2_N2128), .IN2(n3512), .QN(n3515) );
  NAND2X0 U4919 ( .IN1(P2_N391), .IN2(P2_N5503), .QN(n3514) );
  NAND2X0 U4920 ( .IN1(n3516), .IN2(n3517), .QN(P2_N2186) );
  NAND2X0 U4921 ( .IN1(P2_N2127), .IN2(n3512), .QN(n3517) );
  NAND2X0 U4922 ( .IN1(P2_N390), .IN2(P2_N5503), .QN(n3516) );
  NAND2X0 U4923 ( .IN1(n3518), .IN2(n3519), .QN(P2_N2185) );
  NAND2X0 U4924 ( .IN1(P2_N2126), .IN2(n3512), .QN(n3519) );
  NAND2X0 U4925 ( .IN1(P2_N389), .IN2(P2_N5503), .QN(n3518) );
  NAND2X0 U4926 ( .IN1(n3520), .IN2(n3521), .QN(P2_N2184) );
  NAND2X0 U4927 ( .IN1(P2_N2125), .IN2(n3512), .QN(n3521) );
  NAND2X0 U4928 ( .IN1(P2_N388), .IN2(P2_N5503), .QN(n3520) );
  NAND2X0 U4929 ( .IN1(n3522), .IN2(n3523), .QN(P2_N2183) );
  NAND2X0 U4930 ( .IN1(P2_N2124), .IN2(n3512), .QN(n3523) );
  NAND2X0 U4931 ( .IN1(P2_N387), .IN2(P2_N5503), .QN(n3522) );
  NAND2X0 U4932 ( .IN1(n3524), .IN2(n3525), .QN(P2_N2182) );
  NAND2X0 U4933 ( .IN1(P2_N2123), .IN2(n3512), .QN(n3525) );
  NAND2X0 U4934 ( .IN1(P2_N386), .IN2(P2_N5503), .QN(n3524) );
  NAND2X0 U4935 ( .IN1(n3526), .IN2(n3527), .QN(P2_N2181) );
  NAND2X0 U4936 ( .IN1(P2_N2122), .IN2(n3512), .QN(n3527) );
  NAND2X0 U4937 ( .IN1(P2_N385), .IN2(P2_N5503), .QN(n3526) );
  NAND2X0 U4938 ( .IN1(n3528), .IN2(n3529), .QN(P2_N2180) );
  NAND2X0 U4939 ( .IN1(P2_N2121), .IN2(n3512), .QN(n3529) );
  NAND2X0 U4940 ( .IN1(P2_N384), .IN2(P2_N5503), .QN(n3528) );
  NAND2X0 U4941 ( .IN1(n3530), .IN2(n3531), .QN(P2_N2179) );
  NAND2X0 U4942 ( .IN1(P2_N2120), .IN2(n3512), .QN(n3531) );
  NAND2X0 U4943 ( .IN1(P2_N383), .IN2(P2_N5503), .QN(n3530) );
  NAND2X0 U4944 ( .IN1(n3532), .IN2(n3533), .QN(P2_N2178) );
  NAND2X0 U4945 ( .IN1(P2_N2119), .IN2(n3512), .QN(n3533) );
  NAND2X0 U4946 ( .IN1(P2_N382), .IN2(P2_N5503), .QN(n3532) );
  NAND2X0 U4947 ( .IN1(n3534), .IN2(n3535), .QN(P2_N2177) );
  NAND2X0 U4948 ( .IN1(P2_N2118), .IN2(n3512), .QN(n3535) );
  NAND2X0 U4949 ( .IN1(P2_N381), .IN2(P2_N5503), .QN(n3534) );
  NAND2X0 U4950 ( .IN1(n3536), .IN2(n3537), .QN(P2_N2176) );
  NAND2X0 U4951 ( .IN1(P2_N2117), .IN2(n3512), .QN(n3537) );
  NAND2X0 U4952 ( .IN1(P2_N380), .IN2(P2_N5503), .QN(n3536) );
  NAND2X0 U4953 ( .IN1(n3538), .IN2(n3539), .QN(P2_N2175) );
  NAND2X0 U4954 ( .IN1(P2_N2116), .IN2(n3512), .QN(n3539) );
  NAND2X0 U4955 ( .IN1(P2_N379), .IN2(P2_N5503), .QN(n3538) );
  NAND2X0 U4956 ( .IN1(n3540), .IN2(n3541), .QN(P2_N2174) );
  NAND2X0 U4957 ( .IN1(P2_N2115), .IN2(n3512), .QN(n3541) );
  NAND2X0 U4958 ( .IN1(P2_N378), .IN2(P2_N5503), .QN(n3540) );
  NAND2X0 U4959 ( .IN1(n3542), .IN2(n3543), .QN(P2_N2173) );
  NAND2X0 U4960 ( .IN1(P2_N2114), .IN2(n3512), .QN(n3543) );
  NAND2X0 U4961 ( .IN1(P2_N377), .IN2(P2_N5503), .QN(n3542) );
  NAND2X0 U4962 ( .IN1(n3544), .IN2(n3545), .QN(P2_N2172) );
  NAND2X0 U4963 ( .IN1(P2_N2113), .IN2(n3512), .QN(n3545) );
  NAND2X0 U4964 ( .IN1(P2_N376), .IN2(P2_N5503), .QN(n3544) );
  NAND2X0 U4965 ( .IN1(n3546), .IN2(n3547), .QN(P2_N2171) );
  NAND2X0 U4966 ( .IN1(P2_N2112), .IN2(n3512), .QN(n3547) );
  NAND2X0 U4967 ( .IN1(P2_N375), .IN2(P2_N5503), .QN(n3546) );
  NAND2X0 U4968 ( .IN1(n3548), .IN2(n3549), .QN(P2_N2170) );
  NAND2X0 U4969 ( .IN1(P2_N2111), .IN2(n3512), .QN(n3549) );
  NAND2X0 U4970 ( .IN1(P2_N374), .IN2(P2_N5503), .QN(n3548) );
  NAND2X0 U4971 ( .IN1(n3550), .IN2(n3551), .QN(P2_N2169) );
  NAND2X0 U4972 ( .IN1(P2_N2110), .IN2(n3512), .QN(n3551) );
  NAND2X0 U4973 ( .IN1(P2_N373), .IN2(P2_N5503), .QN(n3550) );
  NAND2X0 U4974 ( .IN1(n3552), .IN2(n3553), .QN(P2_N2168) );
  NAND2X0 U4975 ( .IN1(P2_N2109), .IN2(n3512), .QN(n3553) );
  NAND2X0 U4976 ( .IN1(P2_N372), .IN2(P2_N5503), .QN(n3552) );
  NAND2X0 U4977 ( .IN1(n3554), .IN2(n3555), .QN(P2_N2167) );
  NAND2X0 U4978 ( .IN1(P2_N2108), .IN2(n3512), .QN(n3555) );
  NAND2X0 U4979 ( .IN1(P2_N371), .IN2(P2_N5503), .QN(n3554) );
  NAND2X0 U4980 ( .IN1(n3556), .IN2(n3557), .QN(P2_N2166) );
  NAND2X0 U4981 ( .IN1(P2_N2107), .IN2(n3512), .QN(n3557) );
  NAND2X0 U4982 ( .IN1(P2_N370), .IN2(P2_N5503), .QN(n3556) );
  NAND2X0 U4983 ( .IN1(n3558), .IN2(n3559), .QN(P2_N2165) );
  NAND2X0 U4984 ( .IN1(P2_N2106), .IN2(n3512), .QN(n3559) );
  NAND2X0 U4985 ( .IN1(P2_N369), .IN2(P2_N5503), .QN(n3558) );
  NAND2X0 U4986 ( .IN1(n3560), .IN2(n3561), .QN(P2_N2164) );
  NAND2X0 U4987 ( .IN1(P2_N2105), .IN2(n3512), .QN(n3561) );
  NAND2X0 U4988 ( .IN1(P2_N368), .IN2(P2_N5503), .QN(n3560) );
  NAND2X0 U4989 ( .IN1(n3562), .IN2(n3563), .QN(P2_N2163) );
  NAND2X0 U4990 ( .IN1(P2_N2104), .IN2(n3512), .QN(n3563) );
  NAND2X0 U4991 ( .IN1(n18813), .IN2(P2_N5503), .QN(n3562) );
  NAND2X0 U4798 ( .IN1(P2_N373), .IN2(P2_N5504), .QN(n3441) );
  NAND2X0 U4799 ( .IN1(n3443), .IN2(n3444), .QN(P2_N2541) );
  NAND2X0 U4800 ( .IN1(P2_N2482), .IN2(n3403), .QN(n3444) );
  NAND2X0 U4801 ( .IN1(P2_N372), .IN2(P2_N5504), .QN(n3443) );
  NAND2X0 U4802 ( .IN1(n3445), .IN2(n3446), .QN(P2_N2540) );
  NAND2X0 U4803 ( .IN1(P2_N2481), .IN2(n3403), .QN(n3446) );
  NAND2X0 U4804 ( .IN1(P2_N371), .IN2(P2_N5504), .QN(n3445) );
  NAND2X0 U4805 ( .IN1(n3447), .IN2(n3448), .QN(P2_N2539) );
  NAND2X0 U4806 ( .IN1(P2_N2480), .IN2(n3403), .QN(n3448) );
  NAND2X0 U4807 ( .IN1(P2_N370), .IN2(P2_N5504), .QN(n3447) );
  NAND2X0 U4808 ( .IN1(n3449), .IN2(n3450), .QN(P2_N2538) );
  NAND2X0 U4809 ( .IN1(P2_N2479), .IN2(n3403), .QN(n3450) );
  NAND2X0 U4810 ( .IN1(P2_N369), .IN2(P2_N5504), .QN(n3449) );
  NAND2X0 U4811 ( .IN1(n3451), .IN2(n3452), .QN(P2_N2537) );
  NAND2X0 U4812 ( .IN1(P2_N2478), .IN2(n3403), .QN(n3452) );
  NAND2X0 U4813 ( .IN1(P2_N368), .IN2(P2_N5504), .QN(n3451) );
  NAND2X0 U4814 ( .IN1(n3453), .IN2(n3454), .QN(P2_N2536) );
  NAND2X0 U4815 ( .IN1(P2_N2477), .IN2(n3403), .QN(n3454) );
  NAND2X0 U4816 ( .IN1(n18813), .IN2(P2_N5504), .QN(n3453) );
  NAND2X0 U4817 ( .IN1(n3455), .IN2(n3456), .QN(P2_N2535) );
  NAND2X0 U4818 ( .IN1(P2_N2476), .IN2(n3403), .QN(n3456) );
  NAND2X0 U4819 ( .IN1(n6683), .IN2(P2_N5504), .QN(n3455) );
  NAND2X0 U4820 ( .IN1(n3457), .IN2(n3458), .QN(P2_N2534) );
  NAND2X0 U4821 ( .IN1(P2_N2475), .IN2(n3403), .QN(n3458) );
  NAND2X0 U4822 ( .IN1(n6682), .IN2(P2_N5504), .QN(n3457) );
  NAND2X0 U4823 ( .IN1(n3459), .IN2(n3460), .QN(P2_N2533) );
  NAND2X0 U4824 ( .IN1(P2_N2474), .IN2(n3403), .QN(n3460) );
  NAND2X0 U4827 ( .IN1(n6681), .IN2(P2_N5504), .QN(n3459) );
  AND2X1 U4832 ( .IN1(P2_N193), .IN2(n3463), .Q(P2_N244) );
  NAND2X0 U4833 ( .IN1(n3464), .IN2(n3465), .QN(n3463) );
  NOR2X0 U4834 ( .QN(n3465), .IN1(n3466), .IN2(n3467) );
  NAND2X0 U4835 ( .IN1(n3468), .IN2(n3469), .QN(n3467) );
  NOR2X0 U4836 ( .QN(n3469), .IN1(P2_N212), .IN2(n3470) );
  OR2X1 U4837 ( .IN2(P2_N213), .IN1(P2_N214), .Q(n3470) );
  NOR2X0 U4838 ( .QN(n3468), .IN1(P2_N209), .IN2(n3471) );
  OR2X1 U4839 ( .IN2(P2_N210), .IN1(P2_N211), .Q(n3471) );
  NAND2X0 U4840 ( .IN1(n3472), .IN2(n3473), .QN(n3466) );
  NOR2X0 U4841 ( .QN(n3473), .IN1(P2_N218), .IN2(n3474) );
  OR2X1 U4842 ( .IN2(P2_N219), .IN1(P2_N220), .Q(n3474) );
  NOR2X0 U4843 ( .QN(n3472), .IN1(P2_N215), .IN2(n3475) );
  OR2X1 U4844 ( .IN2(P2_N216), .IN1(P2_N217), .Q(n3475) );
  NOR2X0 U4845 ( .QN(n3464), .IN1(n3476), .IN2(n3477) );
  NAND2X0 U4846 ( .IN1(n3478), .IN2(n3479), .QN(n3477) );
  NOR2X0 U4847 ( .QN(n3479), .IN1(P2_N200), .IN2(n3480) );
  OR2X1 U4848 ( .IN2(P2_N201), .IN1(P2_N202), .Q(n3480) );
  NOR2X0 U4849 ( .QN(n3478), .IN1(P2_N197), .IN2(n3481) );
  OR2X1 U4850 ( .IN2(P2_N198), .IN1(P2_N199), .Q(n3481) );
  NAND2X0 U4851 ( .IN1(n3482), .IN2(n3483), .QN(n3476) );
  NOR2X0 U4852 ( .QN(n3483), .IN1(P2_N206), .IN2(n3484) );
  OR2X1 U4853 ( .IN2(P2_N207), .IN1(P2_N208), .Q(n3484) );
  NOR2X0 U4854 ( .QN(n3482), .IN1(P2_N203), .IN2(n3485) );
  OR2X1 U4855 ( .IN2(P2_N204), .IN1(P2_N205), .Q(n3485) );
  NAND2X0 U4856 ( .IN1(n7386), .IN2(n3486), .QN(P2_N2381) );
  NAND2X0 U4857 ( .IN1(n7385), .IN2(n3487), .QN(P2_N2379) );
  NOR2X0 U4858 ( .QN(P2_N2562), .IN1(n3487), .IN2(n3486) );
  INVX0 U4859 ( .ZN(n3486), .INP(n7385) );
  INVX0 U4860 ( .ZN(n3487), .INP(n7386) );
  NOR2X0 U4861 ( .QN(P2_N2261), .IN1(n7329), .IN2(n7007) );
  NOR2X0 U4862 ( .QN(P2_N2260), .IN1(n7327), .IN2(n7007) );
  NOR2X0 U4863 ( .QN(P2_N2259), .IN1(n7325), .IN2(n7007) );
  NOR2X0 U4864 ( .QN(P2_N2258), .IN1(n7323), .IN2(n7011) );
  NOR2X0 U4865 ( .QN(P2_N2257), .IN1(n7321), .IN2(n7011) );
  NOR2X0 U4866 ( .QN(P2_N2256), .IN1(n7319), .IN2(n7011) );
  NOR2X0 U4867 ( .QN(P2_N2255), .IN1(n7317), .IN2(n7011) );
  NOR2X0 U4868 ( .QN(P2_N2254), .IN1(n7315), .IN2(n7015) );
  NOR2X0 U4869 ( .QN(P2_N2253), .IN1(n7313), .IN2(n7015) );
  NOR2X0 U4870 ( .QN(P2_N2252), .IN1(n7311), .IN2(n7015) );
  NAND2X0 U4872 ( .IN1(n2006), .IN2(n3489), .QN(P2_N2251) );
  NAND2X0 U4873 ( .IN1(n7012), .IN2(n2008), .QN(n3489) );
  NAND2X0 U4874 ( .IN1(n2009), .IN2(n3490), .QN(P2_N2250) );
  NAND2X0 U4875 ( .IN1(n7012), .IN2(n2011), .QN(n3490) );
  NAND2X0 U4876 ( .IN1(n2012), .IN2(n3491), .QN(P2_N2249) );
  NAND2X0 U4877 ( .IN1(n7012), .IN2(n2014), .QN(n3491) );
  NAND2X0 U4878 ( .IN1(n2015), .IN2(n3492), .QN(P2_N2248) );
  NAND2X0 U4879 ( .IN1(n7012), .IN2(n2017), .QN(n3492) );
  NAND2X0 U4880 ( .IN1(n2018), .IN2(n3493), .QN(P2_N2247) );
  NAND2X0 U4881 ( .IN1(n7009), .IN2(n2020), .QN(n3493) );
  NAND2X0 U4882 ( .IN1(n2021), .IN2(n3494), .QN(P2_N2246) );
  NAND2X0 U4883 ( .IN1(n7009), .IN2(n2023), .QN(n3494) );
  NAND2X0 U4884 ( .IN1(n2024), .IN2(n3495), .QN(P2_N2245) );
  NAND2X0 U4885 ( .IN1(n7009), .IN2(n2026), .QN(n3495) );
  NAND2X0 U4886 ( .IN1(n2027), .IN2(n3496), .QN(P2_N2244) );
  NAND2X0 U4887 ( .IN1(n7009), .IN2(n2029), .QN(n3496) );
  NAND2X0 U4888 ( .IN1(n2030), .IN2(n3497), .QN(P2_N2243) );
  NAND2X0 U4889 ( .IN1(n7010), .IN2(n2032), .QN(n3497) );
  NAND2X0 U4890 ( .IN1(n2033), .IN2(n3498), .QN(P2_N2242) );
  NAND2X0 U4891 ( .IN1(n7010), .IN2(n2035), .QN(n3498) );
  NAND2X0 U4892 ( .IN1(n2036), .IN2(n3499), .QN(P2_N2241) );
  NAND2X0 U4893 ( .IN1(n7016), .IN2(n2038), .QN(n3499) );
  NAND2X0 U4894 ( .IN1(n2039), .IN2(n3500), .QN(P2_N2240) );
  NAND2X0 U4895 ( .IN1(n7016), .IN2(n2041), .QN(n3500) );
  NAND2X0 U4896 ( .IN1(n2042), .IN2(n3501), .QN(P2_N2239) );
  NAND2X0 U4703 ( .IN1(n2015), .IN2(n3383), .QN(P2_N2621) );
  NAND2X0 U4704 ( .IN1(n7012), .IN2(n2017), .QN(n3383) );
  NAND2X0 U4705 ( .IN1(n2018), .IN2(n3384), .QN(P2_N2620) );
  NAND2X0 U4706 ( .IN1(n7009), .IN2(n2020), .QN(n3384) );
  NAND2X0 U4707 ( .IN1(n2021), .IN2(n3385), .QN(P2_N2619) );
  NAND2X0 U4708 ( .IN1(n7009), .IN2(n2023), .QN(n3385) );
  NAND2X0 U4709 ( .IN1(n2024), .IN2(n3386), .QN(P2_N2618) );
  NAND2X0 U4710 ( .IN1(n7009), .IN2(n2026), .QN(n3386) );
  NAND2X0 U4711 ( .IN1(n2027), .IN2(n3387), .QN(P2_N2617) );
  NAND2X0 U4712 ( .IN1(n7009), .IN2(n2029), .QN(n3387) );
  NAND2X0 U4713 ( .IN1(n2030), .IN2(n3388), .QN(P2_N2616) );
  NAND2X0 U4714 ( .IN1(n7010), .IN2(n2032), .QN(n3388) );
  NAND2X0 U4715 ( .IN1(n2033), .IN2(n3389), .QN(P2_N2615) );
  NAND2X0 U4716 ( .IN1(n7010), .IN2(n2035), .QN(n3389) );
  NAND2X0 U4717 ( .IN1(n2036), .IN2(n3390), .QN(P2_N2614) );
  NAND2X0 U4718 ( .IN1(n7016), .IN2(n2038), .QN(n3390) );
  NAND2X0 U4719 ( .IN1(n2039), .IN2(n3391), .QN(P2_N2613) );
  NAND2X0 U4720 ( .IN1(n7016), .IN2(n2041), .QN(n3391) );
  NAND2X0 U4721 ( .IN1(n2042), .IN2(n3392), .QN(P2_N2612) );
  NAND2X0 U4722 ( .IN1(n7016), .IN2(n2044), .QN(n3392) );
  NAND2X0 U4723 ( .IN1(n2045), .IN2(n3393), .QN(P2_N2611) );
  NAND2X0 U4724 ( .IN1(n7016), .IN2(n2047), .QN(n3393) );
  NAND2X0 U4725 ( .IN1(n2048), .IN2(n3394), .QN(P2_N2610) );
  NAND2X0 U4726 ( .IN1(n7006), .IN2(n2050), .QN(n3394) );
  NAND2X0 U4727 ( .IN1(n2051), .IN2(n3395), .QN(P2_N2609) );
  NAND2X0 U4728 ( .IN1(n7006), .IN2(n2053), .QN(n3395) );
  NAND2X0 U4729 ( .IN1(n2054), .IN2(n3396), .QN(P2_N2608) );
  NAND2X0 U4730 ( .IN1(n7006), .IN2(n2056), .QN(n3396) );
  NAND2X0 U4731 ( .IN1(n2057), .IN2(n3397), .QN(P2_N2607) );
  NAND2X0 U4732 ( .IN1(n7462), .IN2(n2059), .QN(n3397) );
  NAND2X0 U4733 ( .IN1(n2060), .IN2(n3398), .QN(P2_N2606) );
  NAND2X0 U4734 ( .IN1(n7462), .IN2(n2062), .QN(n3398) );
  NAND2X0 U4735 ( .IN1(n2063), .IN2(n3399), .QN(P2_N2605) );
  NAND2X0 U4736 ( .IN1(n7462), .IN2(n2065), .QN(n3399) );
  NAND2X0 U4739 ( .IN1(n3401), .IN2(n3402), .QN(P2_N2561) );
  NAND2X0 U4740 ( .IN1(P2_N2502), .IN2(n3403), .QN(n3402) );
  NAND2X0 U4741 ( .IN1(P2_N392), .IN2(P2_N5504), .QN(n3401) );
  NAND2X0 U4742 ( .IN1(n3405), .IN2(n3406), .QN(P2_N2560) );
  NAND2X0 U4743 ( .IN1(P2_N2501), .IN2(n3403), .QN(n3406) );
  NAND2X0 U4744 ( .IN1(P2_N391), .IN2(P2_N5504), .QN(n3405) );
  NAND2X0 U4745 ( .IN1(n3407), .IN2(n3408), .QN(P2_N2559) );
  NAND2X0 U4746 ( .IN1(P2_N2500), .IN2(n3403), .QN(n3408) );
  NAND2X0 U4747 ( .IN1(P2_N390), .IN2(P2_N5504), .QN(n3407) );
  NAND2X0 U4748 ( .IN1(n3409), .IN2(n3410), .QN(P2_N2558) );
  NAND2X0 U4749 ( .IN1(P2_N2499), .IN2(n3403), .QN(n3410) );
  NAND2X0 U4750 ( .IN1(P2_N389), .IN2(P2_N5504), .QN(n3409) );
  NAND2X0 U4751 ( .IN1(n3411), .IN2(n3412), .QN(P2_N2557) );
  NAND2X0 U4752 ( .IN1(P2_N2498), .IN2(n3403), .QN(n3412) );
  NAND2X0 U4753 ( .IN1(P2_N388), .IN2(P2_N5504), .QN(n3411) );
  NAND2X0 U4754 ( .IN1(n3413), .IN2(n3414), .QN(P2_N2556) );
  NAND2X0 U4755 ( .IN1(P2_N2497), .IN2(n3403), .QN(n3414) );
  NAND2X0 U4756 ( .IN1(P2_N387), .IN2(P2_N5504), .QN(n3413) );
  NAND2X0 U4757 ( .IN1(n3415), .IN2(n3416), .QN(P2_N2555) );
  NAND2X0 U4758 ( .IN1(P2_N2496), .IN2(n3403), .QN(n3416) );
  NAND2X0 U4759 ( .IN1(P2_N386), .IN2(P2_N5504), .QN(n3415) );
  NAND2X0 U4760 ( .IN1(n3417), .IN2(n3418), .QN(P2_N2554) );
  NAND2X0 U4761 ( .IN1(P2_N2495), .IN2(n3403), .QN(n3418) );
  NAND2X0 U4762 ( .IN1(P2_N385), .IN2(P2_N5504), .QN(n3417) );
  NAND2X0 U4763 ( .IN1(n3419), .IN2(n3420), .QN(P2_N2553) );
  NAND2X0 U4764 ( .IN1(P2_N2494), .IN2(n3403), .QN(n3420) );
  NAND2X0 U4765 ( .IN1(P2_N384), .IN2(P2_N5504), .QN(n3419) );
  NAND2X0 U4766 ( .IN1(n3421), .IN2(n3422), .QN(P2_N2552) );
  NAND2X0 U4767 ( .IN1(P2_N2493), .IN2(n3403), .QN(n3422) );
  NAND2X0 U4768 ( .IN1(P2_N383), .IN2(P2_N5504), .QN(n3421) );
  NAND2X0 U4769 ( .IN1(n3423), .IN2(n3424), .QN(P2_N2551) );
  NAND2X0 U4770 ( .IN1(P2_N2492), .IN2(n3403), .QN(n3424) );
  NAND2X0 U4771 ( .IN1(P2_N382), .IN2(P2_N5504), .QN(n3423) );
  NAND2X0 U4772 ( .IN1(n3425), .IN2(n3426), .QN(P2_N2550) );
  NAND2X0 U4773 ( .IN1(P2_N2491), .IN2(n3403), .QN(n3426) );
  NAND2X0 U4774 ( .IN1(P2_N381), .IN2(P2_N5504), .QN(n3425) );
  NAND2X0 U4775 ( .IN1(n3427), .IN2(n3428), .QN(P2_N2549) );
  NAND2X0 U4776 ( .IN1(P2_N2490), .IN2(n3403), .QN(n3428) );
  NAND2X0 U4777 ( .IN1(P2_N380), .IN2(P2_N5504), .QN(n3427) );
  NAND2X0 U4778 ( .IN1(n3429), .IN2(n3430), .QN(P2_N2548) );
  NAND2X0 U4779 ( .IN1(P2_N2489), .IN2(n3403), .QN(n3430) );
  NAND2X0 U4780 ( .IN1(P2_N379), .IN2(P2_N5504), .QN(n3429) );
  NAND2X0 U4781 ( .IN1(n3431), .IN2(n3432), .QN(P2_N2547) );
  NAND2X0 U4782 ( .IN1(P2_N2488), .IN2(n3403), .QN(n3432) );
  NAND2X0 U4783 ( .IN1(P2_N378), .IN2(P2_N5504), .QN(n3431) );
  NAND2X0 U4784 ( .IN1(n3433), .IN2(n3434), .QN(P2_N2546) );
  NAND2X0 U4785 ( .IN1(P2_N2487), .IN2(n3403), .QN(n3434) );
  NAND2X0 U4786 ( .IN1(P2_N377), .IN2(P2_N5504), .QN(n3433) );
  NAND2X0 U4787 ( .IN1(n3435), .IN2(n3436), .QN(P2_N2545) );
  NAND2X0 U4788 ( .IN1(P2_N2486), .IN2(n3403), .QN(n3436) );
  NAND2X0 U4789 ( .IN1(P2_N376), .IN2(P2_N5504), .QN(n3435) );
  NAND2X0 U4790 ( .IN1(n3437), .IN2(n3438), .QN(P2_N2544) );
  NAND2X0 U4791 ( .IN1(P2_N2485), .IN2(n3403), .QN(n3438) );
  NAND2X0 U4792 ( .IN1(P2_N375), .IN2(P2_N5504), .QN(n3437) );
  NAND2X0 U4793 ( .IN1(n3439), .IN2(n3440), .QN(P2_N2543) );
  NAND2X0 U4794 ( .IN1(P2_N2484), .IN2(n3403), .QN(n3440) );
  NAND2X0 U4795 ( .IN1(P2_N374), .IN2(P2_N5504), .QN(n3439) );
  NAND2X0 U4796 ( .IN1(n3441), .IN2(n3442), .QN(P2_N2542) );
  NAND2X0 U4797 ( .IN1(P2_N2483), .IN2(n3403), .QN(n3442) );
  NAND2X0 U4604 ( .IN1(P2_N381), .IN2(P2_N5505), .QN(n3321) );
  NAND2X0 U4605 ( .IN1(n3323), .IN2(n3324), .QN(P2_N2922) );
  NAND2X0 U4606 ( .IN1(P2_N2863), .IN2(n3299), .QN(n3324) );
  NAND2X0 U4607 ( .IN1(P2_N380), .IN2(P2_N5505), .QN(n3323) );
  NAND2X0 U4608 ( .IN1(n3325), .IN2(n3326), .QN(P2_N2921) );
  NAND2X0 U4609 ( .IN1(P2_N2862), .IN2(n3299), .QN(n3326) );
  NAND2X0 U4610 ( .IN1(P2_N379), .IN2(P2_N5505), .QN(n3325) );
  NAND2X0 U4611 ( .IN1(n3327), .IN2(n3328), .QN(P2_N2920) );
  NAND2X0 U4612 ( .IN1(P2_N2861), .IN2(n3299), .QN(n3328) );
  NAND2X0 U4613 ( .IN1(P2_N378), .IN2(P2_N5505), .QN(n3327) );
  NAND2X0 U4614 ( .IN1(n3329), .IN2(n3330), .QN(P2_N2919) );
  NAND2X0 U4615 ( .IN1(P2_N2860), .IN2(n3299), .QN(n3330) );
  NAND2X0 U4616 ( .IN1(P2_N377), .IN2(P2_N5505), .QN(n3329) );
  NAND2X0 U4617 ( .IN1(n3331), .IN2(n3332), .QN(P2_N2918) );
  NAND2X0 U4618 ( .IN1(P2_N2859), .IN2(n3299), .QN(n3332) );
  NAND2X0 U4619 ( .IN1(P2_N376), .IN2(P2_N5505), .QN(n3331) );
  NAND2X0 U4620 ( .IN1(n3333), .IN2(n3334), .QN(P2_N2917) );
  NAND2X0 U4621 ( .IN1(P2_N2858), .IN2(n3299), .QN(n3334) );
  NAND2X0 U4622 ( .IN1(P2_N375), .IN2(P2_N5505), .QN(n3333) );
  NAND2X0 U4623 ( .IN1(n3335), .IN2(n3336), .QN(P2_N2916) );
  NAND2X0 U4624 ( .IN1(P2_N2857), .IN2(n3299), .QN(n3336) );
  NAND2X0 U4625 ( .IN1(P2_N374), .IN2(P2_N5505), .QN(n3335) );
  NAND2X0 U4626 ( .IN1(n3337), .IN2(n3338), .QN(P2_N2915) );
  NAND2X0 U4627 ( .IN1(P2_N2856), .IN2(n3299), .QN(n3338) );
  NAND2X0 U4628 ( .IN1(P2_N373), .IN2(P2_N5505), .QN(n3337) );
  NAND2X0 U4629 ( .IN1(n3339), .IN2(n3340), .QN(P2_N2914) );
  NAND2X0 U4630 ( .IN1(P2_N2855), .IN2(n3299), .QN(n3340) );
  NAND2X0 U4631 ( .IN1(P2_N372), .IN2(P2_N5505), .QN(n3339) );
  NAND2X0 U4632 ( .IN1(n3341), .IN2(n3342), .QN(P2_N2913) );
  NAND2X0 U4633 ( .IN1(P2_N2854), .IN2(n3299), .QN(n3342) );
  NAND2X0 U4634 ( .IN1(P2_N371), .IN2(P2_N5505), .QN(n3341) );
  NAND2X0 U4635 ( .IN1(n3343), .IN2(n3344), .QN(P2_N2912) );
  NAND2X0 U4636 ( .IN1(P2_N2853), .IN2(n3299), .QN(n3344) );
  NAND2X0 U4637 ( .IN1(P2_N370), .IN2(P2_N5505), .QN(n3343) );
  NAND2X0 U4638 ( .IN1(n3345), .IN2(n3346), .QN(P2_N2911) );
  NAND2X0 U4639 ( .IN1(P2_N2852), .IN2(n3299), .QN(n3346) );
  NAND2X0 U4640 ( .IN1(P2_N369), .IN2(P2_N5505), .QN(n3345) );
  NAND2X0 U4641 ( .IN1(n3347), .IN2(n3348), .QN(P2_N2910) );
  NAND2X0 U4642 ( .IN1(P2_N2851), .IN2(n3299), .QN(n3348) );
  NAND2X0 U4643 ( .IN1(P2_N368), .IN2(P2_N5505), .QN(n3347) );
  NAND2X0 U4644 ( .IN1(n3349), .IN2(n3350), .QN(P2_N2909) );
  NAND2X0 U4645 ( .IN1(P2_N2850), .IN2(n3299), .QN(n3350) );
  NAND2X0 U4646 ( .IN1(n18813), .IN2(P2_N5505), .QN(n3349) );
  NAND2X0 U4647 ( .IN1(n3351), .IN2(n3352), .QN(P2_N2908) );
  NAND2X0 U4648 ( .IN1(P2_N2849), .IN2(n3299), .QN(n3352) );
  NAND2X0 U4649 ( .IN1(n6683), .IN2(P2_N5505), .QN(n3351) );
  NAND2X0 U4650 ( .IN1(n3353), .IN2(n3354), .QN(P2_N2907) );
  NAND2X0 U4651 ( .IN1(P2_N2848), .IN2(n3299), .QN(n3354) );
  NAND2X0 U4652 ( .IN1(n6682), .IN2(P2_N5505), .QN(n3353) );
  NAND2X0 U4653 ( .IN1(n3355), .IN2(n3356), .QN(P2_N2906) );
  NAND2X0 U4654 ( .IN1(P2_N2847), .IN2(n3299), .QN(n3356) );
  NAND2X0 U4657 ( .IN1(n6681), .IN2(P2_N5505), .QN(n3355) );
  AND2X1 U4662 ( .IN1(P2_N248), .IN2(n3359), .Q(P2_N290) );
  NAND2X0 U4663 ( .IN1(n3360), .IN2(n3361), .QN(n3359) );
  NOR2X0 U4664 ( .QN(n3361), .IN1(n3362), .IN2(n3363) );
  NAND2X0 U4665 ( .IN1(n3364), .IN2(n3365), .QN(n3363) );
  NOR2X0 U4666 ( .QN(n3365), .IN1(P2_N264), .IN2(n3366) );
  OR2X1 U4667 ( .IN2(P2_N265), .IN1(P2_N266), .Q(n3366) );
  NOR2X0 U4668 ( .QN(n3364), .IN1(P2_N263), .IN2(P2_N262) );
  NAND2X0 U4669 ( .IN1(n3367), .IN2(n3368), .QN(n3362) );
  NOR2X0 U4670 ( .QN(n3368), .IN1(P2_N269), .IN2(n3369) );
  OR2X1 U4671 ( .IN2(P2_N270), .IN1(P2_N271), .Q(n3369) );
  NOR2X0 U4672 ( .QN(n3367), .IN1(P2_N268), .IN2(P2_N267) );
  NOR2X0 U4673 ( .QN(n3360), .IN1(n3370), .IN2(n3371) );
  NAND2X0 U4674 ( .IN1(n3372), .IN2(n3373), .QN(n3371) );
  NOR2X0 U4675 ( .QN(n3373), .IN1(P2_N256), .IN2(P2_N255) );
  NOR2X0 U4676 ( .QN(n3372), .IN1(P2_N254), .IN2(P2_N253) );
  NAND2X0 U4677 ( .IN1(n3374), .IN2(n3375), .QN(n3370) );
  NOR2X0 U4678 ( .QN(n3375), .IN1(P2_N259), .IN2(n3376) );
  OR2X1 U4679 ( .IN2(P2_N260), .IN1(P2_N261), .Q(n3376) );
  NOR2X0 U4680 ( .QN(n3374), .IN1(P2_N258), .IN2(P2_N257) );
  NAND2X0 U4681 ( .IN1(n7388), .IN2(n3377), .QN(P2_N2754) );
  NAND2X0 U4682 ( .IN1(n7387), .IN2(n3378), .QN(P2_N2752) );
  NOR2X0 U4683 ( .QN(P2_N2935), .IN1(n3378), .IN2(n3377) );
  INVX0 U4684 ( .ZN(n3377), .INP(n7387) );
  INVX0 U4685 ( .ZN(n3378), .INP(n7388) );
  NOR2X0 U4686 ( .QN(P2_N2634), .IN1(n7329), .IN2(n7007) );
  NOR2X0 U4687 ( .QN(P2_N2633), .IN1(n7327), .IN2(n7007) );
  NOR2X0 U4688 ( .QN(P2_N2632), .IN1(n7325), .IN2(n7007) );
  NOR2X0 U4689 ( .QN(P2_N2631), .IN1(n7323), .IN2(n7011) );
  NOR2X0 U4690 ( .QN(P2_N2630), .IN1(n7321), .IN2(n7011) );
  NOR2X0 U4691 ( .QN(P2_N2629), .IN1(n7319), .IN2(n7011) );
  NOR2X0 U4692 ( .QN(P2_N2628), .IN1(n7317), .IN2(n7011) );
  NOR2X0 U4693 ( .QN(P2_N2627), .IN1(n7315), .IN2(n7015) );
  NOR2X0 U4694 ( .QN(P2_N2626), .IN1(n7313), .IN2(n7015) );
  NOR2X0 U4695 ( .QN(P2_N2625), .IN1(n7311), .IN2(n7011) );
  NAND2X0 U4697 ( .IN1(n2006), .IN2(n3380), .QN(P2_N2624) );
  NAND2X0 U4698 ( .IN1(n7012), .IN2(n2008), .QN(n3380) );
  NAND2X0 U4699 ( .IN1(n2009), .IN2(n3381), .QN(P2_N2623) );
  NAND2X0 U4700 ( .IN1(n7012), .IN2(n2011), .QN(n3381) );
  NAND2X0 U4701 ( .IN1(n2012), .IN2(n3382), .QN(P2_N2622) );
  NAND2X0 U4702 ( .IN1(P2_N914), .IN2(n2014), .QN(n3382) );
  NAND2X0 U4503 ( .IN1(P2_N3220), .IN2(n3213), .QN(n3270) );
  NAND2X0 U4506 ( .IN1(n6681), .IN2(P2_N5506), .QN(n3269) );
  NAND2X0 U4511 ( .IN1(n7390), .IN2(n3273), .QN(P2_N3127) );
  NAND2X0 U4512 ( .IN1(n7389), .IN2(n3274), .QN(P2_N3125) );
  NOR2X0 U4513 ( .QN(P2_N3308), .IN1(n3274), .IN2(n3273) );
  INVX0 U4514 ( .ZN(n3273), .INP(n7389) );
  INVX0 U4515 ( .ZN(n3274), .INP(n7390) );
  NOR2X0 U4516 ( .QN(P2_N3007), .IN1(n7329), .IN2(n7007) );
  NOR2X0 U4517 ( .QN(P2_N3006), .IN1(n7327), .IN2(n7007) );
  NOR2X0 U4518 ( .QN(P2_N3005), .IN1(n7325), .IN2(n7007) );
  NOR2X0 U4519 ( .QN(P2_N3004), .IN1(n7323), .IN2(n7011) );
  NOR2X0 U4520 ( .QN(P2_N3003), .IN1(n7321), .IN2(n7011) );
  NOR2X0 U4521 ( .QN(P2_N3002), .IN1(n7319), .IN2(n7011) );
  NOR2X0 U4522 ( .QN(P2_N3001), .IN1(n7317), .IN2(n7011) );
  NOR2X0 U4523 ( .QN(P2_N3000), .IN1(n7315), .IN2(n7015) );
  NOR2X0 U4524 ( .QN(P2_N2999), .IN1(n7313), .IN2(n7015) );
  NOR2X0 U4525 ( .QN(P2_N2998), .IN1(n7311), .IN2(n7015) );
  NAND2X0 U4527 ( .IN1(n2006), .IN2(n3276), .QN(P2_N2997) );
  NAND2X0 U4528 ( .IN1(n7012), .IN2(n2008), .QN(n3276) );
  NAND2X0 U4529 ( .IN1(n2009), .IN2(n3277), .QN(P2_N2996) );
  NAND2X0 U4530 ( .IN1(n7012), .IN2(n2011), .QN(n3277) );
  NAND2X0 U4531 ( .IN1(n2012), .IN2(n3278), .QN(P2_N2995) );
  NAND2X0 U4532 ( .IN1(n7012), .IN2(n2014), .QN(n3278) );
  NAND2X0 U4533 ( .IN1(n2015), .IN2(n3279), .QN(P2_N2994) );
  NAND2X0 U4534 ( .IN1(n7012), .IN2(n2017), .QN(n3279) );
  NAND2X0 U4535 ( .IN1(n2018), .IN2(n3280), .QN(P2_N2993) );
  NAND2X0 U4536 ( .IN1(n7009), .IN2(n2020), .QN(n3280) );
  NAND2X0 U4537 ( .IN1(n2021), .IN2(n3281), .QN(P2_N2992) );
  NAND2X0 U4538 ( .IN1(n7009), .IN2(n2023), .QN(n3281) );
  NAND2X0 U4539 ( .IN1(n2024), .IN2(n3282), .QN(P2_N2991) );
  NAND2X0 U4540 ( .IN1(n7009), .IN2(n2026), .QN(n3282) );
  NAND2X0 U4541 ( .IN1(n2027), .IN2(n3283), .QN(P2_N2990) );
  NAND2X0 U4542 ( .IN1(n7009), .IN2(n2029), .QN(n3283) );
  NAND2X0 U4543 ( .IN1(n2030), .IN2(n3284), .QN(P2_N2989) );
  NAND2X0 U4544 ( .IN1(n7010), .IN2(n2032), .QN(n3284) );
  NAND2X0 U4545 ( .IN1(n2033), .IN2(n3285), .QN(P2_N2988) );
  NAND2X0 U4546 ( .IN1(n7010), .IN2(n2035), .QN(n3285) );
  NAND2X0 U4547 ( .IN1(n2036), .IN2(n3286), .QN(P2_N2987) );
  NAND2X0 U4548 ( .IN1(n7016), .IN2(n2038), .QN(n3286) );
  NAND2X0 U4549 ( .IN1(n2039), .IN2(n3287), .QN(P2_N2986) );
  NAND2X0 U4550 ( .IN1(n7016), .IN2(n2041), .QN(n3287) );
  NAND2X0 U4551 ( .IN1(n2042), .IN2(n3288), .QN(P2_N2985) );
  NAND2X0 U4552 ( .IN1(n7016), .IN2(n2044), .QN(n3288) );
  NAND2X0 U4553 ( .IN1(n2045), .IN2(n3289), .QN(P2_N2984) );
  NAND2X0 U4554 ( .IN1(n7016), .IN2(n2047), .QN(n3289) );
  NAND2X0 U4555 ( .IN1(n2048), .IN2(n3290), .QN(P2_N2983) );
  NAND2X0 U4556 ( .IN1(n7016), .IN2(n2050), .QN(n3290) );
  NAND2X0 U4557 ( .IN1(n2051), .IN2(n3291), .QN(P2_N2982) );
  NAND2X0 U4558 ( .IN1(n7006), .IN2(n2053), .QN(n3291) );
  NAND2X0 U4559 ( .IN1(n2054), .IN2(n3292), .QN(P2_N2981) );
  NAND2X0 U4560 ( .IN1(n7006), .IN2(n2056), .QN(n3292) );
  NAND2X0 U4561 ( .IN1(n2057), .IN2(n3293), .QN(P2_N2980) );
  NAND2X0 U4562 ( .IN1(n7006), .IN2(n2059), .QN(n3293) );
  NAND2X0 U4563 ( .IN1(n2060), .IN2(n3294), .QN(P2_N2979) );
  NAND2X0 U4564 ( .IN1(n7006), .IN2(n2062), .QN(n3294) );
  NAND2X0 U4565 ( .IN1(n2063), .IN2(n3295), .QN(P2_N2978) );
  NAND2X0 U4566 ( .IN1(n7006), .IN2(n2065), .QN(n3295) );
  NAND2X0 U4569 ( .IN1(n3297), .IN2(n3298), .QN(P2_N2934) );
  NAND2X0 U4570 ( .IN1(P2_N2875), .IN2(n3299), .QN(n3298) );
  NAND2X0 U4571 ( .IN1(P2_N392), .IN2(P2_N5505), .QN(n3297) );
  NAND2X0 U4572 ( .IN1(n3301), .IN2(n3302), .QN(P2_N2933) );
  NAND2X0 U4573 ( .IN1(P2_N2874), .IN2(n3299), .QN(n3302) );
  NAND2X0 U4574 ( .IN1(P2_N391), .IN2(P2_N5505), .QN(n3301) );
  NAND2X0 U4575 ( .IN1(n3303), .IN2(n3304), .QN(P2_N2932) );
  NAND2X0 U4576 ( .IN1(P2_N2873), .IN2(n3299), .QN(n3304) );
  NAND2X0 U4577 ( .IN1(P2_N390), .IN2(P2_N5505), .QN(n3303) );
  NAND2X0 U4578 ( .IN1(n3305), .IN2(n3306), .QN(P2_N2931) );
  NAND2X0 U4579 ( .IN1(P2_N2872), .IN2(n3299), .QN(n3306) );
  NAND2X0 U4580 ( .IN1(P2_N389), .IN2(P2_N5505), .QN(n3305) );
  NAND2X0 U4581 ( .IN1(n3307), .IN2(n3308), .QN(P2_N2930) );
  NAND2X0 U4582 ( .IN1(P2_N2871), .IN2(n3299), .QN(n3308) );
  NAND2X0 U4583 ( .IN1(P2_N388), .IN2(P2_N5505), .QN(n3307) );
  NAND2X0 U4584 ( .IN1(n3309), .IN2(n3310), .QN(P2_N2929) );
  NAND2X0 U4585 ( .IN1(P2_N2870), .IN2(n3299), .QN(n3310) );
  NAND2X0 U4586 ( .IN1(P2_N387), .IN2(P2_N5505), .QN(n3309) );
  NAND2X0 U4587 ( .IN1(n3311), .IN2(n3312), .QN(P2_N2928) );
  NAND2X0 U4588 ( .IN1(P2_N2869), .IN2(n3299), .QN(n3312) );
  NAND2X0 U4589 ( .IN1(P2_N386), .IN2(P2_N5505), .QN(n3311) );
  NAND2X0 U4590 ( .IN1(n3313), .IN2(n3314), .QN(P2_N2927) );
  NAND2X0 U4591 ( .IN1(P2_N2868), .IN2(n3299), .QN(n3314) );
  NAND2X0 U4592 ( .IN1(P2_N385), .IN2(P2_N5505), .QN(n3313) );
  NAND2X0 U4593 ( .IN1(n3315), .IN2(n3316), .QN(P2_N2926) );
  NAND2X0 U4594 ( .IN1(P2_N2867), .IN2(n3299), .QN(n3316) );
  NAND2X0 U4595 ( .IN1(P2_N384), .IN2(P2_N5505), .QN(n3315) );
  NAND2X0 U4596 ( .IN1(n3317), .IN2(n3318), .QN(P2_N2925) );
  NAND2X0 U4597 ( .IN1(P2_N2866), .IN2(n3299), .QN(n3318) );
  NAND2X0 U4598 ( .IN1(P2_N383), .IN2(P2_N5505), .QN(n3317) );
  NAND2X0 U4599 ( .IN1(n3319), .IN2(n3320), .QN(P2_N2924) );
  NAND2X0 U4600 ( .IN1(P2_N2865), .IN2(n3299), .QN(n3320) );
  NAND2X0 U4601 ( .IN1(P2_N382), .IN2(P2_N5505), .QN(n3319) );
  NAND2X0 U4602 ( .IN1(n3321), .IN2(n3322), .QN(P2_N2923) );
  NAND2X0 U4603 ( .IN1(P2_N2864), .IN2(n3299), .QN(n3322) );
  NAND2X0 U4408 ( .IN1(n2054), .IN2(n3206), .QN(P2_N3354) );
  NAND2X0 U4409 ( .IN1(n7006), .IN2(n2056), .QN(n3206) );
  NAND2X0 U4410 ( .IN1(n2057), .IN2(n3207), .QN(P2_N3353) );
  NAND2X0 U4411 ( .IN1(n7006), .IN2(n2059), .QN(n3207) );
  NAND2X0 U4412 ( .IN1(n2060), .IN2(n3208), .QN(P2_N3352) );
  NAND2X0 U4413 ( .IN1(n7006), .IN2(n2062), .QN(n3208) );
  NAND2X0 U4414 ( .IN1(n2063), .IN2(n3209), .QN(P2_N3351) );
  NAND2X0 U4415 ( .IN1(n7462), .IN2(n2065), .QN(n3209) );
  NAND2X0 U4418 ( .IN1(n3211), .IN2(n3212), .QN(P2_N3307) );
  NAND2X0 U4419 ( .IN1(P2_N3248), .IN2(n3213), .QN(n3212) );
  NAND2X0 U4420 ( .IN1(P2_N392), .IN2(P2_N5506), .QN(n3211) );
  NAND2X0 U4421 ( .IN1(n3215), .IN2(n3216), .QN(P2_N3306) );
  NAND2X0 U4422 ( .IN1(P2_N3247), .IN2(n3213), .QN(n3216) );
  NAND2X0 U4423 ( .IN1(P2_N391), .IN2(P2_N5506), .QN(n3215) );
  NAND2X0 U4424 ( .IN1(n3217), .IN2(n3218), .QN(P2_N3305) );
  NAND2X0 U4425 ( .IN1(P2_N3246), .IN2(n3213), .QN(n3218) );
  NAND2X0 U4426 ( .IN1(P2_N390), .IN2(P2_N5506), .QN(n3217) );
  NAND2X0 U4427 ( .IN1(n3219), .IN2(n3220), .QN(P2_N3304) );
  NAND2X0 U4428 ( .IN1(P2_N3245), .IN2(n3213), .QN(n3220) );
  NAND2X0 U4429 ( .IN1(P2_N389), .IN2(P2_N5506), .QN(n3219) );
  NAND2X0 U4430 ( .IN1(n3221), .IN2(n3222), .QN(P2_N3303) );
  NAND2X0 U4431 ( .IN1(P2_N3244), .IN2(n3213), .QN(n3222) );
  NAND2X0 U4432 ( .IN1(P2_N388), .IN2(P2_N5506), .QN(n3221) );
  NAND2X0 U4433 ( .IN1(n3223), .IN2(n3224), .QN(P2_N3302) );
  NAND2X0 U4434 ( .IN1(P2_N3243), .IN2(n3213), .QN(n3224) );
  NAND2X0 U4435 ( .IN1(P2_N387), .IN2(P2_N5506), .QN(n3223) );
  NAND2X0 U4436 ( .IN1(n3225), .IN2(n3226), .QN(P2_N3301) );
  NAND2X0 U4437 ( .IN1(P2_N3242), .IN2(n3213), .QN(n3226) );
  NAND2X0 U4438 ( .IN1(P2_N386), .IN2(P2_N5506), .QN(n3225) );
  NAND2X0 U4439 ( .IN1(n3227), .IN2(n3228), .QN(P2_N3300) );
  NAND2X0 U4440 ( .IN1(P2_N3241), .IN2(n3213), .QN(n3228) );
  NAND2X0 U4441 ( .IN1(P2_N385), .IN2(P2_N5506), .QN(n3227) );
  NAND2X0 U4442 ( .IN1(n3229), .IN2(n3230), .QN(P2_N3299) );
  NAND2X0 U4443 ( .IN1(P2_N3240), .IN2(n3213), .QN(n3230) );
  NAND2X0 U4444 ( .IN1(P2_N384), .IN2(P2_N5506), .QN(n3229) );
  NAND2X0 U4445 ( .IN1(n3231), .IN2(n3232), .QN(P2_N3298) );
  NAND2X0 U4446 ( .IN1(P2_N3239), .IN2(n3213), .QN(n3232) );
  NAND2X0 U4447 ( .IN1(P2_N383), .IN2(P2_N5506), .QN(n3231) );
  NAND2X0 U4448 ( .IN1(n3233), .IN2(n3234), .QN(P2_N3297) );
  NAND2X0 U4449 ( .IN1(P2_N3238), .IN2(n3213), .QN(n3234) );
  NAND2X0 U4450 ( .IN1(P2_N382), .IN2(P2_N5506), .QN(n3233) );
  NAND2X0 U4451 ( .IN1(n3235), .IN2(n3236), .QN(P2_N3296) );
  NAND2X0 U4452 ( .IN1(P2_N3237), .IN2(n3213), .QN(n3236) );
  NAND2X0 U4453 ( .IN1(P2_N381), .IN2(P2_N5506), .QN(n3235) );
  NAND2X0 U4454 ( .IN1(n3237), .IN2(n3238), .QN(P2_N3295) );
  NAND2X0 U4455 ( .IN1(P2_N3236), .IN2(n3213), .QN(n3238) );
  NAND2X0 U4456 ( .IN1(P2_N380), .IN2(P2_N5506), .QN(n3237) );
  NAND2X0 U4457 ( .IN1(n3239), .IN2(n3240), .QN(P2_N3294) );
  NAND2X0 U4458 ( .IN1(P2_N3235), .IN2(n3213), .QN(n3240) );
  NAND2X0 U4459 ( .IN1(P2_N379), .IN2(P2_N5506), .QN(n3239) );
  NAND2X0 U4460 ( .IN1(n3241), .IN2(n3242), .QN(P2_N3293) );
  NAND2X0 U4461 ( .IN1(P2_N3234), .IN2(n3213), .QN(n3242) );
  NAND2X0 U4462 ( .IN1(P2_N378), .IN2(P2_N5506), .QN(n3241) );
  NAND2X0 U4463 ( .IN1(n3243), .IN2(n3244), .QN(P2_N3292) );
  NAND2X0 U4464 ( .IN1(P2_N3233), .IN2(n3213), .QN(n3244) );
  NAND2X0 U4465 ( .IN1(P2_N377), .IN2(P2_N5506), .QN(n3243) );
  NAND2X0 U4466 ( .IN1(n3245), .IN2(n3246), .QN(P2_N3291) );
  NAND2X0 U4467 ( .IN1(P2_N3232), .IN2(n3213), .QN(n3246) );
  NAND2X0 U4468 ( .IN1(P2_N376), .IN2(P2_N5506), .QN(n3245) );
  NAND2X0 U4469 ( .IN1(n3247), .IN2(n3248), .QN(P2_N3290) );
  NAND2X0 U4470 ( .IN1(P2_N3231), .IN2(n3213), .QN(n3248) );
  NAND2X0 U4471 ( .IN1(P2_N375), .IN2(P2_N5506), .QN(n3247) );
  NAND2X0 U4472 ( .IN1(n3249), .IN2(n3250), .QN(P2_N3289) );
  NAND2X0 U4473 ( .IN1(P2_N3230), .IN2(n3213), .QN(n3250) );
  NAND2X0 U4474 ( .IN1(P2_N374), .IN2(P2_N5506), .QN(n3249) );
  NAND2X0 U4475 ( .IN1(n3251), .IN2(n3252), .QN(P2_N3288) );
  NAND2X0 U4476 ( .IN1(P2_N3229), .IN2(n3213), .QN(n3252) );
  NAND2X0 U4477 ( .IN1(P2_N373), .IN2(P2_N5506), .QN(n3251) );
  NAND2X0 U4478 ( .IN1(n3253), .IN2(n3254), .QN(P2_N3287) );
  NAND2X0 U4479 ( .IN1(P2_N3228), .IN2(n3213), .QN(n3254) );
  NAND2X0 U4480 ( .IN1(P2_N372), .IN2(P2_N5506), .QN(n3253) );
  NAND2X0 U4481 ( .IN1(n3255), .IN2(n3256), .QN(P2_N3286) );
  NAND2X0 U4482 ( .IN1(P2_N3227), .IN2(n3213), .QN(n3256) );
  NAND2X0 U4483 ( .IN1(P2_N371), .IN2(P2_N5506), .QN(n3255) );
  NAND2X0 U4484 ( .IN1(n3257), .IN2(n3258), .QN(P2_N3285) );
  NAND2X0 U4485 ( .IN1(P2_N3226), .IN2(n3213), .QN(n3258) );
  NAND2X0 U4486 ( .IN1(P2_N370), .IN2(P2_N5506), .QN(n3257) );
  NAND2X0 U4487 ( .IN1(n3259), .IN2(n3260), .QN(P2_N3284) );
  NAND2X0 U4488 ( .IN1(P2_N3225), .IN2(n3213), .QN(n3260) );
  NAND2X0 U4489 ( .IN1(P2_N369), .IN2(P2_N5506), .QN(n3259) );
  NAND2X0 U4490 ( .IN1(n3261), .IN2(n3262), .QN(P2_N3283) );
  NAND2X0 U4491 ( .IN1(P2_N3224), .IN2(n3213), .QN(n3262) );
  NAND2X0 U4492 ( .IN1(P2_N368), .IN2(P2_N5506), .QN(n3261) );
  NAND2X0 U4493 ( .IN1(n3263), .IN2(n3264), .QN(P2_N3282) );
  NAND2X0 U4494 ( .IN1(P2_N3223), .IN2(n3213), .QN(n3264) );
  NAND2X0 U4495 ( .IN1(n18813), .IN2(P2_N5506), .QN(n3263) );
  NAND2X0 U4496 ( .IN1(n3265), .IN2(n3266), .QN(P2_N3281) );
  NAND2X0 U4497 ( .IN1(P2_N3222), .IN2(n3213), .QN(n3266) );
  NAND2X0 U4498 ( .IN1(n6683), .IN2(P2_N5506), .QN(n3265) );
  NAND2X0 U4499 ( .IN1(n3267), .IN2(n3268), .QN(P2_N3280) );
  NAND2X0 U4500 ( .IN1(P2_N3221), .IN2(n3213), .QN(n3268) );
  NAND2X0 U4501 ( .IN1(n6682), .IN2(P2_N5506), .QN(n3267) );
  NAND2X0 U4502 ( .IN1(n3269), .IN2(n3270), .QN(P2_N3279) );
  NAND2X0 U4309 ( .IN1(P2_N371), .IN2(P2_N5507), .QN(n3147) );
  NAND2X0 U4310 ( .IN1(n3149), .IN2(n3150), .QN(P2_N3658) );
  NAND2X0 U4311 ( .IN1(P2_N3599), .IN2(n3105), .QN(n3150) );
  NAND2X0 U4312 ( .IN1(P2_N370), .IN2(P2_N5507), .QN(n3149) );
  NAND2X0 U4313 ( .IN1(n3151), .IN2(n3152), .QN(P2_N3657) );
  NAND2X0 U4314 ( .IN1(P2_N3598), .IN2(n3105), .QN(n3152) );
  NAND2X0 U4315 ( .IN1(P2_N369), .IN2(P2_N5507), .QN(n3151) );
  NAND2X0 U4316 ( .IN1(n3153), .IN2(n3154), .QN(P2_N3656) );
  NAND2X0 U4317 ( .IN1(P2_N3597), .IN2(n3105), .QN(n3154) );
  NAND2X0 U4318 ( .IN1(P2_N368), .IN2(P2_N5507), .QN(n3153) );
  NAND2X0 U4319 ( .IN1(n3155), .IN2(n3156), .QN(P2_N3655) );
  NAND2X0 U4320 ( .IN1(P2_N3596), .IN2(n3105), .QN(n3156) );
  NAND2X0 U4321 ( .IN1(n18813), .IN2(P2_N5507), .QN(n3155) );
  NAND2X0 U4322 ( .IN1(n3157), .IN2(n3158), .QN(P2_N3654) );
  NAND2X0 U4323 ( .IN1(P2_N3595), .IN2(n3105), .QN(n3158) );
  NAND2X0 U4324 ( .IN1(n6683), .IN2(P2_N5507), .QN(n3157) );
  NAND2X0 U4325 ( .IN1(n3159), .IN2(n3160), .QN(P2_N3653) );
  NAND2X0 U4326 ( .IN1(P2_N3594), .IN2(n3105), .QN(n3160) );
  NAND2X0 U4327 ( .IN1(n6682), .IN2(P2_N5507), .QN(n3159) );
  NAND2X0 U4328 ( .IN1(n3161), .IN2(n3162), .QN(P2_N3652) );
  NAND2X0 U4329 ( .IN1(P2_N3593), .IN2(n3105), .QN(n3162) );
  NAND2X0 U4332 ( .IN1(n6681), .IN2(P2_N5507), .QN(n3161) );
  NAND2X0 U4337 ( .IN1(n7392), .IN2(n3165), .QN(P2_N3500) );
  NAND2X0 U4338 ( .IN1(n7391), .IN2(n3166), .QN(P2_N3498) );
  NOR2X0 U4339 ( .QN(P2_N3681), .IN1(n3166), .IN2(n3165) );
  INVX0 U4340 ( .ZN(n3165), .INP(n7391) );
  INVX0 U4341 ( .ZN(n3166), .INP(n7392) );
  AND2X1 U4342 ( .IN1(P2_N295), .IN2(n3167), .Q(P2_N342) );
  NAND2X0 U4343 ( .IN1(n3168), .IN2(n3169), .QN(n3167) );
  NOR2X0 U4344 ( .QN(n3169), .IN1(n3170), .IN2(n3171) );
  NAND2X0 U4345 ( .IN1(n3172), .IN2(n3173), .QN(n3171) );
  NOR2X0 U4346 ( .QN(n3173), .IN1(P2_N311), .IN2(n3174) );
  OR2X1 U4347 ( .IN2(P2_N312), .IN1(P2_N313), .Q(n3174) );
  NOR2X0 U4348 ( .QN(n3172), .IN1(P2_N308), .IN2(n3175) );
  OR2X1 U4349 ( .IN2(P2_N309), .IN1(P2_N310), .Q(n3175) );
  NAND2X0 U4350 ( .IN1(n3176), .IN2(n3177), .QN(n3170) );
  NOR2X0 U4351 ( .QN(n3177), .IN1(P2_N317), .IN2(n3178) );
  OR2X1 U4352 ( .IN2(P2_N318), .IN1(P2_N319), .Q(n3178) );
  NOR2X0 U4353 ( .QN(n3176), .IN1(P2_N314), .IN2(n3179) );
  OR2X1 U4354 ( .IN2(P2_N315), .IN1(P2_N316), .Q(n3179) );
  NOR2X0 U4355 ( .QN(n3168), .IN1(n3180), .IN2(n3181) );
  NAND2X0 U4356 ( .IN1(n3182), .IN2(n3183), .QN(n3181) );
  NOR2X0 U4357 ( .QN(n3183), .IN1(P2_N299), .IN2(n3184) );
  OR2X1 U4358 ( .IN2(P2_N300), .IN1(P2_N301), .Q(n3184) );
  NOR2X0 U4359 ( .QN(n3182), .IN1(P2_N298), .IN2(P2_N297) );
  NAND2X0 U4360 ( .IN1(n3185), .IN2(n3186), .QN(n3180) );
  NOR2X0 U4361 ( .QN(n3186), .IN1(P2_N305), .IN2(n3187) );
  OR2X1 U4362 ( .IN2(P2_N306), .IN1(P2_N307), .Q(n3187) );
  NOR2X0 U4363 ( .QN(n3185), .IN1(P2_N302), .IN2(n3188) );
  OR2X1 U4364 ( .IN2(P2_N303), .IN1(P2_N304), .Q(n3188) );
  NOR2X0 U4365 ( .QN(P2_N3380), .IN1(n7329), .IN2(n7007) );
  NOR2X0 U4366 ( .QN(P2_N3379), .IN1(n7327), .IN2(n7007) );
  NOR2X0 U4367 ( .QN(P2_N3378), .IN1(n7325), .IN2(n7007) );
  NOR2X0 U4368 ( .QN(P2_N3377), .IN1(n7323), .IN2(n7011) );
  NOR2X0 U4369 ( .QN(P2_N3376), .IN1(n7321), .IN2(n7011) );
  NOR2X0 U4370 ( .QN(P2_N3375), .IN1(n7319), .IN2(n7011) );
  NOR2X0 U4371 ( .QN(P2_N3374), .IN1(n7317), .IN2(n7011) );
  NOR2X0 U4372 ( .QN(P2_N3373), .IN1(n7315), .IN2(n7015) );
  NOR2X0 U4373 ( .QN(P2_N3372), .IN1(n7313), .IN2(n7015) );
  NOR2X0 U4374 ( .QN(P2_N3371), .IN1(n7311), .IN2(n7011) );
  NAND2X0 U4376 ( .IN1(n2006), .IN2(n3190), .QN(P2_N3370) );
  NAND2X0 U4377 ( .IN1(n7012), .IN2(n2008), .QN(n3190) );
  NAND2X0 U4378 ( .IN1(n2009), .IN2(n3191), .QN(P2_N3369) );
  NAND2X0 U4379 ( .IN1(n7012), .IN2(n2011), .QN(n3191) );
  NAND2X0 U4380 ( .IN1(n2012), .IN2(n3192), .QN(P2_N3368) );
  NAND2X0 U4381 ( .IN1(n7012), .IN2(n2014), .QN(n3192) );
  NAND2X0 U4382 ( .IN1(n2015), .IN2(n3193), .QN(P2_N3367) );
  NAND2X0 U4383 ( .IN1(n7012), .IN2(n2017), .QN(n3193) );
  NAND2X0 U4384 ( .IN1(n2018), .IN2(n3194), .QN(P2_N3366) );
  NAND2X0 U4385 ( .IN1(n7009), .IN2(n2020), .QN(n3194) );
  NAND2X0 U4386 ( .IN1(n2021), .IN2(n3195), .QN(P2_N3365) );
  NAND2X0 U4387 ( .IN1(n7009), .IN2(n2023), .QN(n3195) );
  NAND2X0 U4388 ( .IN1(n2024), .IN2(n3196), .QN(P2_N3364) );
  NAND2X0 U4389 ( .IN1(n7009), .IN2(n2026), .QN(n3196) );
  NAND2X0 U4390 ( .IN1(n2027), .IN2(n3197), .QN(P2_N3363) );
  NAND2X0 U4391 ( .IN1(n7009), .IN2(n2029), .QN(n3197) );
  NAND2X0 U4392 ( .IN1(n2030), .IN2(n3198), .QN(P2_N3362) );
  NAND2X0 U4393 ( .IN1(n7010), .IN2(n2032), .QN(n3198) );
  NAND2X0 U4394 ( .IN1(n2033), .IN2(n3199), .QN(P2_N3361) );
  NAND2X0 U4395 ( .IN1(n7010), .IN2(n2035), .QN(n3199) );
  NAND2X0 U4396 ( .IN1(n2036), .IN2(n3200), .QN(P2_N3360) );
  NAND2X0 U4397 ( .IN1(n7016), .IN2(n2038), .QN(n3200) );
  NAND2X0 U4398 ( .IN1(n2039), .IN2(n3201), .QN(P2_N3359) );
  NAND2X0 U4399 ( .IN1(n7016), .IN2(n2041), .QN(n3201) );
  NAND2X0 U4400 ( .IN1(n2042), .IN2(n3202), .QN(P2_N3358) );
  NAND2X0 U4401 ( .IN1(n7016), .IN2(n2044), .QN(n3202) );
  NAND2X0 U4402 ( .IN1(n2045), .IN2(n3203), .QN(P2_N3357) );
  NAND2X0 U4403 ( .IN1(n7016), .IN2(n2047), .QN(n3203) );
  NAND2X0 U4404 ( .IN1(n2048), .IN2(n3204), .QN(P2_N3356) );
  NAND2X0 U4405 ( .IN1(n7016), .IN2(n2050), .QN(n3204) );
  NAND2X0 U4406 ( .IN1(n2051), .IN2(n3205), .QN(P2_N3355) );
  NAND2X0 U4407 ( .IN1(n7006), .IN2(n2053), .QN(n3205) );
  NAND2X0 U4214 ( .IN1(n2024), .IN2(n3088), .QN(P2_N3737) );
  NAND2X0 U4215 ( .IN1(n7009), .IN2(n2026), .QN(n3088) );
  NAND2X0 U4216 ( .IN1(n2027), .IN2(n3089), .QN(P2_N3736) );
  NAND2X0 U4217 ( .IN1(n7010), .IN2(n2029), .QN(n3089) );
  NAND2X0 U4218 ( .IN1(n2030), .IN2(n3090), .QN(P2_N3735) );
  NAND2X0 U4219 ( .IN1(n7010), .IN2(n2032), .QN(n3090) );
  NAND2X0 U4220 ( .IN1(n2033), .IN2(n3091), .QN(P2_N3734) );
  NAND2X0 U4221 ( .IN1(n7010), .IN2(n2035), .QN(n3091) );
  NAND2X0 U4222 ( .IN1(n2036), .IN2(n3092), .QN(P2_N3733) );
  NAND2X0 U4223 ( .IN1(n7016), .IN2(n2038), .QN(n3092) );
  NAND2X0 U4224 ( .IN1(n2039), .IN2(n3093), .QN(P2_N3732) );
  NAND2X0 U4225 ( .IN1(n7016), .IN2(n2041), .QN(n3093) );
  NAND2X0 U4226 ( .IN1(n2042), .IN2(n3094), .QN(P2_N3731) );
  NAND2X0 U4227 ( .IN1(n7016), .IN2(n2044), .QN(n3094) );
  NAND2X0 U4228 ( .IN1(n2045), .IN2(n3095), .QN(P2_N3730) );
  NAND2X0 U4229 ( .IN1(n7016), .IN2(n2047), .QN(n3095) );
  NAND2X0 U4230 ( .IN1(n2048), .IN2(n3096), .QN(P2_N3729) );
  NAND2X0 U4231 ( .IN1(n7016), .IN2(n2050), .QN(n3096) );
  NAND2X0 U4232 ( .IN1(n2051), .IN2(n3097), .QN(P2_N3728) );
  NAND2X0 U4233 ( .IN1(n7006), .IN2(n2053), .QN(n3097) );
  NAND2X0 U4234 ( .IN1(n2054), .IN2(n3098), .QN(P2_N3727) );
  NAND2X0 U4235 ( .IN1(n7006), .IN2(n2056), .QN(n3098) );
  NAND2X0 U4236 ( .IN1(n2057), .IN2(n3099), .QN(P2_N3726) );
  NAND2X0 U4237 ( .IN1(n7006), .IN2(n2059), .QN(n3099) );
  NAND2X0 U4238 ( .IN1(n2060), .IN2(n3100), .QN(P2_N3725) );
  NAND2X0 U4239 ( .IN1(n7006), .IN2(n2062), .QN(n3100) );
  NAND2X0 U4240 ( .IN1(n2063), .IN2(n3101), .QN(P2_N3724) );
  NAND2X0 U4241 ( .IN1(n7006), .IN2(n2065), .QN(n3101) );
  NAND2X0 U4244 ( .IN1(n3103), .IN2(n3104), .QN(P2_N3680) );
  NAND2X0 U4245 ( .IN1(P2_N3621), .IN2(n3105), .QN(n3104) );
  NAND2X0 U4246 ( .IN1(P2_N392), .IN2(P2_N5507), .QN(n3103) );
  NAND2X0 U4247 ( .IN1(n3107), .IN2(n3108), .QN(P2_N3679) );
  NAND2X0 U4248 ( .IN1(P2_N3620), .IN2(n3105), .QN(n3108) );
  NAND2X0 U4249 ( .IN1(P2_N391), .IN2(P2_N5507), .QN(n3107) );
  NAND2X0 U4250 ( .IN1(n3109), .IN2(n3110), .QN(P2_N3678) );
  NAND2X0 U4251 ( .IN1(P2_N3619), .IN2(n3105), .QN(n3110) );
  NAND2X0 U4252 ( .IN1(P2_N390), .IN2(P2_N5507), .QN(n3109) );
  NAND2X0 U4253 ( .IN1(n3111), .IN2(n3112), .QN(P2_N3677) );
  NAND2X0 U4254 ( .IN1(P2_N3618), .IN2(n3105), .QN(n3112) );
  NAND2X0 U4255 ( .IN1(P2_N389), .IN2(P2_N5507), .QN(n3111) );
  NAND2X0 U4256 ( .IN1(n3113), .IN2(n3114), .QN(P2_N3676) );
  NAND2X0 U4257 ( .IN1(P2_N3617), .IN2(n3105), .QN(n3114) );
  NAND2X0 U4258 ( .IN1(P2_N388), .IN2(P2_N5507), .QN(n3113) );
  NAND2X0 U4259 ( .IN1(n3115), .IN2(n3116), .QN(P2_N3675) );
  NAND2X0 U4260 ( .IN1(P2_N3616), .IN2(n3105), .QN(n3116) );
  NAND2X0 U4261 ( .IN1(P2_N387), .IN2(P2_N5507), .QN(n3115) );
  NAND2X0 U4262 ( .IN1(n3117), .IN2(n3118), .QN(P2_N3674) );
  NAND2X0 U4263 ( .IN1(P2_N3615), .IN2(n3105), .QN(n3118) );
  NAND2X0 U4264 ( .IN1(P2_N386), .IN2(P2_N5507), .QN(n3117) );
  NAND2X0 U4265 ( .IN1(n3119), .IN2(n3120), .QN(P2_N3673) );
  NAND2X0 U4266 ( .IN1(P2_N3614), .IN2(n3105), .QN(n3120) );
  NAND2X0 U4267 ( .IN1(P2_N385), .IN2(P2_N5507), .QN(n3119) );
  NAND2X0 U4268 ( .IN1(n3121), .IN2(n3122), .QN(P2_N3672) );
  NAND2X0 U4269 ( .IN1(P2_N3613), .IN2(n3105), .QN(n3122) );
  NAND2X0 U4270 ( .IN1(P2_N384), .IN2(P2_N5507), .QN(n3121) );
  NAND2X0 U4271 ( .IN1(n3123), .IN2(n3124), .QN(P2_N3671) );
  NAND2X0 U4272 ( .IN1(P2_N3612), .IN2(n3105), .QN(n3124) );
  NAND2X0 U4273 ( .IN1(P2_N383), .IN2(P2_N5507), .QN(n3123) );
  NAND2X0 U4274 ( .IN1(n3125), .IN2(n3126), .QN(P2_N3670) );
  NAND2X0 U4275 ( .IN1(P2_N3611), .IN2(n3105), .QN(n3126) );
  NAND2X0 U4276 ( .IN1(P2_N382), .IN2(P2_N5507), .QN(n3125) );
  NAND2X0 U4277 ( .IN1(n3127), .IN2(n3128), .QN(P2_N3669) );
  NAND2X0 U4278 ( .IN1(P2_N3610), .IN2(n3105), .QN(n3128) );
  NAND2X0 U4279 ( .IN1(P2_N381), .IN2(P2_N5507), .QN(n3127) );
  NAND2X0 U4280 ( .IN1(n3129), .IN2(n3130), .QN(P2_N3668) );
  NAND2X0 U4281 ( .IN1(P2_N3609), .IN2(n3105), .QN(n3130) );
  NAND2X0 U4282 ( .IN1(P2_N380), .IN2(P2_N5507), .QN(n3129) );
  NAND2X0 U4283 ( .IN1(n3131), .IN2(n3132), .QN(P2_N3667) );
  NAND2X0 U4284 ( .IN1(P2_N3608), .IN2(n3105), .QN(n3132) );
  NAND2X0 U4285 ( .IN1(P2_N379), .IN2(P2_N5507), .QN(n3131) );
  NAND2X0 U4286 ( .IN1(n3133), .IN2(n3134), .QN(P2_N3666) );
  NAND2X0 U4287 ( .IN1(P2_N3607), .IN2(n3105), .QN(n3134) );
  NAND2X0 U4288 ( .IN1(P2_N378), .IN2(P2_N5507), .QN(n3133) );
  NAND2X0 U4289 ( .IN1(n3135), .IN2(n3136), .QN(P2_N3665) );
  NAND2X0 U4290 ( .IN1(P2_N3606), .IN2(n3105), .QN(n3136) );
  NAND2X0 U4291 ( .IN1(P2_N377), .IN2(P2_N5507), .QN(n3135) );
  NAND2X0 U4292 ( .IN1(n3137), .IN2(n3138), .QN(P2_N3664) );
  NAND2X0 U4293 ( .IN1(P2_N3605), .IN2(n3105), .QN(n3138) );
  NAND2X0 U4294 ( .IN1(P2_N376), .IN2(P2_N5507), .QN(n3137) );
  NAND2X0 U4295 ( .IN1(n3139), .IN2(n3140), .QN(P2_N3663) );
  NAND2X0 U4296 ( .IN1(P2_N3604), .IN2(n3105), .QN(n3140) );
  NAND2X0 U4297 ( .IN1(P2_N375), .IN2(P2_N5507), .QN(n3139) );
  NAND2X0 U4298 ( .IN1(n3141), .IN2(n3142), .QN(P2_N3662) );
  NAND2X0 U4299 ( .IN1(P2_N3603), .IN2(n3105), .QN(n3142) );
  NAND2X0 U4300 ( .IN1(P2_N374), .IN2(P2_N5507), .QN(n3141) );
  NAND2X0 U4301 ( .IN1(n3143), .IN2(n3144), .QN(P2_N3661) );
  NAND2X0 U4302 ( .IN1(P2_N3602), .IN2(n3105), .QN(n3144) );
  NAND2X0 U4303 ( .IN1(P2_N373), .IN2(P2_N5507), .QN(n3143) );
  NAND2X0 U4304 ( .IN1(n3145), .IN2(n3146), .QN(P2_N3660) );
  NAND2X0 U4305 ( .IN1(P2_N3601), .IN2(n3105), .QN(n3146) );
  NAND2X0 U4306 ( .IN1(P2_N372), .IN2(P2_N5507), .QN(n3145) );
  NAND2X0 U4307 ( .IN1(n3147), .IN2(n3148), .QN(P2_N3659) );
  NAND2X0 U4308 ( .IN1(P2_N3600), .IN2(n3105), .QN(n3148) );
  NAND2X0 U4115 ( .IN1(P2_N3987), .IN2(n3019), .QN(n3034) );
  NAND2X0 U4116 ( .IN1(P2_N385), .IN2(P2_N5508), .QN(n3033) );
  NAND2X0 U4117 ( .IN1(n3035), .IN2(n3036), .QN(P2_N4045) );
  NAND2X0 U4118 ( .IN1(P2_N3986), .IN2(n3019), .QN(n3036) );
  NAND2X0 U4119 ( .IN1(P2_N384), .IN2(P2_N5508), .QN(n3035) );
  NAND2X0 U4120 ( .IN1(n3037), .IN2(n3038), .QN(P2_N4044) );
  NAND2X0 U4121 ( .IN1(P2_N3985), .IN2(n3019), .QN(n3038) );
  NAND2X0 U4122 ( .IN1(P2_N383), .IN2(P2_N5508), .QN(n3037) );
  NAND2X0 U4123 ( .IN1(n3039), .IN2(n3040), .QN(P2_N4043) );
  NAND2X0 U4124 ( .IN1(P2_N3984), .IN2(n3019), .QN(n3040) );
  NAND2X0 U4125 ( .IN1(P2_N382), .IN2(P2_N5508), .QN(n3039) );
  NAND2X0 U4126 ( .IN1(n3041), .IN2(n3042), .QN(P2_N4042) );
  NAND2X0 U4127 ( .IN1(P2_N3983), .IN2(n3019), .QN(n3042) );
  NAND2X0 U4128 ( .IN1(P2_N381), .IN2(P2_N5508), .QN(n3041) );
  NAND2X0 U4129 ( .IN1(n3043), .IN2(n3044), .QN(P2_N4041) );
  NAND2X0 U4130 ( .IN1(P2_N3982), .IN2(n3019), .QN(n3044) );
  NAND2X0 U4131 ( .IN1(P2_N380), .IN2(P2_N5508), .QN(n3043) );
  NAND2X0 U4132 ( .IN1(n3045), .IN2(n3046), .QN(P2_N4040) );
  NAND2X0 U4133 ( .IN1(P2_N3981), .IN2(n3019), .QN(n3046) );
  NAND2X0 U4134 ( .IN1(P2_N379), .IN2(P2_N5508), .QN(n3045) );
  NAND2X0 U4135 ( .IN1(n3047), .IN2(n3048), .QN(P2_N4039) );
  NAND2X0 U4136 ( .IN1(P2_N3980), .IN2(n3019), .QN(n3048) );
  NAND2X0 U4137 ( .IN1(P2_N378), .IN2(P2_N5508), .QN(n3047) );
  NAND2X0 U4138 ( .IN1(n3049), .IN2(n3050), .QN(P2_N4038) );
  NAND2X0 U4139 ( .IN1(P2_N3979), .IN2(n3019), .QN(n3050) );
  NAND2X0 U4140 ( .IN1(P2_N377), .IN2(P2_N5508), .QN(n3049) );
  NAND2X0 U4141 ( .IN1(n3051), .IN2(n3052), .QN(P2_N4037) );
  NAND2X0 U4142 ( .IN1(P2_N3978), .IN2(n3019), .QN(n3052) );
  NAND2X0 U4143 ( .IN1(P2_N376), .IN2(P2_N5508), .QN(n3051) );
  NAND2X0 U4144 ( .IN1(n3053), .IN2(n3054), .QN(P2_N4036) );
  NAND2X0 U4145 ( .IN1(P2_N3977), .IN2(n3019), .QN(n3054) );
  NAND2X0 U4146 ( .IN1(P2_N375), .IN2(P2_N5508), .QN(n3053) );
  NAND2X0 U4147 ( .IN1(n3055), .IN2(n3056), .QN(P2_N4035) );
  NAND2X0 U4148 ( .IN1(P2_N3976), .IN2(n3019), .QN(n3056) );
  NAND2X0 U4149 ( .IN1(P2_N374), .IN2(P2_N5508), .QN(n3055) );
  NAND2X0 U4150 ( .IN1(n3057), .IN2(n3058), .QN(P2_N4034) );
  NAND2X0 U4151 ( .IN1(P2_N3975), .IN2(n3019), .QN(n3058) );
  NAND2X0 U4152 ( .IN1(P2_N373), .IN2(P2_N5508), .QN(n3057) );
  NAND2X0 U4153 ( .IN1(n3059), .IN2(n3060), .QN(P2_N4033) );
  NAND2X0 U4154 ( .IN1(P2_N3974), .IN2(n3019), .QN(n3060) );
  NAND2X0 U4155 ( .IN1(P2_N372), .IN2(P2_N5508), .QN(n3059) );
  NAND2X0 U4156 ( .IN1(n3061), .IN2(n3062), .QN(P2_N4032) );
  NAND2X0 U4157 ( .IN1(P2_N3973), .IN2(n3019), .QN(n3062) );
  NAND2X0 U4158 ( .IN1(P2_N371), .IN2(P2_N5508), .QN(n3061) );
  NAND2X0 U4159 ( .IN1(n3063), .IN2(n3064), .QN(P2_N4031) );
  NAND2X0 U4160 ( .IN1(P2_N3972), .IN2(n3019), .QN(n3064) );
  NAND2X0 U4161 ( .IN1(P2_N370), .IN2(P2_N5508), .QN(n3063) );
  NAND2X0 U4162 ( .IN1(n3065), .IN2(n3066), .QN(P2_N4030) );
  NAND2X0 U4163 ( .IN1(P2_N3971), .IN2(n3019), .QN(n3066) );
  NAND2X0 U4164 ( .IN1(P2_N369), .IN2(P2_N5508), .QN(n3065) );
  NAND2X0 U4165 ( .IN1(n3067), .IN2(n3068), .QN(P2_N4029) );
  NAND2X0 U4166 ( .IN1(P2_N3970), .IN2(n3019), .QN(n3068) );
  NAND2X0 U4167 ( .IN1(P2_N368), .IN2(P2_N5508), .QN(n3067) );
  NAND2X0 U4168 ( .IN1(n3069), .IN2(n3070), .QN(P2_N4028) );
  NAND2X0 U4169 ( .IN1(P2_N3969), .IN2(n3019), .QN(n3070) );
  NAND2X0 U4170 ( .IN1(n18813), .IN2(P2_N5508), .QN(n3069) );
  NAND2X0 U4171 ( .IN1(n3071), .IN2(n3072), .QN(P2_N4027) );
  NAND2X0 U4172 ( .IN1(P2_N3968), .IN2(n3019), .QN(n3072) );
  NAND2X0 U4173 ( .IN1(n6683), .IN2(P2_N5508), .QN(n3071) );
  NAND2X0 U4174 ( .IN1(n3073), .IN2(n3074), .QN(P2_N4026) );
  NAND2X0 U4175 ( .IN1(P2_N3967), .IN2(n3019), .QN(n3074) );
  NAND2X0 U4176 ( .IN1(n6682), .IN2(P2_N5508), .QN(n3073) );
  NAND2X0 U4177 ( .IN1(n3075), .IN2(n3076), .QN(P2_N4025) );
  NAND2X0 U4178 ( .IN1(P2_N3966), .IN2(n3019), .QN(n3076) );
  NAND2X0 U4181 ( .IN1(n6681), .IN2(P2_N5508), .QN(n3075) );
  NAND2X0 U4186 ( .IN1(n7394), .IN2(n3079), .QN(P2_N3873) );
  NAND2X0 U4187 ( .IN1(n7393), .IN2(n3080), .QN(P2_N3871) );
  NOR2X0 U4188 ( .QN(P2_N4054), .IN1(n3080), .IN2(n3079) );
  INVX0 U4189 ( .ZN(n3079), .INP(n7393) );
  INVX0 U4190 ( .ZN(n3080), .INP(n7394) );
  NOR2X0 U4191 ( .QN(P2_N3753), .IN1(n7329), .IN2(n7007) );
  NOR2X0 U4192 ( .QN(P2_N3752), .IN1(n7327), .IN2(n7007) );
  NOR2X0 U4193 ( .QN(P2_N3751), .IN1(n7325), .IN2(n7007) );
  NOR2X0 U4194 ( .QN(P2_N3750), .IN1(n7323), .IN2(n7011) );
  NOR2X0 U4195 ( .QN(P2_N3749), .IN1(n7321), .IN2(n7011) );
  NOR2X0 U4196 ( .QN(P2_N3748), .IN1(n7319), .IN2(n7011) );
  NOR2X0 U4197 ( .QN(P2_N3747), .IN1(n7317), .IN2(n7011) );
  NOR2X0 U4198 ( .QN(P2_N3746), .IN1(n7315), .IN2(n7015) );
  NOR2X0 U4199 ( .QN(P2_N3745), .IN1(n7313), .IN2(n7015) );
  NOR2X0 U4200 ( .QN(P2_N3744), .IN1(n7311), .IN2(n7015) );
  NAND2X0 U4202 ( .IN1(n2006), .IN2(n3082), .QN(P2_N3743) );
  NAND2X0 U4203 ( .IN1(P2_N914), .IN2(n2008), .QN(n3082) );
  NAND2X0 U4204 ( .IN1(n2009), .IN2(n3083), .QN(P2_N3742) );
  NAND2X0 U4205 ( .IN1(P2_N914), .IN2(n2011), .QN(n3083) );
  NAND2X0 U4206 ( .IN1(n2012), .IN2(n3084), .QN(P2_N3741) );
  NAND2X0 U4207 ( .IN1(P2_N914), .IN2(n2014), .QN(n3084) );
  NAND2X0 U4208 ( .IN1(n2015), .IN2(n3085), .QN(P2_N3740) );
  NAND2X0 U4209 ( .IN1(P2_N914), .IN2(n2017), .QN(n3085) );
  NAND2X0 U4210 ( .IN1(n2018), .IN2(n3086), .QN(P2_N3739) );
  NAND2X0 U4211 ( .IN1(n7009), .IN2(n2020), .QN(n3086) );
  NAND2X0 U4212 ( .IN1(n2021), .IN2(n3087), .QN(P2_N3738) );
  NAND2X0 U4213 ( .IN1(n7009), .IN2(n2023), .QN(n3087) );
  NAND2X0 U4013 ( .IN1(P2_N369), .IN2(P2_N5509), .QN(n2980) );
  NAND2X0 U4014 ( .IN1(n2982), .IN2(n2983), .QN(P2_N4403) );
  NAND2X0 U4015 ( .IN1(P2_N4253), .IN2(n2934), .QN(n2983) );
  NAND2X0 U4016 ( .IN1(P2_N368), .IN2(P2_N5509), .QN(n2982) );
  NAND2X0 U4017 ( .IN1(n2984), .IN2(n2985), .QN(P2_N4402) );
  NAND2X0 U4018 ( .IN1(P2_N4252), .IN2(n2934), .QN(n2985) );
  NAND2X0 U4019 ( .IN1(n18813), .IN2(P2_N5509), .QN(n2984) );
  NAND2X0 U4020 ( .IN1(n2986), .IN2(n2987), .QN(P2_N4401) );
  NAND2X0 U4021 ( .IN1(P2_N4251), .IN2(n2934), .QN(n2987) );
  NAND2X0 U4022 ( .IN1(n6683), .IN2(P2_N5509), .QN(n2986) );
  NAND2X0 U4023 ( .IN1(n2988), .IN2(n2989), .QN(P2_N4400) );
  NAND2X0 U4024 ( .IN1(P2_N4250), .IN2(n2934), .QN(n2989) );
  NAND2X0 U4025 ( .IN1(n6682), .IN2(P2_N5509), .QN(n2988) );
  NAND2X0 U4026 ( .IN1(n2990), .IN2(n2991), .QN(P2_N4399) );
  NAND2X0 U4027 ( .IN1(P2_N4249), .IN2(n2934), .QN(n2991) );
  NAND2X0 U4030 ( .IN1(n6681), .IN2(P2_N5509), .QN(n2990) );
  NOR2X0 U4036 ( .QN(P2_N4398), .IN1(n2992), .IN2(n7354) );
  OR2X1 U4038 ( .IN2(n7354), .IN1(P2_N4178), .Q(P2_N4244) );
  NOR2X0 U4040 ( .QN(P2_N4126), .IN1(n7329), .IN2(n7007) );
  NOR2X0 U4041 ( .QN(P2_N4125), .IN1(n7327), .IN2(n7007) );
  NOR2X0 U4042 ( .QN(P2_N4124), .IN1(n7325), .IN2(n7007) );
  NOR2X0 U4043 ( .QN(P2_N4123), .IN1(n7323), .IN2(n7011) );
  NOR2X0 U4044 ( .QN(P2_N4122), .IN1(n7321), .IN2(n7011) );
  NOR2X0 U4045 ( .QN(P2_N4121), .IN1(n7319), .IN2(n7011) );
  NOR2X0 U4046 ( .QN(P2_N4120), .IN1(n7317), .IN2(n7011) );
  NOR2X0 U4047 ( .QN(P2_N4119), .IN1(n7315), .IN2(n7015) );
  NOR2X0 U4048 ( .QN(P2_N4118), .IN1(n7313), .IN2(n7015) );
  NOR2X0 U4049 ( .QN(P2_N4117), .IN1(n7311), .IN2(n7015) );
  NAND2X0 U4051 ( .IN1(n2006), .IN2(n2996), .QN(P2_N4116) );
  NAND2X0 U4052 ( .IN1(P2_N914), .IN2(n2008), .QN(n2996) );
  NAND2X0 U4053 ( .IN1(n2009), .IN2(n2997), .QN(P2_N4115) );
  NAND2X0 U4054 ( .IN1(P2_N914), .IN2(n2011), .QN(n2997) );
  NAND2X0 U4055 ( .IN1(n2012), .IN2(n2998), .QN(P2_N4114) );
  NAND2X0 U4056 ( .IN1(P2_N914), .IN2(n2014), .QN(n2998) );
  NAND2X0 U4057 ( .IN1(n2015), .IN2(n2999), .QN(P2_N4113) );
  NAND2X0 U4058 ( .IN1(P2_N914), .IN2(n2017), .QN(n2999) );
  NAND2X0 U4059 ( .IN1(n2018), .IN2(n3000), .QN(P2_N4112) );
  NAND2X0 U4060 ( .IN1(n7009), .IN2(n2020), .QN(n3000) );
  NAND2X0 U4061 ( .IN1(n2021), .IN2(n3001), .QN(P2_N4111) );
  NAND2X0 U4062 ( .IN1(n7009), .IN2(n2023), .QN(n3001) );
  NAND2X0 U4063 ( .IN1(n2024), .IN2(n3002), .QN(P2_N4110) );
  NAND2X0 U4064 ( .IN1(n7009), .IN2(n2026), .QN(n3002) );
  NAND2X0 U4065 ( .IN1(n2027), .IN2(n3003), .QN(P2_N4109) );
  NAND2X0 U4066 ( .IN1(n7009), .IN2(n2029), .QN(n3003) );
  NAND2X0 U4067 ( .IN1(n2030), .IN2(n3004), .QN(P2_N4108) );
  NAND2X0 U4068 ( .IN1(n7010), .IN2(n2032), .QN(n3004) );
  NAND2X0 U4069 ( .IN1(n2033), .IN2(n3005), .QN(P2_N4107) );
  NAND2X0 U4070 ( .IN1(n7010), .IN2(n2035), .QN(n3005) );
  NAND2X0 U4071 ( .IN1(n2036), .IN2(n3006), .QN(P2_N4106) );
  NAND2X0 U4072 ( .IN1(n7016), .IN2(n2038), .QN(n3006) );
  NAND2X0 U4073 ( .IN1(n2039), .IN2(n3007), .QN(P2_N4105) );
  NAND2X0 U4074 ( .IN1(n7016), .IN2(n2041), .QN(n3007) );
  NAND2X0 U4075 ( .IN1(n2042), .IN2(n3008), .QN(P2_N4104) );
  NAND2X0 U4076 ( .IN1(n7016), .IN2(n2044), .QN(n3008) );
  NAND2X0 U4077 ( .IN1(n2045), .IN2(n3009), .QN(P2_N4103) );
  NAND2X0 U4078 ( .IN1(n7016), .IN2(n2047), .QN(n3009) );
  NAND2X0 U4079 ( .IN1(n2048), .IN2(n3010), .QN(P2_N4102) );
  NAND2X0 U4080 ( .IN1(n7016), .IN2(n2050), .QN(n3010) );
  NAND2X0 U4081 ( .IN1(n2051), .IN2(n3011), .QN(P2_N4101) );
  NAND2X0 U4082 ( .IN1(n7006), .IN2(n2053), .QN(n3011) );
  NAND2X0 U4083 ( .IN1(n2054), .IN2(n3012), .QN(P2_N4100) );
  NAND2X0 U4084 ( .IN1(n7006), .IN2(n2056), .QN(n3012) );
  NAND2X0 U4085 ( .IN1(n2057), .IN2(n3013), .QN(P2_N4099) );
  NAND2X0 U4086 ( .IN1(n7462), .IN2(n2059), .QN(n3013) );
  NAND2X0 U4087 ( .IN1(n2060), .IN2(n3014), .QN(P2_N4098) );
  NAND2X0 U4088 ( .IN1(n7462), .IN2(n2062), .QN(n3014) );
  NAND2X0 U4089 ( .IN1(n2063), .IN2(n3015), .QN(P2_N4097) );
  NAND2X0 U4090 ( .IN1(n7462), .IN2(n2065), .QN(n3015) );
  NAND2X0 U4093 ( .IN1(n3017), .IN2(n3018), .QN(P2_N4053) );
  NAND2X0 U4094 ( .IN1(P2_N3994), .IN2(n3019), .QN(n3018) );
  NAND2X0 U4095 ( .IN1(P2_N392), .IN2(P2_N5508), .QN(n3017) );
  NAND2X0 U4096 ( .IN1(n3021), .IN2(n3022), .QN(P2_N4052) );
  NAND2X0 U4097 ( .IN1(P2_N3993), .IN2(n3019), .QN(n3022) );
  NAND2X0 U4098 ( .IN1(P2_N391), .IN2(P2_N5508), .QN(n3021) );
  NAND2X0 U4099 ( .IN1(n3023), .IN2(n3024), .QN(P2_N4051) );
  NAND2X0 U4100 ( .IN1(P2_N3992), .IN2(n3019), .QN(n3024) );
  NAND2X0 U4101 ( .IN1(P2_N390), .IN2(P2_N5508), .QN(n3023) );
  NAND2X0 U4102 ( .IN1(n3025), .IN2(n3026), .QN(P2_N4050) );
  NAND2X0 U4103 ( .IN1(P2_N3991), .IN2(n3019), .QN(n3026) );
  NAND2X0 U4104 ( .IN1(P2_N389), .IN2(P2_N5508), .QN(n3025) );
  NAND2X0 U4105 ( .IN1(n3027), .IN2(n3028), .QN(P2_N4049) );
  NAND2X0 U4106 ( .IN1(P2_N3990), .IN2(n3019), .QN(n3028) );
  NAND2X0 U4107 ( .IN1(P2_N388), .IN2(P2_N5508), .QN(n3027) );
  NAND2X0 U4108 ( .IN1(n3029), .IN2(n3030), .QN(P2_N4048) );
  NAND2X0 U4109 ( .IN1(P2_N3989), .IN2(n3019), .QN(n3030) );
  NAND2X0 U4110 ( .IN1(P2_N387), .IN2(P2_N5508), .QN(n3029) );
  NAND2X0 U4111 ( .IN1(n3031), .IN2(n3032), .QN(P2_N4047) );
  NAND2X0 U4112 ( .IN1(P2_N3988), .IN2(n3019), .QN(n3032) );
  NAND2X0 U4113 ( .IN1(P2_N386), .IN2(P2_N5508), .QN(n3031) );
  NAND2X0 U4114 ( .IN1(n3033), .IN2(n3034), .QN(P2_N4046) );
  NAND2X0 U3919 ( .IN1(P2_N5493), .IN2(n7035), .QN(n2917) );
  AND2X1 U3921 ( .IN1(P2_N4431), .IN2(n2702), .Q(P2_N4499) );
  OR2X1 U3922 ( .IN2(n2693), .IN1(n7341), .Q(n2702) );
  NOR2X0 U3923 ( .QN(P2_N4430), .IN1(n2562), .IN2(n2919) );
  NAND2X0 U3925 ( .IN1(n2922), .IN2(n2923), .QN(n2921) );
  NAND2X0 U3926 ( .IN1(n9837), .IN2(n7342), .QN(n2923) );
  NAND2X0 U3927 ( .IN1(n9842), .IN2(n7343), .QN(n2922) );
  NAND2X0 U3928 ( .IN1(n2924), .IN2(n2925), .QN(n2920) );
  NAND2X0 U3929 ( .IN1(n9218), .IN2(n2569), .QN(n2925) );
  NAND2X0 U3930 ( .IN1(n7346), .IN2(n6681), .QN(n2924) );
  NOR2X0 U3931 ( .QN(n2562), .IN1(n2926), .IN2(n2927) );
  NAND2X0 U3932 ( .IN1(n2928), .IN2(n2929), .QN(n2927) );
  NAND2X0 U3933 ( .IN1(n9222), .IN2(n7342), .QN(n2929) );
  NAND2X0 U3934 ( .IN1(n9306), .IN2(n7343), .QN(n2928) );
  NAND2X0 U3935 ( .IN1(n2567), .IN2(n2930), .QN(n2926) );
  NAND2X0 U3936 ( .IN1(n9098), .IN2(n2569), .QN(n2930) );
  INVX0 U3938 ( .ZN(n2661), .INP(n7338) );
  INVX0 U3939 ( .ZN(n2660), .INP(n7339) );
  NAND2X0 U3940 ( .IN1(n7346), .IN2(P2_N394), .QN(n2567) );
  NAND2X0 U3942 ( .IN1(n2932), .IN2(n2933), .QN(P2_N4427) );
  NAND2X0 U3943 ( .IN1(P2_N4277), .IN2(n2934), .QN(n2933) );
  NAND2X0 U3944 ( .IN1(P2_N392), .IN2(P2_N5509), .QN(n2932) );
  NAND2X0 U3945 ( .IN1(n2936), .IN2(n2937), .QN(P2_N4426) );
  NAND2X0 U3946 ( .IN1(P2_N4276), .IN2(n2934), .QN(n2937) );
  NAND2X0 U3947 ( .IN1(P2_N391), .IN2(P2_N5509), .QN(n2936) );
  NAND2X0 U3948 ( .IN1(n2938), .IN2(n2939), .QN(P2_N4425) );
  NAND2X0 U3949 ( .IN1(P2_N4275), .IN2(n2934), .QN(n2939) );
  NAND2X0 U3950 ( .IN1(P2_N390), .IN2(P2_N5509), .QN(n2938) );
  NAND2X0 U3951 ( .IN1(n2940), .IN2(n2941), .QN(P2_N4424) );
  NAND2X0 U3952 ( .IN1(P2_N4274), .IN2(n2934), .QN(n2941) );
  NAND2X0 U3953 ( .IN1(P2_N389), .IN2(P2_N5509), .QN(n2940) );
  NAND2X0 U3954 ( .IN1(n2942), .IN2(n2943), .QN(P2_N4423) );
  NAND2X0 U3955 ( .IN1(P2_N4273), .IN2(n2934), .QN(n2943) );
  NAND2X0 U3956 ( .IN1(P2_N388), .IN2(P2_N5509), .QN(n2942) );
  NAND2X0 U3957 ( .IN1(n2944), .IN2(n2945), .QN(P2_N4422) );
  NAND2X0 U3958 ( .IN1(P2_N4272), .IN2(n2934), .QN(n2945) );
  NAND2X0 U3959 ( .IN1(P2_N387), .IN2(P2_N5509), .QN(n2944) );
  NAND2X0 U3960 ( .IN1(n2946), .IN2(n2947), .QN(P2_N4421) );
  NAND2X0 U3961 ( .IN1(P2_N4271), .IN2(n2934), .QN(n2947) );
  NAND2X0 U3962 ( .IN1(P2_N386), .IN2(P2_N5509), .QN(n2946) );
  NAND2X0 U3963 ( .IN1(n2948), .IN2(n2949), .QN(P2_N4420) );
  NAND2X0 U3964 ( .IN1(P2_N4270), .IN2(n2934), .QN(n2949) );
  NAND2X0 U3965 ( .IN1(P2_N385), .IN2(P2_N5509), .QN(n2948) );
  NAND2X0 U3966 ( .IN1(n2950), .IN2(n2951), .QN(P2_N4419) );
  NAND2X0 U3967 ( .IN1(P2_N4269), .IN2(n2934), .QN(n2951) );
  NAND2X0 U3968 ( .IN1(P2_N384), .IN2(P2_N5509), .QN(n2950) );
  NAND2X0 U3969 ( .IN1(n2952), .IN2(n2953), .QN(P2_N4418) );
  NAND2X0 U3970 ( .IN1(P2_N4268), .IN2(n2934), .QN(n2953) );
  NAND2X0 U3971 ( .IN1(P2_N383), .IN2(P2_N5509), .QN(n2952) );
  NAND2X0 U3972 ( .IN1(n2954), .IN2(n2955), .QN(P2_N4417) );
  NAND2X0 U3973 ( .IN1(P2_N4267), .IN2(n2934), .QN(n2955) );
  NAND2X0 U3974 ( .IN1(P2_N382), .IN2(P2_N5509), .QN(n2954) );
  NAND2X0 U3975 ( .IN1(n2956), .IN2(n2957), .QN(P2_N4416) );
  NAND2X0 U3976 ( .IN1(P2_N4266), .IN2(n2934), .QN(n2957) );
  NAND2X0 U3977 ( .IN1(P2_N381), .IN2(P2_N5509), .QN(n2956) );
  NAND2X0 U3978 ( .IN1(n2958), .IN2(n2959), .QN(P2_N4415) );
  NAND2X0 U3979 ( .IN1(P2_N4265), .IN2(n2934), .QN(n2959) );
  NAND2X0 U3980 ( .IN1(P2_N380), .IN2(P2_N5509), .QN(n2958) );
  NAND2X0 U3981 ( .IN1(n2960), .IN2(n2961), .QN(P2_N4414) );
  NAND2X0 U3982 ( .IN1(P2_N4264), .IN2(n2934), .QN(n2961) );
  NAND2X0 U3983 ( .IN1(P2_N379), .IN2(P2_N5509), .QN(n2960) );
  NAND2X0 U3984 ( .IN1(n2962), .IN2(n2963), .QN(P2_N4413) );
  NAND2X0 U3985 ( .IN1(P2_N4263), .IN2(n2934), .QN(n2963) );
  NAND2X0 U3986 ( .IN1(P2_N378), .IN2(P2_N5509), .QN(n2962) );
  NAND2X0 U3987 ( .IN1(n2964), .IN2(n2965), .QN(P2_N4412) );
  NAND2X0 U3988 ( .IN1(P2_N4262), .IN2(n2934), .QN(n2965) );
  NAND2X0 U3989 ( .IN1(P2_N377), .IN2(P2_N5509), .QN(n2964) );
  NAND2X0 U3990 ( .IN1(n2966), .IN2(n2967), .QN(P2_N4411) );
  NAND2X0 U3991 ( .IN1(P2_N4261), .IN2(n2934), .QN(n2967) );
  NAND2X0 U3992 ( .IN1(P2_N376), .IN2(P2_N5509), .QN(n2966) );
  NAND2X0 U3993 ( .IN1(n2968), .IN2(n2969), .QN(P2_N4410) );
  NAND2X0 U3994 ( .IN1(P2_N4260), .IN2(n2934), .QN(n2969) );
  NAND2X0 U3995 ( .IN1(P2_N375), .IN2(P2_N5509), .QN(n2968) );
  NAND2X0 U3996 ( .IN1(n2970), .IN2(n2971), .QN(P2_N4409) );
  NAND2X0 U3997 ( .IN1(P2_N4259), .IN2(n2934), .QN(n2971) );
  NAND2X0 U3998 ( .IN1(P2_N374), .IN2(P2_N5509), .QN(n2970) );
  NAND2X0 U3999 ( .IN1(n2972), .IN2(n2973), .QN(P2_N4408) );
  NAND2X0 U4000 ( .IN1(P2_N4258), .IN2(n2934), .QN(n2973) );
  NAND2X0 U4001 ( .IN1(P2_N373), .IN2(P2_N5509), .QN(n2972) );
  NAND2X0 U4002 ( .IN1(n2974), .IN2(n2975), .QN(P2_N4407) );
  NAND2X0 U4003 ( .IN1(P2_N4257), .IN2(n2934), .QN(n2975) );
  NAND2X0 U4004 ( .IN1(P2_N372), .IN2(P2_N5509), .QN(n2974) );
  NAND2X0 U4005 ( .IN1(n2976), .IN2(n2977), .QN(P2_N4406) );
  NAND2X0 U4006 ( .IN1(P2_N4256), .IN2(n2934), .QN(n2977) );
  NAND2X0 U4007 ( .IN1(P2_N371), .IN2(P2_N5509), .QN(n2976) );
  NAND2X0 U4008 ( .IN1(n2978), .IN2(n2979), .QN(P2_N4405) );
  NAND2X0 U4009 ( .IN1(P2_N4255), .IN2(n2934), .QN(n2979) );
  NAND2X0 U4010 ( .IN1(P2_N370), .IN2(P2_N5509), .QN(n2978) );
  NAND2X0 U4011 ( .IN1(n2980), .IN2(n2981), .QN(P2_N4404) );
  NAND2X0 U4012 ( .IN1(P2_N4254), .IN2(n2934), .QN(n2981) );
  NAND2X0 U3826 ( .IN1(n7346), .IN2(P2_N374), .QN(n2843) );
  NAND2X0 U3827 ( .IN1(n2845), .IN2(n2846), .QN(P2_N4509) );
  NAND2X0 U3828 ( .IN1(P2_N4441), .IN2(n2702), .QN(n2846) );
  NAND2X0 U3829 ( .IN1(P2_N5493), .IN2(P2_N5080), .QN(n2845) );
  OR2X1 U3830 ( .IN2(n2848), .IN1(n2847), .Q(P2_N5080) );
  NAND2X0 U3831 ( .IN1(n2849), .IN2(n2850), .QN(n2848) );
  NAND2X0 U3832 ( .IN1(n6671), .IN2(n7342), .QN(n2850) );
  NAND2X0 U3833 ( .IN1(n6654), .IN2(n7343), .QN(n2849) );
  NAND2X0 U3834 ( .IN1(n2851), .IN2(n2852), .QN(n2847) );
  NAND2X0 U3835 ( .IN1(n9182), .IN2(n2569), .QN(n2852) );
  NAND2X0 U3836 ( .IN1(n7346), .IN2(P2_N373), .QN(n2851) );
  NAND2X0 U3837 ( .IN1(n2853), .IN2(n2854), .QN(P2_N4508) );
  NAND2X0 U3838 ( .IN1(P2_N4440), .IN2(n2702), .QN(n2854) );
  NAND2X0 U3839 ( .IN1(P2_N5493), .IN2(n7154), .QN(n2853) );
  OR2X1 U3840 ( .IN2(n2856), .IN1(n2855), .Q(P2_N5079) );
  NAND2X0 U3841 ( .IN1(n2857), .IN2(n2858), .QN(n2856) );
  NAND2X0 U3842 ( .IN1(n10249), .IN2(n7342), .QN(n2858) );
  NAND2X0 U3843 ( .IN1(n6653), .IN2(n7343), .QN(n2857) );
  NAND2X0 U3844 ( .IN1(n2859), .IN2(n2860), .QN(n2855) );
  NAND2X0 U3845 ( .IN1(n9186), .IN2(n2569), .QN(n2860) );
  NAND2X0 U3846 ( .IN1(n7346), .IN2(P2_N372), .QN(n2859) );
  NAND2X0 U3847 ( .IN1(n2861), .IN2(n2862), .QN(P2_N4507) );
  NAND2X0 U3848 ( .IN1(P2_N4439), .IN2(n2702), .QN(n2862) );
  NAND2X0 U3849 ( .IN1(P2_N5493), .IN2(n7158), .QN(n2861) );
  OR2X1 U3850 ( .IN2(n2864), .IN1(n2863), .Q(P2_N5078) );
  NAND2X0 U3851 ( .IN1(n2865), .IN2(n2866), .QN(n2864) );
  NAND2X0 U3852 ( .IN1(n6670), .IN2(n7342), .QN(n2866) );
  NAND2X0 U3853 ( .IN1(n6652), .IN2(n7343), .QN(n2865) );
  NAND2X0 U3854 ( .IN1(n2867), .IN2(n2868), .QN(n2863) );
  NAND2X0 U3855 ( .IN1(n9190), .IN2(n2569), .QN(n2868) );
  NAND2X0 U3856 ( .IN1(n7346), .IN2(P2_N371), .QN(n2867) );
  NAND2X0 U3857 ( .IN1(n2869), .IN2(n2870), .QN(P2_N4506) );
  NAND2X0 U3858 ( .IN1(P2_N4438), .IN2(n2702), .QN(n2870) );
  NAND2X0 U3859 ( .IN1(P2_N5493), .IN2(n7162), .QN(n2869) );
  OR2X1 U3860 ( .IN2(n2872), .IN1(n2871), .Q(P2_N5077) );
  NAND2X0 U3861 ( .IN1(n2873), .IN2(n2874), .QN(n2872) );
  NAND2X0 U3862 ( .IN1(n6669), .IN2(n7342), .QN(n2874) );
  NAND2X0 U3863 ( .IN1(n6651), .IN2(n7343), .QN(n2873) );
  NAND2X0 U3864 ( .IN1(n2875), .IN2(n2876), .QN(n2871) );
  NAND2X0 U3865 ( .IN1(n9194), .IN2(n2569), .QN(n2876) );
  NAND2X0 U3866 ( .IN1(n7346), .IN2(P2_N370), .QN(n2875) );
  NAND2X0 U3867 ( .IN1(n2877), .IN2(n2878), .QN(P2_N4505) );
  NAND2X0 U3868 ( .IN1(P2_N4437), .IN2(n2702), .QN(n2878) );
  NAND2X0 U3869 ( .IN1(P2_N5493), .IN2(P2_N5076), .QN(n2877) );
  OR2X1 U3870 ( .IN2(n2880), .IN1(n2879), .Q(P2_N5076) );
  NAND2X0 U3871 ( .IN1(n2881), .IN2(n2882), .QN(n2880) );
  NAND2X0 U3872 ( .IN1(n6668), .IN2(n7342), .QN(n2882) );
  NAND2X0 U3873 ( .IN1(n6650), .IN2(n7343), .QN(n2881) );
  NAND2X0 U3874 ( .IN1(n2883), .IN2(n2884), .QN(n2879) );
  NAND2X0 U3875 ( .IN1(n9198), .IN2(n2569), .QN(n2884) );
  NAND2X0 U3876 ( .IN1(n7346), .IN2(P2_N369), .QN(n2883) );
  NAND2X0 U3877 ( .IN1(n2885), .IN2(n2886), .QN(P2_N4504) );
  NAND2X0 U3878 ( .IN1(P2_N4436), .IN2(n2702), .QN(n2886) );
  NAND2X0 U3879 ( .IN1(P2_N5493), .IN2(P2_N5075), .QN(n2885) );
  OR2X1 U3880 ( .IN2(n2888), .IN1(n2887), .Q(P2_N5075) );
  NAND2X0 U3881 ( .IN1(n2889), .IN2(n2890), .QN(n2888) );
  NAND2X0 U3882 ( .IN1(n6667), .IN2(n7342), .QN(n2890) );
  NAND2X0 U3883 ( .IN1(n6649), .IN2(n7343), .QN(n2889) );
  NAND2X0 U3884 ( .IN1(n2891), .IN2(n2892), .QN(n2887) );
  NAND2X0 U3885 ( .IN1(n9202), .IN2(n2569), .QN(n2892) );
  NAND2X0 U3886 ( .IN1(n7346), .IN2(P2_N368), .QN(n2891) );
  NAND2X0 U3887 ( .IN1(n2893), .IN2(n2894), .QN(P2_N4503) );
  NAND2X0 U3888 ( .IN1(P2_N4435), .IN2(n2702), .QN(n2894) );
  NAND2X0 U3889 ( .IN1(P2_N5493), .IN2(n7177), .QN(n2893) );
  OR2X1 U3890 ( .IN2(n2896), .IN1(n2895), .Q(P2_N5074) );
  NAND2X0 U3891 ( .IN1(n2897), .IN2(n2898), .QN(n2896) );
  NAND2X0 U3892 ( .IN1(n6666), .IN2(n7342), .QN(n2898) );
  NAND2X0 U3893 ( .IN1(n6648), .IN2(n7343), .QN(n2897) );
  NAND2X0 U3894 ( .IN1(n2899), .IN2(n2900), .QN(n2895) );
  NAND2X0 U3895 ( .IN1(n9206), .IN2(n2569), .QN(n2900) );
  NAND2X0 U3896 ( .IN1(n7346), .IN2(n18813), .QN(n2899) );
  NAND2X0 U3897 ( .IN1(n2901), .IN2(n2902), .QN(P2_N4502) );
  NAND2X0 U3898 ( .IN1(P2_N4434), .IN2(n2702), .QN(n2902) );
  NAND2X0 U3899 ( .IN1(P2_N5493), .IN2(n7181), .QN(n2901) );
  OR2X1 U3900 ( .IN2(n2904), .IN1(n2903), .Q(P2_N5073) );
  NAND2X0 U3901 ( .IN1(n2905), .IN2(n2906), .QN(n2904) );
  NAND2X0 U3902 ( .IN1(n6665), .IN2(n7342), .QN(n2906) );
  NAND2X0 U3903 ( .IN1(n6721), .IN2(n7343), .QN(n2905) );
  NAND2X0 U3904 ( .IN1(n2907), .IN2(n2908), .QN(n2903) );
  NAND2X0 U3905 ( .IN1(n9210), .IN2(n2569), .QN(n2908) );
  NAND2X0 U3906 ( .IN1(n7346), .IN2(n6683), .QN(n2907) );
  NAND2X0 U3907 ( .IN1(n2909), .IN2(n2910), .QN(P2_N4501) );
  NAND2X0 U3908 ( .IN1(P2_N4433), .IN2(n2702), .QN(n2910) );
  NAND2X0 U3909 ( .IN1(P2_N5493), .IN2(P2_N5072), .QN(n2909) );
  OR2X1 U3910 ( .IN2(n2912), .IN1(n2911), .Q(P2_N5072) );
  NAND2X0 U3911 ( .IN1(n2913), .IN2(n2914), .QN(n2912) );
  NAND2X0 U3912 ( .IN1(n6664), .IN2(n7342), .QN(n2914) );
  NAND2X0 U3913 ( .IN1(n6720), .IN2(n7343), .QN(n2913) );
  NAND2X0 U3914 ( .IN1(n2915), .IN2(n2916), .QN(n2911) );
  NAND2X0 U3915 ( .IN1(n9214), .IN2(n2569), .QN(n2916) );
  NAND2X0 U3916 ( .IN1(n7346), .IN2(n6682), .QN(n2915) );
  NAND2X0 U3917 ( .IN1(n2917), .IN2(n2918), .QN(P2_N4500) );
  NAND2X0 U3918 ( .IN1(P2_N4432), .IN2(n2702), .QN(n2918) );
  NAND2X0 U3733 ( .IN1(n10116), .IN2(n7343), .QN(n2769) );
  NAND2X0 U3734 ( .IN1(n2771), .IN2(n2772), .QN(n2767) );
  NAND2X0 U3735 ( .IN1(n9142), .IN2(n2569), .QN(n2772) );
  NAND2X0 U3736 ( .IN1(n7346), .IN2(P2_N383), .QN(n2771) );
  NAND2X0 U3737 ( .IN1(n2773), .IN2(n2774), .QN(P2_N4518) );
  NAND2X0 U3738 ( .IN1(P2_N4450), .IN2(n2702), .QN(n2774) );
  NAND2X0 U3739 ( .IN1(P2_N5493), .IN2(n7187), .QN(n2773) );
  OR2X1 U3740 ( .IN2(n2776), .IN1(n2775), .Q(P2_N5089) );
  NAND2X0 U3741 ( .IN1(n2777), .IN2(n2778), .QN(n2776) );
  NAND2X0 U3742 ( .IN1(n6680), .IN2(n7342), .QN(n2778) );
  NAND2X0 U3743 ( .IN1(n6663), .IN2(n7343), .QN(n2777) );
  NAND2X0 U3744 ( .IN1(n2779), .IN2(n2780), .QN(n2775) );
  NAND2X0 U3745 ( .IN1(n9146), .IN2(n2569), .QN(n2780) );
  NAND2X0 U3746 ( .IN1(n7346), .IN2(P2_N382), .QN(n2779) );
  NAND2X0 U3747 ( .IN1(n2781), .IN2(n2782), .QN(P2_N4517) );
  NAND2X0 U3748 ( .IN1(P2_N4449), .IN2(n2702), .QN(n2782) );
  NAND2X0 U3749 ( .IN1(P2_N5493), .IN2(n7194), .QN(n2781) );
  OR2X1 U3750 ( .IN2(n2784), .IN1(n2783), .Q(P2_N5088) );
  NAND2X0 U3751 ( .IN1(n2785), .IN2(n2786), .QN(n2784) );
  NAND2X0 U3752 ( .IN1(n6679), .IN2(n7342), .QN(n2786) );
  NAND2X0 U3753 ( .IN1(n6662), .IN2(n7343), .QN(n2785) );
  NAND2X0 U3754 ( .IN1(n2787), .IN2(n2788), .QN(n2783) );
  NAND2X0 U3755 ( .IN1(n9150), .IN2(n2569), .QN(n2788) );
  NAND2X0 U3756 ( .IN1(n7346), .IN2(P2_N381), .QN(n2787) );
  NAND2X0 U3757 ( .IN1(n2789), .IN2(n2790), .QN(P2_N4516) );
  NAND2X0 U3758 ( .IN1(P2_N4448), .IN2(n2702), .QN(n2790) );
  NAND2X0 U3759 ( .IN1(P2_N5493), .IN2(n7198), .QN(n2789) );
  OR2X1 U3760 ( .IN2(n2792), .IN1(n2791), .Q(P2_N5087) );
  NAND2X0 U3761 ( .IN1(n2793), .IN2(n2794), .QN(n2792) );
  NAND2X0 U3762 ( .IN1(n6678), .IN2(n7342), .QN(n2794) );
  NAND2X0 U3763 ( .IN1(n6661), .IN2(n7343), .QN(n2793) );
  NAND2X0 U3764 ( .IN1(n2795), .IN2(n2796), .QN(n2791) );
  NAND2X0 U3765 ( .IN1(n9154), .IN2(n2569), .QN(n2796) );
  NAND2X0 U3766 ( .IN1(n7346), .IN2(P2_N380), .QN(n2795) );
  NAND2X0 U3767 ( .IN1(n2797), .IN2(n2798), .QN(P2_N4515) );
  NAND2X0 U3768 ( .IN1(P2_N4447), .IN2(n2702), .QN(n2798) );
  NAND2X0 U3769 ( .IN1(P2_N5493), .IN2(n7202), .QN(n2797) );
  OR2X1 U3770 ( .IN2(n2800), .IN1(n2799), .Q(P2_N5086) );
  NAND2X0 U3771 ( .IN1(n2801), .IN2(n2802), .QN(n2800) );
  NAND2X0 U3772 ( .IN1(n6677), .IN2(n7342), .QN(n2802) );
  NAND2X0 U3773 ( .IN1(n6660), .IN2(n7343), .QN(n2801) );
  NAND2X0 U3774 ( .IN1(n2803), .IN2(n2804), .QN(n2799) );
  NAND2X0 U3775 ( .IN1(n9158), .IN2(n2569), .QN(n2804) );
  NAND2X0 U3776 ( .IN1(n7346), .IN2(P2_N379), .QN(n2803) );
  NAND2X0 U3777 ( .IN1(n2805), .IN2(n2806), .QN(P2_N4514) );
  NAND2X0 U3778 ( .IN1(P2_N4446), .IN2(n2702), .QN(n2806) );
  NAND2X0 U3779 ( .IN1(P2_N5493), .IN2(n7206), .QN(n2805) );
  OR2X1 U3780 ( .IN2(n2808), .IN1(n2807), .Q(P2_N5085) );
  NAND2X0 U3781 ( .IN1(n2809), .IN2(n2810), .QN(n2808) );
  NAND2X0 U3782 ( .IN1(n6676), .IN2(n7342), .QN(n2810) );
  NAND2X0 U3783 ( .IN1(n6659), .IN2(n7343), .QN(n2809) );
  NAND2X0 U3784 ( .IN1(n2811), .IN2(n2812), .QN(n2807) );
  NAND2X0 U3785 ( .IN1(n9162), .IN2(n2569), .QN(n2812) );
  NAND2X0 U3786 ( .IN1(n7346), .IN2(P2_N378), .QN(n2811) );
  NAND2X0 U3787 ( .IN1(n2813), .IN2(n2814), .QN(P2_N4513) );
  NAND2X0 U3788 ( .IN1(P2_N4445), .IN2(n2702), .QN(n2814) );
  NAND2X0 U3789 ( .IN1(P2_N5493), .IN2(n7209), .QN(n2813) );
  OR2X1 U3790 ( .IN2(n2816), .IN1(n2815), .Q(P2_N5084) );
  NAND2X0 U3791 ( .IN1(n2817), .IN2(n2818), .QN(n2816) );
  NAND2X0 U3792 ( .IN1(n6675), .IN2(n7342), .QN(n2818) );
  NAND2X0 U3793 ( .IN1(n6658), .IN2(n7343), .QN(n2817) );
  NAND2X0 U3794 ( .IN1(n2819), .IN2(n2820), .QN(n2815) );
  NAND2X0 U3795 ( .IN1(n9166), .IN2(n2569), .QN(n2820) );
  NAND2X0 U3796 ( .IN1(n7346), .IN2(P2_N377), .QN(n2819) );
  NAND2X0 U3797 ( .IN1(n2821), .IN2(n2822), .QN(P2_N4512) );
  NAND2X0 U3798 ( .IN1(P2_N4444), .IN2(n2702), .QN(n2822) );
  NAND2X0 U3799 ( .IN1(P2_N5493), .IN2(P2_N5083), .QN(n2821) );
  OR2X1 U3800 ( .IN2(n2824), .IN1(n2823), .Q(P2_N5083) );
  NAND2X0 U3801 ( .IN1(n2825), .IN2(n2826), .QN(n2824) );
  NAND2X0 U3802 ( .IN1(n6674), .IN2(n7342), .QN(n2826) );
  NAND2X0 U3803 ( .IN1(n6657), .IN2(n7343), .QN(n2825) );
  NAND2X0 U3804 ( .IN1(n2827), .IN2(n2828), .QN(n2823) );
  NAND2X0 U3805 ( .IN1(n9170), .IN2(n2569), .QN(n2828) );
  NAND2X0 U3806 ( .IN1(n7346), .IN2(P2_N376), .QN(n2827) );
  NAND2X0 U3807 ( .IN1(n2829), .IN2(n2830), .QN(P2_N4511) );
  NAND2X0 U3808 ( .IN1(P2_N4443), .IN2(n2702), .QN(n2830) );
  NAND2X0 U3809 ( .IN1(P2_N5493), .IN2(n7216), .QN(n2829) );
  OR2X1 U3810 ( .IN2(n2832), .IN1(n2831), .Q(P2_N5082) );
  NAND2X0 U3811 ( .IN1(n2833), .IN2(n2834), .QN(n2832) );
  NAND2X0 U3812 ( .IN1(n6673), .IN2(n7342), .QN(n2834) );
  NAND2X0 U3813 ( .IN1(n6656), .IN2(n7343), .QN(n2833) );
  NAND2X0 U3814 ( .IN1(n2835), .IN2(n2836), .QN(n2831) );
  NAND2X0 U3815 ( .IN1(n9174), .IN2(n2569), .QN(n2836) );
  NAND2X0 U3816 ( .IN1(n7346), .IN2(P2_N375), .QN(n2835) );
  NAND2X0 U3817 ( .IN1(n2837), .IN2(n2838), .QN(P2_N4510) );
  NAND2X0 U3818 ( .IN1(P2_N4442), .IN2(n2702), .QN(n2838) );
  NAND2X0 U3819 ( .IN1(P2_N5493), .IN2(n7220), .QN(n2837) );
  OR2X1 U3820 ( .IN2(n2840), .IN1(n2839), .Q(P2_N5081) );
  NAND2X0 U3821 ( .IN1(n2841), .IN2(n2842), .QN(n2840) );
  NAND2X0 U3822 ( .IN1(n6672), .IN2(n7342), .QN(n2842) );
  NAND2X0 U3823 ( .IN1(n6655), .IN2(n7343), .QN(n2841) );
  NAND2X0 U3824 ( .IN1(n2843), .IN2(n2844), .QN(n2839) );
  NAND2X0 U3825 ( .IN1(n9178), .IN2(n2569), .QN(n2844) );
  OR2X1 U3640 ( .IN2(n2695), .IN1(n2694), .Q(P2_N5099) );
  NAND2X0 U3641 ( .IN1(n2696), .IN2(n2697), .QN(n2695) );
  NAND2X0 U3642 ( .IN1(n9230), .IN2(n7342), .QN(n2697) );
  NAND2X0 U3643 ( .IN1(n9270), .IN2(n7343), .QN(n2696) );
  NAND2X0 U3644 ( .IN1(n2698), .IN2(n2699), .QN(n2694) );
  NAND2X0 U3645 ( .IN1(n9106), .IN2(n2569), .QN(n2699) );
  NAND2X0 U3646 ( .IN1(n7346), .IN2(P2_N392), .QN(n2698) );
  NAND2X0 U3647 ( .IN1(n2700), .IN2(n2701), .QN(P2_N4527) );
  NAND2X0 U3648 ( .IN1(P2_N4459), .IN2(n2702), .QN(n2701) );
  NAND2X0 U3649 ( .IN1(P2_N5493), .IN2(n7227), .QN(n2700) );
  OR2X1 U3650 ( .IN2(n2704), .IN1(n2703), .Q(P2_N5098) );
  NAND2X0 U3651 ( .IN1(n2705), .IN2(n2706), .QN(n2704) );
  NAND2X0 U3652 ( .IN1(n9234), .IN2(n7342), .QN(n2706) );
  NAND2X0 U3653 ( .IN1(n9274), .IN2(n7343), .QN(n2705) );
  NAND2X0 U3654 ( .IN1(n2707), .IN2(n2708), .QN(n2703) );
  NAND2X0 U3655 ( .IN1(n9110), .IN2(n2569), .QN(n2708) );
  NAND2X0 U3656 ( .IN1(n7346), .IN2(P2_N391), .QN(n2707) );
  NAND2X0 U3657 ( .IN1(n2709), .IN2(n2710), .QN(P2_N4526) );
  NAND2X0 U3658 ( .IN1(P2_N4458), .IN2(n2702), .QN(n2710) );
  NAND2X0 U3659 ( .IN1(P2_N5493), .IN2(P2_N5097), .QN(n2709) );
  OR2X1 U3660 ( .IN2(n2712), .IN1(n2711), .Q(P2_N5097) );
  NAND2X0 U3661 ( .IN1(n2713), .IN2(n2714), .QN(n2712) );
  NAND2X0 U3662 ( .IN1(n9238), .IN2(n7342), .QN(n2714) );
  NAND2X0 U3663 ( .IN1(n9278), .IN2(n7343), .QN(n2713) );
  NAND2X0 U3664 ( .IN1(n2715), .IN2(n2716), .QN(n2711) );
  NAND2X0 U3665 ( .IN1(n9114), .IN2(n2569), .QN(n2716) );
  NAND2X0 U3666 ( .IN1(n7346), .IN2(P2_N390), .QN(n2715) );
  NAND2X0 U3667 ( .IN1(n2717), .IN2(n2718), .QN(P2_N4525) );
  NAND2X0 U3668 ( .IN1(P2_N4457), .IN2(n2702), .QN(n2718) );
  NAND2X0 U3669 ( .IN1(P2_N5493), .IN2(P2_N5096), .QN(n2717) );
  OR2X1 U3670 ( .IN2(n2720), .IN1(n2719), .Q(P2_N5096) );
  NAND2X0 U3671 ( .IN1(n2721), .IN2(n2722), .QN(n2720) );
  NAND2X0 U3672 ( .IN1(n9242), .IN2(n7342), .QN(n2722) );
  NAND2X0 U3673 ( .IN1(n9282), .IN2(n7343), .QN(n2721) );
  NAND2X0 U3674 ( .IN1(n2723), .IN2(n2724), .QN(n2719) );
  NAND2X0 U3675 ( .IN1(n9118), .IN2(n2569), .QN(n2724) );
  NAND2X0 U3676 ( .IN1(n7346), .IN2(P2_N389), .QN(n2723) );
  NAND2X0 U3677 ( .IN1(n2725), .IN2(n2726), .QN(P2_N4524) );
  NAND2X0 U3678 ( .IN1(P2_N4456), .IN2(n2702), .QN(n2726) );
  NAND2X0 U3679 ( .IN1(P2_N5493), .IN2(P2_N5095), .QN(n2725) );
  OR2X1 U3680 ( .IN2(n2728), .IN1(n2727), .Q(P2_N5095) );
  NAND2X0 U3681 ( .IN1(n2729), .IN2(n2730), .QN(n2728) );
  NAND2X0 U3682 ( .IN1(n9246), .IN2(n7342), .QN(n2730) );
  NAND2X0 U3683 ( .IN1(n9286), .IN2(n7343), .QN(n2729) );
  NAND2X0 U3684 ( .IN1(n2731), .IN2(n2732), .QN(n2727) );
  NAND2X0 U3685 ( .IN1(n9122), .IN2(n2569), .QN(n2732) );
  NAND2X0 U3686 ( .IN1(n7346), .IN2(P2_N388), .QN(n2731) );
  NAND2X0 U3687 ( .IN1(n2733), .IN2(n2734), .QN(P2_N4523) );
  NAND2X0 U3688 ( .IN1(P2_N4455), .IN2(n2702), .QN(n2734) );
  NAND2X0 U3689 ( .IN1(P2_N5493), .IN2(P2_N5094), .QN(n2733) );
  OR2X1 U3690 ( .IN2(n2736), .IN1(n2735), .Q(P2_N5094) );
  NAND2X0 U3691 ( .IN1(n2737), .IN2(n2738), .QN(n2736) );
  NAND2X0 U3692 ( .IN1(n9250), .IN2(n7342), .QN(n2738) );
  NAND2X0 U3693 ( .IN1(n9290), .IN2(n7343), .QN(n2737) );
  NAND2X0 U3694 ( .IN1(n2739), .IN2(n2740), .QN(n2735) );
  NAND2X0 U3695 ( .IN1(n9126), .IN2(n2569), .QN(n2740) );
  NAND2X0 U3696 ( .IN1(n7346), .IN2(P2_N387), .QN(n2739) );
  NAND2X0 U3697 ( .IN1(n2741), .IN2(n2742), .QN(P2_N4522) );
  NAND2X0 U3698 ( .IN1(P2_N4454), .IN2(n2702), .QN(n2742) );
  NAND2X0 U3699 ( .IN1(P2_N5493), .IN2(P2_N5093), .QN(n2741) );
  OR2X1 U3700 ( .IN2(n2744), .IN1(n2743), .Q(P2_N5093) );
  NAND2X0 U3701 ( .IN1(n2745), .IN2(n2746), .QN(n2744) );
  NAND2X0 U3702 ( .IN1(n9254), .IN2(n7342), .QN(n2746) );
  NAND2X0 U3703 ( .IN1(n9294), .IN2(n7343), .QN(n2745) );
  NAND2X0 U3704 ( .IN1(n2747), .IN2(n2748), .QN(n2743) );
  NAND2X0 U3705 ( .IN1(n9130), .IN2(n2569), .QN(n2748) );
  NAND2X0 U3706 ( .IN1(n7346), .IN2(P2_N386), .QN(n2747) );
  NAND2X0 U3707 ( .IN1(n2749), .IN2(n2750), .QN(P2_N4521) );
  NAND2X0 U3708 ( .IN1(P2_N4453), .IN2(n2702), .QN(n2750) );
  NAND2X0 U3709 ( .IN1(P2_N5493), .IN2(n7252), .QN(n2749) );
  OR2X1 U3710 ( .IN2(n2752), .IN1(n2751), .Q(P2_N5092) );
  NAND2X0 U3711 ( .IN1(n2753), .IN2(n2754), .QN(n2752) );
  NAND2X0 U3712 ( .IN1(n9258), .IN2(n7342), .QN(n2754) );
  NAND2X0 U3713 ( .IN1(n9298), .IN2(n7343), .QN(n2753) );
  NAND2X0 U3714 ( .IN1(n2755), .IN2(n2756), .QN(n2751) );
  NAND2X0 U3715 ( .IN1(n9134), .IN2(n2569), .QN(n2756) );
  NAND2X0 U3716 ( .IN1(n7346), .IN2(P2_N385), .QN(n2755) );
  NAND2X0 U3717 ( .IN1(n2757), .IN2(n2758), .QN(P2_N4520) );
  NAND2X0 U3718 ( .IN1(P2_N4452), .IN2(n2702), .QN(n2758) );
  NAND2X0 U3719 ( .IN1(P2_N5493), .IN2(n7259), .QN(n2757) );
  OR2X1 U3720 ( .IN2(n2760), .IN1(n2759), .Q(P2_N5091) );
  NAND2X0 U3721 ( .IN1(n2761), .IN2(n2762), .QN(n2760) );
  NAND2X0 U3722 ( .IN1(n9262), .IN2(n7342), .QN(n2762) );
  NAND2X0 U3723 ( .IN1(n9302), .IN2(n7343), .QN(n2761) );
  NAND2X0 U3724 ( .IN1(n2763), .IN2(n2764), .QN(n2759) );
  NAND2X0 U3725 ( .IN1(n9138), .IN2(n2569), .QN(n2764) );
  NAND2X0 U3726 ( .IN1(n7346), .IN2(P2_N384), .QN(n2763) );
  NAND2X0 U3727 ( .IN1(n2765), .IN2(n2766), .QN(P2_N4519) );
  NAND2X0 U3728 ( .IN1(P2_N4451), .IN2(n2702), .QN(n2766) );
  NAND2X0 U3729 ( .IN1(P2_N5493), .IN2(n7263), .QN(n2765) );
  OR2X1 U3730 ( .IN2(n2768), .IN1(n2767), .Q(P2_N5090) );
  NAND2X0 U3731 ( .IN1(n2769), .IN2(n2770), .QN(n2768) );
  NAND2X0 U3732 ( .IN1(n10111), .IN2(n7342), .QN(n2770) );
  NAND2X0 U3541 ( .IN1(n2599), .IN2(P2_N4515), .QN(n2624) );
  NAND2X0 U3542 ( .IN1(P2_N380), .IN2(P2_N5497), .QN(n2623) );
  NAND2X0 U3543 ( .IN1(n2625), .IN2(n2626), .QN(P2_N4677) );
  NAND2X0 U3544 ( .IN1(n2599), .IN2(P2_N4514), .QN(n2626) );
  NAND2X0 U3545 ( .IN1(P2_N379), .IN2(P2_N5497), .QN(n2625) );
  NAND2X0 U3546 ( .IN1(n2627), .IN2(n2628), .QN(P2_N4676) );
  NAND2X0 U3547 ( .IN1(n2599), .IN2(P2_N4513), .QN(n2628) );
  NAND2X0 U3548 ( .IN1(P2_N378), .IN2(P2_N5497), .QN(n2627) );
  NAND2X0 U3549 ( .IN1(n2629), .IN2(n2630), .QN(P2_N4675) );
  NAND2X0 U3550 ( .IN1(n2599), .IN2(P2_N4512), .QN(n2630) );
  NAND2X0 U3551 ( .IN1(P2_N377), .IN2(P2_N5497), .QN(n2629) );
  NAND2X0 U3552 ( .IN1(n2631), .IN2(n2632), .QN(P2_N4674) );
  NAND2X0 U3553 ( .IN1(n2599), .IN2(P2_N4511), .QN(n2632) );
  NAND2X0 U3554 ( .IN1(P2_N376), .IN2(P2_N5497), .QN(n2631) );
  NAND2X0 U3555 ( .IN1(n2633), .IN2(n2634), .QN(P2_N4673) );
  NAND2X0 U3556 ( .IN1(n2599), .IN2(P2_N4510), .QN(n2634) );
  NAND2X0 U3557 ( .IN1(P2_N375), .IN2(P2_N5497), .QN(n2633) );
  NAND2X0 U3558 ( .IN1(n2635), .IN2(n2636), .QN(P2_N4672) );
  NAND2X0 U3559 ( .IN1(n2599), .IN2(P2_N4509), .QN(n2636) );
  NAND2X0 U3560 ( .IN1(P2_N374), .IN2(P2_N5497), .QN(n2635) );
  NAND2X0 U3561 ( .IN1(n2637), .IN2(n2638), .QN(P2_N4671) );
  NAND2X0 U3562 ( .IN1(n2599), .IN2(P2_N4508), .QN(n2638) );
  NAND2X0 U3563 ( .IN1(P2_N373), .IN2(P2_N5497), .QN(n2637) );
  NAND2X0 U3564 ( .IN1(n2639), .IN2(n2640), .QN(P2_N4670) );
  NAND2X0 U3565 ( .IN1(n2599), .IN2(P2_N4507), .QN(n2640) );
  NAND2X0 U3566 ( .IN1(P2_N372), .IN2(P2_N5497), .QN(n2639) );
  NAND2X0 U3567 ( .IN1(n2641), .IN2(n2642), .QN(P2_N4669) );
  NAND2X0 U3568 ( .IN1(n2599), .IN2(P2_N4506), .QN(n2642) );
  NAND2X0 U3569 ( .IN1(P2_N371), .IN2(P2_N5497), .QN(n2641) );
  NAND2X0 U3570 ( .IN1(n2643), .IN2(n2644), .QN(P2_N4668) );
  NAND2X0 U3571 ( .IN1(n2599), .IN2(P2_N4505), .QN(n2644) );
  NAND2X0 U3572 ( .IN1(P2_N370), .IN2(P2_N5497), .QN(n2643) );
  NAND2X0 U3573 ( .IN1(n2645), .IN2(n2646), .QN(P2_N4667) );
  NAND2X0 U3574 ( .IN1(n2599), .IN2(P2_N4504), .QN(n2646) );
  NAND2X0 U3575 ( .IN1(P2_N369), .IN2(P2_N5497), .QN(n2645) );
  NAND2X0 U3576 ( .IN1(n2647), .IN2(n2648), .QN(P2_N4666) );
  NAND2X0 U3577 ( .IN1(n2599), .IN2(P2_N4503), .QN(n2648) );
  NAND2X0 U3578 ( .IN1(P2_N368), .IN2(P2_N5497), .QN(n2647) );
  NAND2X0 U3579 ( .IN1(n2649), .IN2(n2650), .QN(P2_N4665) );
  NAND2X0 U3580 ( .IN1(n2599), .IN2(P2_N4502), .QN(n2650) );
  NAND2X0 U3581 ( .IN1(n18813), .IN2(P2_N5497), .QN(n2649) );
  NAND2X0 U3582 ( .IN1(n2651), .IN2(n2652), .QN(P2_N4664) );
  NAND2X0 U3583 ( .IN1(n2599), .IN2(P2_N4501), .QN(n2652) );
  NAND2X0 U3584 ( .IN1(n6683), .IN2(P2_N5497), .QN(n2651) );
  NAND2X0 U3585 ( .IN1(n2653), .IN2(n2654), .QN(P2_N4663) );
  NAND2X0 U3586 ( .IN1(n2599), .IN2(P2_N4500), .QN(n2654) );
  NAND2X0 U3587 ( .IN1(n6682), .IN2(P2_N5497), .QN(n2653) );
  NAND2X0 U3588 ( .IN1(n2655), .IN2(n2656), .QN(P2_N4662) );
  NAND2X0 U3589 ( .IN1(P2_N4499), .IN2(n2599), .QN(n2656) );
  AND2X1 U3590 ( .IN1(n2657), .IN2(n7398), .Q(n2599) );
  NAND2X0 U3592 ( .IN1(n6681), .IN2(P2_N5497), .QN(n2655) );
  NOR2X0 U3599 ( .QN(P2_N4661), .IN1(n2657), .IN2(n7398) );
  OR2X1 U3602 ( .IN2(n7398), .IN1(P2_N4561), .Q(P2_N4626) );
  AND2X1 U3605 ( .IN1(P2_N395), .IN2(n2662), .Q(P2_N455) );
  NAND2X0 U3606 ( .IN1(n2663), .IN2(n2664), .QN(n2662) );
  NOR2X0 U3607 ( .QN(n2664), .IN1(n2665), .IN2(n2666) );
  NAND2X0 U3608 ( .IN1(n2667), .IN2(n2668), .QN(n2666) );
  AND2X1 U3609 ( .IN1(n2669), .IN2(n2670), .Q(n2668) );
  NOR2X0 U3610 ( .QN(n2670), .IN1(P2_N418), .IN2(P2_N417) );
  NOR2X0 U3611 ( .QN(n2669), .IN1(P2_N416), .IN2(P2_N415) );
  NOR2X0 U3612 ( .QN(n2667), .IN1(P2_N412), .IN2(n2671) );
  OR2X1 U3613 ( .IN2(P2_N413), .IN1(P2_N414), .Q(n2671) );
  OR2X1 U3614 ( .IN2(n2673), .IN1(n2672), .Q(n2665) );
  NAND2X0 U3615 ( .IN1(n2674), .IN2(n2675), .QN(n2673) );
  NOR2X0 U3616 ( .QN(n2675), .IN1(P2_N422), .IN2(P2_N421) );
  NOR2X0 U3617 ( .QN(n2674), .IN1(P2_N420), .IN2(P2_N419) );
  NAND2X0 U3618 ( .IN1(n2676), .IN2(n2677), .QN(n2672) );
  NOR2X0 U3619 ( .QN(n2677), .IN1(P2_N426), .IN2(P2_N425) );
  NOR2X0 U3620 ( .QN(n2676), .IN1(P2_N424), .IN2(P2_N423) );
  NOR2X0 U3621 ( .QN(n2663), .IN1(n2678), .IN2(n2679) );
  NAND2X0 U3622 ( .IN1(n2680), .IN2(n2681), .QN(n2679) );
  AND2X1 U3623 ( .IN1(n2682), .IN2(n2683), .Q(n2681) );
  NOR2X0 U3624 ( .QN(n2683), .IN1(P2_N404), .IN2(P2_N403) );
  NOR2X0 U3625 ( .QN(n2682), .IN1(P2_N402), .IN2(P2_N401) );
  NOR2X0 U3626 ( .QN(n2680), .IN1(P2_N398), .IN2(n2684) );
  OR2X1 U3627 ( .IN2(P2_N399), .IN1(P2_N400), .Q(n2684) );
  NAND2X0 U3628 ( .IN1(n2685), .IN2(n2686), .QN(n2678) );
  AND2X1 U3629 ( .IN1(n2687), .IN2(n2688), .Q(n2686) );
  NOR2X0 U3630 ( .QN(n2688), .IN1(P2_N411), .IN2(P2_N410) );
  NOR2X0 U3631 ( .QN(n2687), .IN1(P2_N409), .IN2(P2_N408) );
  NOR2X0 U3632 ( .QN(n2685), .IN1(P2_N405), .IN2(n2689) );
  OR2X1 U3633 ( .IN2(P2_N406), .IN1(P2_N407), .Q(n2689) );
  NAND2X0 U3634 ( .IN1(n2690), .IN2(n2691), .QN(P2_N4528) );
  NAND2X0 U3635 ( .IN1(P2_N4460), .IN2(n2589), .QN(n2691) );
  NAND2X0 U3636 ( .IN1(n6993), .IN2(n2692), .QN(n2589) );
  NAND2X0 U3637 ( .IN1(P2_N506), .IN2(n7341), .QN(n2692) );
  NAND2X0 U3639 ( .IN1(P2_N5493), .IN2(P2_N5099), .QN(n2690) );
  NAND2X0 U3447 ( .IN1(n2042), .IN2(n2554), .QN(P2_N5013) );
  NAND2X0 U3448 ( .IN1(n7016), .IN2(n2044), .QN(n2554) );
  NAND2X0 U3449 ( .IN1(n2045), .IN2(n2555), .QN(P2_N5012) );
  NAND2X0 U3450 ( .IN1(n7016), .IN2(n2047), .QN(n2555) );
  NAND2X0 U3451 ( .IN1(n2048), .IN2(n2556), .QN(P2_N5011) );
  NAND2X0 U3452 ( .IN1(n7016), .IN2(n2050), .QN(n2556) );
  NAND2X0 U3453 ( .IN1(n2051), .IN2(n2557), .QN(P2_N5010) );
  NAND2X0 U3454 ( .IN1(n7006), .IN2(n2053), .QN(n2557) );
  NAND2X0 U3455 ( .IN1(n2054), .IN2(n2558), .QN(P2_N5009) );
  NAND2X0 U3456 ( .IN1(n7006), .IN2(n2056), .QN(n2558) );
  NAND2X0 U3457 ( .IN1(n2057), .IN2(n2559), .QN(P2_N5008) );
  NAND2X0 U3458 ( .IN1(n7006), .IN2(n2059), .QN(n2559) );
  NAND2X0 U3459 ( .IN1(n2060), .IN2(n2560), .QN(P2_N5007) );
  NAND2X0 U3460 ( .IN1(n7006), .IN2(n2062), .QN(n2560) );
  NAND2X0 U3461 ( .IN1(n2063), .IN2(n2561), .QN(P2_N5006) );
  NAND2X0 U3462 ( .IN1(n7006), .IN2(n2065), .QN(n2561) );
  OR2X1 U3464 ( .IN2(n2564), .IN1(n2563), .Q(P2_N497) );
  NAND2X0 U3465 ( .IN1(n2565), .IN2(n2566), .QN(n2564) );
  NAND2X0 U3466 ( .IN1(n8878), .IN2(n7342), .QN(n2566) );
  NAND2X0 U3467 ( .IN1(n8870), .IN2(n7343), .QN(n2565) );
  NAND2X0 U3468 ( .IN1(n2567), .IN2(n2568), .QN(n2563) );
  NAND2X0 U3469 ( .IN1(n8874), .IN2(n2569), .QN(n2568) );
  OR2X1 U3470 ( .IN2(n2571), .IN1(n2570), .Q(P2_N5100) );
  NAND2X0 U3471 ( .IN1(n2572), .IN2(n2573), .QN(n2571) );
  NAND2X0 U3472 ( .IN1(n9226), .IN2(n7342), .QN(n2573) );
  NAND2X0 U3473 ( .IN1(n9266), .IN2(n7343), .QN(n2572) );
  NAND2X0 U3474 ( .IN1(n2574), .IN2(n2575), .QN(n2570) );
  NAND2X0 U3475 ( .IN1(n9102), .IN2(n2569), .QN(n2575) );
  NAND2X0 U3476 ( .IN1(P2_N393), .IN2(n7346), .QN(n2574) );
  NAND2X0 U3477 ( .IN1(n2576), .IN2(n7446), .QN(P2_N4809) );
  NAND2X0 U3479 ( .IN1(n2576), .IN2(n7447), .QN(P2_N4808) );
  NAND2X0 U3481 ( .IN1(n7423), .IN2(P2_N394), .QN(n2576) );
  NAND2X0 U3483 ( .IN1(n2581), .IN2(P2_N4462), .QN(n2580) );
  NAND2X0 U3484 ( .IN1(n2582), .IN2(n2172), .QN(n2579) );
  NAND2X0 U3485 ( .IN1(n2583), .IN2(n2584), .QN(n2172) );
  NAND2X0 U3486 ( .IN1(N70), .IN2(n6739), .QN(n2584) );
  NAND2X0 U3487 ( .IN1(n9345), .IN2(N5), .QN(n2583) );
  NAND2X0 U3489 ( .IN1(n2581), .IN2(P2_N4461), .QN(n2587) );
  NOR2X0 U3490 ( .QN(n2581), .IN1(n2588), .IN2(n7421) );
  INVX0 U3492 ( .ZN(n2588), .INP(n2589) );
  NAND2X0 U3493 ( .IN1(n2582), .IN2(n2175), .QN(n2586) );
  NAND2X0 U3494 ( .IN1(n2590), .IN2(n2591), .QN(n2175) );
  NAND2X0 U3495 ( .IN1(N69), .IN2(n6739), .QN(n2591) );
  NAND2X0 U3496 ( .IN1(n10103), .IN2(N5), .QN(n2590) );
  NAND2X0 U3497 ( .IN1(n2592), .IN2(n2593), .QN(n2582) );
  NAND2X0 U3498 ( .IN1(n7420), .IN2(n7012), .QN(n2593) );
  AND2X1 U3499 ( .IN1(n2594), .IN2(n2595), .Q(n2592) );
  NAND2X0 U3500 ( .IN1(P2_N543), .IN2(n7012), .QN(n2595) );
  AND2X1 U3501 ( .IN1(P2_N542), .IN2(P2_N541), .Q(P2_N543) );
  NAND2X0 U3502 ( .IN1(n7418), .IN2(n7012), .QN(n2594) );
  NAND2X0 U3504 ( .IN1(n2597), .IN2(n2598), .QN(P2_N4690) );
  NAND2X0 U3505 ( .IN1(n2599), .IN2(P2_N4527), .QN(n2598) );
  NAND2X0 U3506 ( .IN1(P2_N392), .IN2(P2_N5497), .QN(n2597) );
  NAND2X0 U3507 ( .IN1(n2601), .IN2(n2602), .QN(P2_N4689) );
  NAND2X0 U3508 ( .IN1(n2599), .IN2(P2_N4526), .QN(n2602) );
  NAND2X0 U3509 ( .IN1(P2_N391), .IN2(P2_N5497), .QN(n2601) );
  NAND2X0 U3510 ( .IN1(n2603), .IN2(n2604), .QN(P2_N4688) );
  NAND2X0 U3511 ( .IN1(n2599), .IN2(P2_N4525), .QN(n2604) );
  NAND2X0 U3512 ( .IN1(P2_N390), .IN2(P2_N5497), .QN(n2603) );
  NAND2X0 U3513 ( .IN1(n2605), .IN2(n2606), .QN(P2_N4687) );
  NAND2X0 U3514 ( .IN1(n2599), .IN2(P2_N4524), .QN(n2606) );
  NAND2X0 U3515 ( .IN1(P2_N389), .IN2(P2_N5497), .QN(n2605) );
  NAND2X0 U3516 ( .IN1(n2607), .IN2(n2608), .QN(P2_N4686) );
  NAND2X0 U3517 ( .IN1(n2599), .IN2(P2_N4523), .QN(n2608) );
  NAND2X0 U3518 ( .IN1(P2_N388), .IN2(P2_N5497), .QN(n2607) );
  NAND2X0 U3519 ( .IN1(n2609), .IN2(n2610), .QN(P2_N4685) );
  NAND2X0 U3520 ( .IN1(n2599), .IN2(P2_N4522), .QN(n2610) );
  NAND2X0 U3521 ( .IN1(P2_N387), .IN2(P2_N5497), .QN(n2609) );
  NAND2X0 U3522 ( .IN1(n2611), .IN2(n2612), .QN(P2_N4684) );
  NAND2X0 U3523 ( .IN1(n2599), .IN2(P2_N4521), .QN(n2612) );
  NAND2X0 U3524 ( .IN1(P2_N386), .IN2(P2_N5497), .QN(n2611) );
  NAND2X0 U3525 ( .IN1(n2613), .IN2(n2614), .QN(P2_N4683) );
  NAND2X0 U3526 ( .IN1(n2599), .IN2(P2_N4520), .QN(n2614) );
  NAND2X0 U3527 ( .IN1(P2_N385), .IN2(P2_N5497), .QN(n2613) );
  NAND2X0 U3528 ( .IN1(n2615), .IN2(n2616), .QN(P2_N4682) );
  NAND2X0 U3529 ( .IN1(n2599), .IN2(P2_N4519), .QN(n2616) );
  NAND2X0 U3530 ( .IN1(P2_N384), .IN2(P2_N5497), .QN(n2615) );
  NAND2X0 U3531 ( .IN1(n2617), .IN2(n2618), .QN(P2_N4681) );
  NAND2X0 U3532 ( .IN1(n2599), .IN2(P2_N4518), .QN(n2618) );
  NAND2X0 U3533 ( .IN1(P2_N383), .IN2(P2_N5497), .QN(n2617) );
  NAND2X0 U3534 ( .IN1(n2619), .IN2(n2620), .QN(P2_N4680) );
  NAND2X0 U3535 ( .IN1(n2599), .IN2(P2_N4517), .QN(n2620) );
  NAND2X0 U3536 ( .IN1(P2_N382), .IN2(P2_N5497), .QN(n2619) );
  NAND2X0 U3537 ( .IN1(n2621), .IN2(n2622), .QN(P2_N4679) );
  NAND2X0 U3538 ( .IN1(n2599), .IN2(P2_N4516), .QN(n2622) );
  NAND2X0 U3539 ( .IN1(P2_N381), .IN2(P2_N5497), .QN(n2621) );
  NAND2X0 U3540 ( .IN1(n2623), .IN2(n2624), .QN(P2_N4678) );
  NAND2X0 U3353 ( .IN1(P2_N5089), .IN2(n7279), .QN(n2505) );
  NAND2X0 U3354 ( .IN1(P2_N5089), .IN2(P2_N5069), .QN(n2504) );
  NAND2X0 U3355 ( .IN1(n2506), .IN2(n2507), .QN(P2_N5338) );
  NAND2X0 U3356 ( .IN1(P2_N5088), .IN2(n7279), .QN(n2507) );
  NAND2X0 U3357 ( .IN1(P2_N5088), .IN2(P2_N5069), .QN(n2506) );
  NAND2X0 U3358 ( .IN1(n2508), .IN2(n2509), .QN(P2_N5337) );
  NAND2X0 U3359 ( .IN1(P2_N5087), .IN2(n7279), .QN(n2509) );
  NAND2X0 U3360 ( .IN1(n7198), .IN2(P2_N5069), .QN(n2508) );
  NAND2X0 U3361 ( .IN1(n2510), .IN2(n2511), .QN(P2_N5336) );
  NAND2X0 U3362 ( .IN1(P2_N5086), .IN2(n7279), .QN(n2511) );
  NAND2X0 U3363 ( .IN1(n7202), .IN2(P2_N5069), .QN(n2510) );
  NAND2X0 U3364 ( .IN1(n2512), .IN2(n2513), .QN(P2_N5335) );
  NAND2X0 U3365 ( .IN1(P2_N5085), .IN2(n7279), .QN(n2513) );
  NAND2X0 U3366 ( .IN1(P2_N5085), .IN2(P2_N5069), .QN(n2512) );
  NAND2X0 U3367 ( .IN1(n2514), .IN2(n2515), .QN(P2_N5334) );
  NAND2X0 U3368 ( .IN1(P2_N5084), .IN2(n7279), .QN(n2515) );
  NAND2X0 U3369 ( .IN1(P2_N5084), .IN2(P2_N5069), .QN(n2514) );
  NAND2X0 U3370 ( .IN1(n2516), .IN2(n2517), .QN(P2_N5333) );
  NAND2X0 U3371 ( .IN1(n7210), .IN2(n7279), .QN(n2517) );
  NAND2X0 U3372 ( .IN1(n7210), .IN2(P2_N5069), .QN(n2516) );
  NAND2X0 U3373 ( .IN1(n2518), .IN2(n2519), .QN(P2_N5332) );
  NAND2X0 U3374 ( .IN1(n7216), .IN2(n7279), .QN(n2519) );
  NAND2X0 U3375 ( .IN1(n7216), .IN2(P2_N5069), .QN(n2518) );
  NAND2X0 U3376 ( .IN1(n2520), .IN2(n2521), .QN(P2_N5331) );
  NAND2X0 U3377 ( .IN1(P2_N5081), .IN2(n7279), .QN(n2521) );
  NAND2X0 U3378 ( .IN1(P2_N5081), .IN2(P2_N5069), .QN(n2520) );
  NAND2X0 U3379 ( .IN1(n2522), .IN2(n2523), .QN(P2_N5330) );
  NAND2X0 U3380 ( .IN1(P2_N5080), .IN2(n7279), .QN(n2523) );
  NAND2X0 U3381 ( .IN1(P2_N5080), .IN2(P2_N5069), .QN(n2522) );
  NAND2X0 U3382 ( .IN1(n2524), .IN2(n2525), .QN(P2_N5329) );
  NAND2X0 U3383 ( .IN1(P2_N5079), .IN2(n7279), .QN(n2525) );
  NAND2X0 U3384 ( .IN1(P2_N5079), .IN2(P2_N5069), .QN(n2524) );
  NAND2X0 U3385 ( .IN1(n2526), .IN2(n2527), .QN(P2_N5328) );
  NAND2X0 U3386 ( .IN1(P2_N5078), .IN2(n7279), .QN(n2527) );
  NAND2X0 U3387 ( .IN1(n7158), .IN2(P2_N5069), .QN(n2526) );
  NAND2X0 U3388 ( .IN1(n2528), .IN2(n2529), .QN(P2_N5327) );
  NAND2X0 U3389 ( .IN1(n7162), .IN2(n7279), .QN(n2529) );
  NAND2X0 U3390 ( .IN1(n7162), .IN2(P2_N5069), .QN(n2528) );
  NAND2X0 U3391 ( .IN1(n2530), .IN2(n2531), .QN(P2_N5326) );
  NAND2X0 U3392 ( .IN1(P2_N5076), .IN2(n7279), .QN(n2531) );
  NAND2X0 U3393 ( .IN1(P2_N5076), .IN2(P2_N5069), .QN(n2530) );
  NAND2X0 U3394 ( .IN1(n2532), .IN2(n2533), .QN(P2_N5325) );
  NAND2X0 U3395 ( .IN1(P2_N5075), .IN2(n7279), .QN(n2533) );
  NAND2X0 U3396 ( .IN1(P2_N5075), .IN2(P2_N5069), .QN(n2532) );
  NAND2X0 U3397 ( .IN1(n2534), .IN2(n2535), .QN(P2_N5324) );
  NAND2X0 U3398 ( .IN1(P2_N5074), .IN2(n7279), .QN(n2535) );
  NAND2X0 U3399 ( .IN1(P2_N5074), .IN2(P2_N5069), .QN(n2534) );
  NAND2X0 U3400 ( .IN1(n2536), .IN2(n2537), .QN(P2_N5323) );
  NAND2X0 U3401 ( .IN1(P2_N5073), .IN2(n7279), .QN(n2537) );
  NAND2X0 U3402 ( .IN1(P2_N5073), .IN2(P2_N5069), .QN(n2536) );
  NAND2X0 U3403 ( .IN1(n2538), .IN2(n2539), .QN(P2_N5322) );
  NAND2X0 U3404 ( .IN1(P2_N5072), .IN2(n7279), .QN(n2539) );
  NAND2X0 U3405 ( .IN1(P2_N5072), .IN2(P2_N5069), .QN(n2538) );
  NAND2X0 U3406 ( .IN1(n2540), .IN2(n2541), .QN(P2_N5321) );
  NAND2X0 U3407 ( .IN1(n7035), .IN2(n7279), .QN(n2541) );
  NAND2X0 U3409 ( .IN1(n7035), .IN2(P2_N5069), .QN(n2540) );
  AND2X1 U3410 ( .IN1(n2172), .IN2(n7012), .Q(P2_N5037) );
  AND2X1 U3411 ( .IN1(n2175), .IN2(n7012), .Q(P2_N5036) );
  NOR2X0 U3412 ( .QN(P2_N5035), .IN1(n7329), .IN2(n7007) );
  NOR2X0 U3413 ( .QN(P2_N5034), .IN1(n7327), .IN2(n7007) );
  NOR2X0 U3414 ( .QN(P2_N5033), .IN1(n7325), .IN2(n7007) );
  NOR2X0 U3415 ( .QN(P2_N5032), .IN1(n7323), .IN2(n7007) );
  NOR2X0 U3416 ( .QN(P2_N5031), .IN1(n7321), .IN2(n7007) );
  NOR2X0 U3417 ( .QN(P2_N5030), .IN1(n7319), .IN2(n7007) );
  NOR2X0 U3418 ( .QN(P2_N5029), .IN1(n7317), .IN2(n7011) );
  NOR2X0 U3419 ( .QN(P2_N5028), .IN1(n7315), .IN2(n7015) );
  NOR2X0 U3420 ( .QN(P2_N5027), .IN1(n7313), .IN2(n7013) );
  NOR2X0 U3421 ( .QN(P2_N5026), .IN1(n7311), .IN2(n7011) );
  NAND2X0 U3423 ( .IN1(n2006), .IN2(n2542), .QN(P2_N5025) );
  NAND2X0 U3424 ( .IN1(n7012), .IN2(n2008), .QN(n2542) );
  NAND2X0 U3425 ( .IN1(n2009), .IN2(n2543), .QN(P2_N5024) );
  NAND2X0 U3426 ( .IN1(n7012), .IN2(n2011), .QN(n2543) );
  NAND2X0 U3427 ( .IN1(n2012), .IN2(n2544), .QN(P2_N5023) );
  NAND2X0 U3428 ( .IN1(n7012), .IN2(n2014), .QN(n2544) );
  NAND2X0 U3429 ( .IN1(n2015), .IN2(n2545), .QN(P2_N5022) );
  NAND2X0 U3430 ( .IN1(n7012), .IN2(n2017), .QN(n2545) );
  NAND2X0 U3431 ( .IN1(n2018), .IN2(n2546), .QN(P2_N5021) );
  NAND2X0 U3432 ( .IN1(n7009), .IN2(n2020), .QN(n2546) );
  NAND2X0 U3433 ( .IN1(n2021), .IN2(n2547), .QN(P2_N5020) );
  NAND2X0 U3434 ( .IN1(n7009), .IN2(n2023), .QN(n2547) );
  NAND2X0 U3435 ( .IN1(n2024), .IN2(n2548), .QN(P2_N5019) );
  NAND2X0 U3436 ( .IN1(n7009), .IN2(n2026), .QN(n2548) );
  NAND2X0 U3437 ( .IN1(n2027), .IN2(n2549), .QN(P2_N5018) );
  NAND2X0 U3438 ( .IN1(n7009), .IN2(n2029), .QN(n2549) );
  NAND2X0 U3439 ( .IN1(n2030), .IN2(n2550), .QN(P2_N5017) );
  NAND2X0 U3440 ( .IN1(n7010), .IN2(n2032), .QN(n2550) );
  NAND2X0 U3441 ( .IN1(n2033), .IN2(n2551), .QN(P2_N5016) );
  NAND2X0 U3442 ( .IN1(n7010), .IN2(n2035), .QN(n2551) );
  NAND2X0 U3443 ( .IN1(n2036), .IN2(n2552), .QN(P2_N5015) );
  NAND2X0 U3444 ( .IN1(n7016), .IN2(n2038), .QN(n2552) );
  NAND2X0 U3445 ( .IN1(n2039), .IN2(n2553), .QN(P2_N5014) );
  NAND2X0 U3446 ( .IN1(n7016), .IN2(n2041), .QN(n2553) );
  NAND2X0 U3258 ( .IN1(P2_N4844), .IN2(n2252), .QN(n2434) );
  NAND2X0 U3259 ( .IN1(n2253), .IN2(P2_N362), .QN(n2433) );
  AND2X1 U3260 ( .IN1(P2_N4864), .IN2(n2254), .Q(n2431) );
  NOR2X0 U3261 ( .QN(n2429), .IN1(n2435), .IN2(n2436) );
  NAND2X0 U3262 ( .IN1(n2437), .IN2(n2438), .QN(n2436) );
  NAND2X0 U3263 ( .IN1(n2168), .IN2(P2_N916), .QN(n2438) );
  NAND2X0 U3264 ( .IN1(P2_N4694), .IN2(n2161), .QN(n2437) );
  AND2X1 U3265 ( .IN1(n6682), .IN2(n2166), .Q(n2435) );
  NAND2X0 U3266 ( .IN1(n2439), .IN2(n2440), .QN(P2_N5420) );
  NOR2X0 U3267 ( .QN(n2440), .IN1(n2441), .IN2(n2442) );
  NAND2X0 U3268 ( .IN1(n2443), .IN2(n2444), .QN(n2442) );
  NAND2X0 U3269 ( .IN1(P2_N4843), .IN2(n2252), .QN(n2444) );
  NOR2X0 U3270 ( .QN(n2252), .IN1(n2445), .IN2(n6993) );
  NAND2X0 U3271 ( .IN1(n2253), .IN2(P2_N363), .QN(n2443) );
  AND2X1 U3272 ( .IN1(P2_N5492), .IN2(n2169), .Q(n2253) );
  AND2X1 U3273 ( .IN1(P2_N4863), .IN2(n2254), .Q(n2441) );
  AND2X1 U3274 ( .IN1(n2169), .IN2(n6999), .Q(n2254) );
  INVX0 U3275 ( .ZN(n2169), .INP(n2445) );
  NAND2X0 U3276 ( .IN1(n2447), .IN2(n6590), .QN(n2445) );
  NOR2X0 U3277 ( .QN(n2439), .IN1(n2448), .IN2(n2449) );
  NAND2X0 U3278 ( .IN1(n2450), .IN2(n2451), .QN(n2449) );
  NAND2X0 U3279 ( .IN1(n2168), .IN2(P2_N915), .QN(n2451) );
  NAND2X0 U3281 ( .IN1(P2_N4693), .IN2(n2161), .QN(n2450) );
  NOR2X0 U3282 ( .QN(n2161), .IN1(n6589), .IN2(n2452) );
  AND2X1 U3283 ( .IN1(n6681), .IN2(n6589), .Q(n2448) );
  NAND2X0 U3284 ( .IN1(n2453), .IN2(n2454), .QN(P2_N5419) );
  INVX0 U3285 ( .ZN(n2454), .INP(P2_N5440) );
  NAND2X0 U3286 ( .IN1(n2455), .IN2(n6590), .QN(P2_N5440) );
  NOR2X0 U3287 ( .QN(n2455), .IN1(n2456), .IN2(n2457) );
  NOR2X0 U3288 ( .QN(n2457), .IN1(P2_N499), .IN2(n7013) );
  AND2X1 U3289 ( .IN1(P2_N4692), .IN2(n2459), .Q(n2456) );
  NAND2X0 U3290 ( .IN1(n2447), .IN2(P2_N4841), .QN(n2453) );
  NOR2X0 U3291 ( .QN(n2447), .IN1(n7415), .IN2(n2460) );
  INVX0 U3295 ( .ZN(n2460), .INP(P2_N499) );
  NAND2X0 U3296 ( .IN1(n2463), .IN2(n2464), .QN(P2_N531) );
  NAND2X0 U3297 ( .IN1(n2463), .IN2(n2465), .QN(P2_N530) );
  NAND2X0 U3298 ( .IN1(P2_N517), .IN2(n2464), .QN(n2465) );
  INVX0 U3299 ( .ZN(n2464), .INP(P2_N514) );
  AND2X1 U3300 ( .IN1(n2466), .IN2(n2467), .Q(n2463) );
  NOR2X0 U3301 ( .QN(n2466), .IN1(P2_N511), .IN2(P2_N508) );
  NAND2X0 U3303 ( .IN1(n2470), .IN2(n2467), .QN(n2469) );
  INVX0 U3304 ( .ZN(n2467), .INP(P2_N504) );
  NAND2X0 U3305 ( .IN1(n2471), .IN2(n2472), .QN(n2470) );
  NAND2X0 U3306 ( .IN1(n2473), .IN2(n2474), .QN(n2472) );
  NAND2X0 U3307 ( .IN1(n2475), .IN2(n2476), .QN(n2473) );
  NOR2X0 U3308 ( .QN(n2476), .IN1(P2_N519), .IN2(P2_N517) );
  NOR2X0 U3309 ( .QN(n2475), .IN1(P2_N514), .IN2(P2_N511) );
  OR2X1 U3310 ( .IN2(P2_N506), .IN1(n2474), .Q(n2471) );
  INVX0 U3311 ( .ZN(n2474), .INP(P2_N508) );
  NAND2X0 U3312 ( .IN1(P2_N506), .IN2(P2_N504), .QN(n2468) );
  NAND2X0 U3313 ( .IN1(n2477), .IN2(n2478), .QN(P2_N5352) );
  NAND2X0 U3314 ( .IN1(n7147), .IN2(n7279), .QN(n2478) );
  NAND2X0 U3315 ( .IN1(P2_N5102), .IN2(P2_N5069), .QN(n2477) );
  NAND2X0 U3316 ( .IN1(n2480), .IN2(n2481), .QN(P2_N5351) );
  NAND2X0 U3317 ( .IN1(P2_N497), .IN2(n7279), .QN(n2481) );
  NAND2X0 U3318 ( .IN1(n7265), .IN2(P2_N5069), .QN(n2480) );
  NAND2X0 U3319 ( .IN1(n2482), .IN2(n2483), .QN(P2_N5350) );
  NAND2X0 U3320 ( .IN1(P2_N5100), .IN2(n7279), .QN(n2483) );
  NAND2X0 U3321 ( .IN1(P2_N5100), .IN2(P2_N5069), .QN(n2482) );
  NAND2X0 U3322 ( .IN1(n2484), .IN2(n2485), .QN(P2_N5349) );
  NAND2X0 U3323 ( .IN1(P2_N5099), .IN2(n7279), .QN(n2485) );
  NAND2X0 U3324 ( .IN1(P2_N5099), .IN2(P2_N5069), .QN(n2484) );
  NAND2X0 U3325 ( .IN1(n2486), .IN2(n2487), .QN(P2_N5348) );
  NAND2X0 U3326 ( .IN1(P2_N5098), .IN2(n7279), .QN(n2487) );
  NAND2X0 U3327 ( .IN1(P2_N5098), .IN2(P2_N5069), .QN(n2486) );
  NAND2X0 U3328 ( .IN1(n2488), .IN2(n2489), .QN(P2_N5347) );
  NAND2X0 U3329 ( .IN1(P2_N5097), .IN2(n7279), .QN(n2489) );
  NAND2X0 U3330 ( .IN1(P2_N5097), .IN2(P2_N5069), .QN(n2488) );
  NAND2X0 U3331 ( .IN1(n2490), .IN2(n2491), .QN(P2_N5346) );
  NAND2X0 U3332 ( .IN1(P2_N5096), .IN2(n7279), .QN(n2491) );
  NAND2X0 U3333 ( .IN1(P2_N5096), .IN2(P2_N5069), .QN(n2490) );
  NAND2X0 U3334 ( .IN1(n2492), .IN2(n2493), .QN(P2_N5345) );
  NAND2X0 U3335 ( .IN1(P2_N5095), .IN2(n7279), .QN(n2493) );
  NAND2X0 U3336 ( .IN1(P2_N5095), .IN2(P2_N5069), .QN(n2492) );
  NAND2X0 U3337 ( .IN1(n2494), .IN2(n2495), .QN(P2_N5344) );
  NAND2X0 U3338 ( .IN1(n7242), .IN2(n7279), .QN(n2495) );
  NAND2X0 U3339 ( .IN1(P2_N5094), .IN2(P2_N5069), .QN(n2494) );
  NAND2X0 U3340 ( .IN1(n2496), .IN2(n2497), .QN(P2_N5343) );
  NAND2X0 U3341 ( .IN1(P2_N5093), .IN2(n7279), .QN(n2497) );
  NAND2X0 U3342 ( .IN1(n7247), .IN2(P2_N5069), .QN(n2496) );
  NAND2X0 U3343 ( .IN1(n2498), .IN2(n2499), .QN(P2_N5342) );
  NAND2X0 U3344 ( .IN1(P2_N5092), .IN2(n7279), .QN(n2499) );
  NAND2X0 U3345 ( .IN1(P2_N5092), .IN2(P2_N5069), .QN(n2498) );
  NAND2X0 U3346 ( .IN1(n2500), .IN2(n2501), .QN(P2_N5341) );
  NAND2X0 U3347 ( .IN1(n7259), .IN2(n7279), .QN(n2501) );
  NAND2X0 U3348 ( .IN1(P2_N5091), .IN2(P2_N5069), .QN(n2500) );
  NAND2X0 U3349 ( .IN1(n2502), .IN2(n2503), .QN(P2_N5340) );
  NAND2X0 U3350 ( .IN1(P2_N5090), .IN2(n7279), .QN(n2503) );
  NAND2X0 U3351 ( .IN1(P2_N5090), .IN2(P2_N5069), .QN(n2502) );
  NAND2X0 U3352 ( .IN1(n2504), .IN2(n2505), .QN(P2_N5339) );
  NAND2X0 U3165 ( .IN1(P2_N4703), .IN2(n2161), .QN(n2347) );
  AND2X1 U3166 ( .IN1(n9537), .IN2(n2166), .Q(n2345) );
  NAND2X0 U3167 ( .IN1(n2349), .IN2(n2350), .QN(P2_N5429) );
  NOR2X0 U3168 ( .QN(n2350), .IN1(n2351), .IN2(n2352) );
  NAND2X0 U3169 ( .IN1(n2353), .IN2(n2354), .QN(n2352) );
  NAND2X0 U3170 ( .IN1(P2_N4852), .IN2(n2252), .QN(n2354) );
  NAND2X0 U3171 ( .IN1(n2253), .IN2(P2_N354), .QN(n2353) );
  AND2X1 U3172 ( .IN1(P2_N4872), .IN2(n2254), .Q(n2351) );
  NOR2X0 U3173 ( .QN(n2349), .IN1(n2355), .IN2(n2356) );
  NAND2X0 U3174 ( .IN1(n2357), .IN2(n2358), .QN(n2356) );
  NAND2X0 U3175 ( .IN1(n2168), .IN2(P2_N924), .QN(n2358) );
  NAND2X0 U3176 ( .IN1(P2_N4702), .IN2(n2161), .QN(n2357) );
  AND2X1 U3177 ( .IN1(n9541), .IN2(n2166), .Q(n2355) );
  NAND2X0 U3178 ( .IN1(n2359), .IN2(n2360), .QN(P2_N5428) );
  NOR2X0 U3179 ( .QN(n2360), .IN1(n2361), .IN2(n2362) );
  NAND2X0 U3180 ( .IN1(n2363), .IN2(n2364), .QN(n2362) );
  NAND2X0 U3181 ( .IN1(P2_N4851), .IN2(n2252), .QN(n2364) );
  NAND2X0 U3182 ( .IN1(n2253), .IN2(P2_N355), .QN(n2363) );
  AND2X1 U3183 ( .IN1(P2_N4871), .IN2(n2254), .Q(n2361) );
  NOR2X0 U3184 ( .QN(n2359), .IN1(n2365), .IN2(n2366) );
  NAND2X0 U3185 ( .IN1(n2367), .IN2(n2368), .QN(n2366) );
  NAND2X0 U3186 ( .IN1(n2168), .IN2(P2_N923), .QN(n2368) );
  NAND2X0 U3187 ( .IN1(P2_N4701), .IN2(n2161), .QN(n2367) );
  AND2X1 U3188 ( .IN1(n9545), .IN2(n2166), .Q(n2365) );
  NAND2X0 U3189 ( .IN1(n2369), .IN2(n2370), .QN(P2_N5427) );
  NOR2X0 U3190 ( .QN(n2370), .IN1(n2371), .IN2(n2372) );
  NAND2X0 U3191 ( .IN1(n2373), .IN2(n2374), .QN(n2372) );
  NAND2X0 U3192 ( .IN1(P2_N4850), .IN2(n2252), .QN(n2374) );
  NAND2X0 U3193 ( .IN1(n2253), .IN2(P2_N356), .QN(n2373) );
  AND2X1 U3194 ( .IN1(P2_N4870), .IN2(n2254), .Q(n2371) );
  NOR2X0 U3195 ( .QN(n2369), .IN1(n2375), .IN2(n2376) );
  NAND2X0 U3196 ( .IN1(n2377), .IN2(n2378), .QN(n2376) );
  NAND2X0 U3197 ( .IN1(n2168), .IN2(P2_N922), .QN(n2378) );
  NAND2X0 U3198 ( .IN1(P2_N4700), .IN2(n2161), .QN(n2377) );
  AND2X1 U3199 ( .IN1(n9549), .IN2(n2166), .Q(n2375) );
  NAND2X0 U3200 ( .IN1(n2379), .IN2(n2380), .QN(P2_N5426) );
  NOR2X0 U3201 ( .QN(n2380), .IN1(n2381), .IN2(n2382) );
  NAND2X0 U3202 ( .IN1(n2383), .IN2(n2384), .QN(n2382) );
  NAND2X0 U3203 ( .IN1(P2_N4849), .IN2(n2252), .QN(n2384) );
  NAND2X0 U3204 ( .IN1(n2253), .IN2(P2_N357), .QN(n2383) );
  AND2X1 U3205 ( .IN1(P2_N4869), .IN2(n2254), .Q(n2381) );
  NOR2X0 U3206 ( .QN(n2379), .IN1(n2385), .IN2(n2386) );
  NAND2X0 U3207 ( .IN1(n2387), .IN2(n2388), .QN(n2386) );
  NAND2X0 U3208 ( .IN1(n2168), .IN2(P2_N921), .QN(n2388) );
  NAND2X0 U3209 ( .IN1(P2_N4699), .IN2(n2161), .QN(n2387) );
  AND2X1 U3210 ( .IN1(n9553), .IN2(n2166), .Q(n2385) );
  NAND2X0 U3211 ( .IN1(n2389), .IN2(n2390), .QN(P2_N5425) );
  NOR2X0 U3212 ( .QN(n2390), .IN1(n2391), .IN2(n2392) );
  NAND2X0 U3213 ( .IN1(n2393), .IN2(n2394), .QN(n2392) );
  NAND2X0 U3214 ( .IN1(P2_N4848), .IN2(n2252), .QN(n2394) );
  NAND2X0 U3215 ( .IN1(n2253), .IN2(P2_N358), .QN(n2393) );
  AND2X1 U3216 ( .IN1(P2_N4868), .IN2(n2254), .Q(n2391) );
  NOR2X0 U3217 ( .QN(n2389), .IN1(n2395), .IN2(n2396) );
  NAND2X0 U3218 ( .IN1(n2397), .IN2(n2398), .QN(n2396) );
  NAND2X0 U3219 ( .IN1(n2168), .IN2(P2_N920), .QN(n2398) );
  NAND2X0 U3220 ( .IN1(P2_N4698), .IN2(n2161), .QN(n2397) );
  AND2X1 U3221 ( .IN1(n9557), .IN2(n2166), .Q(n2395) );
  NAND2X0 U3222 ( .IN1(n2399), .IN2(n2400), .QN(P2_N5424) );
  NOR2X0 U3223 ( .QN(n2400), .IN1(n2401), .IN2(n2402) );
  NAND2X0 U3224 ( .IN1(n2403), .IN2(n2404), .QN(n2402) );
  NAND2X0 U3225 ( .IN1(P2_N4847), .IN2(n2252), .QN(n2404) );
  NAND2X0 U3226 ( .IN1(n2253), .IN2(P2_N359), .QN(n2403) );
  AND2X1 U3227 ( .IN1(P2_N4867), .IN2(n2254), .Q(n2401) );
  NOR2X0 U3228 ( .QN(n2399), .IN1(n2405), .IN2(n2406) );
  NAND2X0 U3229 ( .IN1(n2407), .IN2(n2408), .QN(n2406) );
  NAND2X0 U3230 ( .IN1(n2168), .IN2(P2_N919), .QN(n2408) );
  NAND2X0 U3231 ( .IN1(P2_N4697), .IN2(n2161), .QN(n2407) );
  AND2X1 U3232 ( .IN1(n9397), .IN2(n2166), .Q(n2405) );
  NAND2X0 U3233 ( .IN1(n2409), .IN2(n2410), .QN(P2_N5423) );
  NOR2X0 U3234 ( .QN(n2410), .IN1(n2411), .IN2(n2412) );
  NAND2X0 U3235 ( .IN1(n2413), .IN2(n2414), .QN(n2412) );
  NAND2X0 U3236 ( .IN1(P2_N4846), .IN2(n2252), .QN(n2414) );
  NAND2X0 U3237 ( .IN1(n2253), .IN2(P2_N360), .QN(n2413) );
  AND2X1 U3238 ( .IN1(P2_N4866), .IN2(n2254), .Q(n2411) );
  NOR2X0 U3239 ( .QN(n2409), .IN1(n2415), .IN2(n2416) );
  NAND2X0 U3240 ( .IN1(n2417), .IN2(n2418), .QN(n2416) );
  NAND2X0 U3241 ( .IN1(n2168), .IN2(P2_N918), .QN(n2418) );
  NAND2X0 U3242 ( .IN1(P2_N4696), .IN2(n2161), .QN(n2417) );
  AND2X1 U3243 ( .IN1(n6684), .IN2(n2166), .Q(n2415) );
  NAND2X0 U3244 ( .IN1(n2419), .IN2(n2420), .QN(P2_N5422) );
  NOR2X0 U3245 ( .QN(n2420), .IN1(n2421), .IN2(n2422) );
  NAND2X0 U3246 ( .IN1(n2423), .IN2(n2424), .QN(n2422) );
  NAND2X0 U3247 ( .IN1(P2_N4845), .IN2(n2252), .QN(n2424) );
  NAND2X0 U3248 ( .IN1(n2253), .IN2(P2_N361), .QN(n2423) );
  AND2X1 U3249 ( .IN1(P2_N4865), .IN2(n2254), .Q(n2421) );
  NOR2X0 U3250 ( .QN(n2419), .IN1(n2425), .IN2(n2426) );
  NAND2X0 U3251 ( .IN1(n2427), .IN2(n2428), .QN(n2426) );
  NAND2X0 U3252 ( .IN1(n2168), .IN2(P2_N917), .QN(n2428) );
  NAND2X0 U3253 ( .IN1(P2_N4695), .IN2(n2161), .QN(n2427) );
  AND2X1 U3254 ( .IN1(n6683), .IN2(n2166), .Q(n2425) );
  NAND2X0 U3255 ( .IN1(n2429), .IN2(n2430), .QN(P2_N5421) );
  NOR2X0 U3256 ( .QN(n2430), .IN1(n2431), .IN2(n2432) );
  NAND2X0 U3257 ( .IN1(n2433), .IN2(n2434), .QN(n2432) );
  NAND2X0 U3072 ( .IN1(n2253), .IN2(P2_N345), .QN(n2263) );
  AND2X1 U3073 ( .IN1(P2_N4881), .IN2(n2254), .Q(n2261) );
  NOR2X0 U3074 ( .QN(n2259), .IN1(n2265), .IN2(n2266) );
  NAND2X0 U3075 ( .IN1(n2267), .IN2(n2268), .QN(n2266) );
  NAND2X0 U3076 ( .IN1(n2168), .IN2(P2_N933), .QN(n2268) );
  NAND2X0 U3077 ( .IN1(P2_N4711), .IN2(n2161), .QN(n2267) );
  AND2X1 U3078 ( .IN1(n9505), .IN2(n6589), .Q(n2265) );
  NAND2X0 U3079 ( .IN1(n2269), .IN2(n2270), .QN(P2_N5437) );
  NOR2X0 U3080 ( .QN(n2270), .IN1(n2271), .IN2(n2272) );
  NAND2X0 U3081 ( .IN1(n2273), .IN2(n2274), .QN(n2272) );
  NAND2X0 U3082 ( .IN1(P2_N4860), .IN2(n2252), .QN(n2274) );
  NAND2X0 U3083 ( .IN1(n2253), .IN2(P2_N346), .QN(n2273) );
  AND2X1 U3084 ( .IN1(P2_N4880), .IN2(n2254), .Q(n2271) );
  NOR2X0 U3085 ( .QN(n2269), .IN1(n2275), .IN2(n2276) );
  NAND2X0 U3086 ( .IN1(n2277), .IN2(n2278), .QN(n2276) );
  NAND2X0 U3087 ( .IN1(n2168), .IN2(P2_N932), .QN(n2278) );
  NAND2X0 U3088 ( .IN1(P2_N4710), .IN2(n2161), .QN(n2277) );
  AND2X1 U3089 ( .IN1(n9509), .IN2(n6589), .Q(n2275) );
  NAND2X0 U3090 ( .IN1(n2279), .IN2(n2280), .QN(P2_N5436) );
  NOR2X0 U3091 ( .QN(n2280), .IN1(n2281), .IN2(n2282) );
  NAND2X0 U3092 ( .IN1(n2283), .IN2(n2284), .QN(n2282) );
  NAND2X0 U3093 ( .IN1(P2_N4859), .IN2(n2252), .QN(n2284) );
  NAND2X0 U3094 ( .IN1(n2253), .IN2(P2_N347), .QN(n2283) );
  AND2X1 U3095 ( .IN1(P2_N4879), .IN2(n2254), .Q(n2281) );
  NOR2X0 U3096 ( .QN(n2279), .IN1(n2285), .IN2(n2286) );
  NAND2X0 U3097 ( .IN1(n2287), .IN2(n2288), .QN(n2286) );
  NAND2X0 U3098 ( .IN1(n2168), .IN2(P2_N931), .QN(n2288) );
  NAND2X0 U3099 ( .IN1(P2_N4709), .IN2(n2161), .QN(n2287) );
  AND2X1 U3100 ( .IN1(n9513), .IN2(n2166), .Q(n2285) );
  NAND2X0 U3101 ( .IN1(n2289), .IN2(n2290), .QN(P2_N5435) );
  NOR2X0 U3102 ( .QN(n2290), .IN1(n2291), .IN2(n2292) );
  NAND2X0 U3103 ( .IN1(n2293), .IN2(n2294), .QN(n2292) );
  NAND2X0 U3104 ( .IN1(P2_N4858), .IN2(n2252), .QN(n2294) );
  NAND2X0 U3105 ( .IN1(n2253), .IN2(P2_N348), .QN(n2293) );
  AND2X1 U3106 ( .IN1(P2_N4878), .IN2(n2254), .Q(n2291) );
  NOR2X0 U3107 ( .QN(n2289), .IN1(n2295), .IN2(n2296) );
  NAND2X0 U3108 ( .IN1(n2297), .IN2(n2298), .QN(n2296) );
  NAND2X0 U3109 ( .IN1(n2168), .IN2(P2_N930), .QN(n2298) );
  NAND2X0 U3110 ( .IN1(P2_N4708), .IN2(n2161), .QN(n2297) );
  AND2X1 U3111 ( .IN1(n9517), .IN2(n2166), .Q(n2295) );
  NAND2X0 U3112 ( .IN1(n2299), .IN2(n2300), .QN(P2_N5434) );
  NOR2X0 U3113 ( .QN(n2300), .IN1(n2301), .IN2(n2302) );
  NAND2X0 U3114 ( .IN1(n2303), .IN2(n2304), .QN(n2302) );
  NAND2X0 U3115 ( .IN1(P2_N4857), .IN2(n2252), .QN(n2304) );
  NAND2X0 U3116 ( .IN1(n2253), .IN2(P2_N349), .QN(n2303) );
  AND2X1 U3117 ( .IN1(P2_N4877), .IN2(n2254), .Q(n2301) );
  NOR2X0 U3118 ( .QN(n2299), .IN1(n2305), .IN2(n2306) );
  NAND2X0 U3119 ( .IN1(n2307), .IN2(n2308), .QN(n2306) );
  NAND2X0 U3120 ( .IN1(n2168), .IN2(P2_N929), .QN(n2308) );
  NAND2X0 U3121 ( .IN1(P2_N4707), .IN2(n2161), .QN(n2307) );
  AND2X1 U3122 ( .IN1(n9521), .IN2(n2166), .Q(n2305) );
  NAND2X0 U3123 ( .IN1(n2309), .IN2(n2310), .QN(P2_N5433) );
  NOR2X0 U3124 ( .QN(n2310), .IN1(n2311), .IN2(n2312) );
  NAND2X0 U3125 ( .IN1(n2313), .IN2(n2314), .QN(n2312) );
  NAND2X0 U3126 ( .IN1(P2_N4856), .IN2(n2252), .QN(n2314) );
  NAND2X0 U3127 ( .IN1(n2253), .IN2(P2_N350), .QN(n2313) );
  AND2X1 U3128 ( .IN1(P2_N4876), .IN2(n2254), .Q(n2311) );
  NOR2X0 U3129 ( .QN(n2309), .IN1(n2315), .IN2(n2316) );
  NAND2X0 U3130 ( .IN1(n2317), .IN2(n2318), .QN(n2316) );
  NAND2X0 U3131 ( .IN1(n2168), .IN2(P2_N928), .QN(n2318) );
  NAND2X0 U3132 ( .IN1(P2_N4706), .IN2(n2161), .QN(n2317) );
  AND2X1 U3133 ( .IN1(n9525), .IN2(n2166), .Q(n2315) );
  NAND2X0 U3134 ( .IN1(n2319), .IN2(n2320), .QN(P2_N5432) );
  NOR2X0 U3135 ( .QN(n2320), .IN1(n2321), .IN2(n2322) );
  NAND2X0 U3136 ( .IN1(n2323), .IN2(n2324), .QN(n2322) );
  NAND2X0 U3137 ( .IN1(P2_N4855), .IN2(n2252), .QN(n2324) );
  NAND2X0 U3138 ( .IN1(n2253), .IN2(P2_N351), .QN(n2323) );
  AND2X1 U3139 ( .IN1(P2_N4875), .IN2(n2254), .Q(n2321) );
  NOR2X0 U3140 ( .QN(n2319), .IN1(n2325), .IN2(n2326) );
  NAND2X0 U3141 ( .IN1(n2327), .IN2(n2328), .QN(n2326) );
  NAND2X0 U3142 ( .IN1(n2168), .IN2(P2_N927), .QN(n2328) );
  NAND2X0 U3143 ( .IN1(P2_N4705), .IN2(n2161), .QN(n2327) );
  AND2X1 U3144 ( .IN1(n9529), .IN2(n2166), .Q(n2325) );
  NAND2X0 U3145 ( .IN1(n2329), .IN2(n2330), .QN(P2_N5431) );
  NOR2X0 U3146 ( .QN(n2330), .IN1(n2331), .IN2(n2332) );
  NAND2X0 U3147 ( .IN1(n2333), .IN2(n2334), .QN(n2332) );
  NAND2X0 U3148 ( .IN1(P2_N4854), .IN2(n2252), .QN(n2334) );
  NAND2X0 U3149 ( .IN1(n2253), .IN2(P2_N352), .QN(n2333) );
  AND2X1 U3150 ( .IN1(P2_N4874), .IN2(n2254), .Q(n2331) );
  NOR2X0 U3151 ( .QN(n2329), .IN1(n2335), .IN2(n2336) );
  NAND2X0 U3152 ( .IN1(n2337), .IN2(n2338), .QN(n2336) );
  NAND2X0 U3153 ( .IN1(n2168), .IN2(P2_N926), .QN(n2338) );
  NAND2X0 U3154 ( .IN1(P2_N4704), .IN2(n2161), .QN(n2337) );
  AND2X1 U3155 ( .IN1(n9533), .IN2(n2166), .Q(n2335) );
  NAND2X0 U3156 ( .IN1(n2339), .IN2(n2340), .QN(P2_N5430) );
  NOR2X0 U3157 ( .QN(n2340), .IN1(n2341), .IN2(n2342) );
  NAND2X0 U3158 ( .IN1(n2343), .IN2(n2344), .QN(n2342) );
  NAND2X0 U3159 ( .IN1(P2_N4853), .IN2(n2252), .QN(n2344) );
  NAND2X0 U3160 ( .IN1(n2253), .IN2(P2_N353), .QN(n2343) );
  AND2X1 U3161 ( .IN1(P2_N4873), .IN2(n2254), .Q(n2341) );
  NOR2X0 U3162 ( .QN(n2339), .IN1(n2345), .IN2(n2346) );
  NAND2X0 U3163 ( .IN1(n2347), .IN2(n2348), .QN(n2346) );
  NAND2X0 U3164 ( .IN1(n2168), .IN2(P2_N925), .QN(n2348) );
  NAND2X0 U2979 ( .IN1(n2193), .IN2(n6589), .QN(n2192) );
  NAND2X0 U2980 ( .IN1(P2_N126), .IN2(n6588), .QN(n2191) );
  NAND2X0 U2981 ( .IN1(n2194), .IN2(n2195), .QN(P2_N5466) );
  NAND2X0 U2982 ( .IN1(n2196), .IN2(n6589), .QN(n2195) );
  NAND2X0 U2983 ( .IN1(P2_N125), .IN2(n6586), .QN(n2194) );
  NAND2X0 U2984 ( .IN1(n2197), .IN2(n2198), .QN(P2_N5465) );
  NAND2X0 U2985 ( .IN1(n2199), .IN2(n6589), .QN(n2198) );
  NAND2X0 U2986 ( .IN1(P2_N124), .IN2(n6586), .QN(n2197) );
  NAND2X0 U2987 ( .IN1(n2200), .IN2(n2201), .QN(P2_N5464) );
  NAND2X0 U2988 ( .IN1(n2202), .IN2(n6589), .QN(n2201) );
  NAND2X0 U2989 ( .IN1(P2_N123), .IN2(n6586), .QN(n2200) );
  NAND2X0 U2990 ( .IN1(n2203), .IN2(n2204), .QN(P2_N5463) );
  NAND2X0 U2991 ( .IN1(n2205), .IN2(n6589), .QN(n2204) );
  NAND2X0 U2992 ( .IN1(P2_N122), .IN2(n6586), .QN(n2203) );
  NAND2X0 U2993 ( .IN1(n2206), .IN2(n2207), .QN(P2_N5462) );
  NAND2X0 U2994 ( .IN1(n2008), .IN2(n6585), .QN(n2207) );
  NAND2X0 U2995 ( .IN1(P2_N121), .IN2(n6586), .QN(n2206) );
  NAND2X0 U2996 ( .IN1(n2208), .IN2(n2209), .QN(P2_N5461) );
  NAND2X0 U2997 ( .IN1(n2011), .IN2(n6585), .QN(n2209) );
  NAND2X0 U2998 ( .IN1(P2_N120), .IN2(n6586), .QN(n2208) );
  NAND2X0 U2999 ( .IN1(n2210), .IN2(n2211), .QN(P2_N5460) );
  NAND2X0 U3000 ( .IN1(n2014), .IN2(n6585), .QN(n2211) );
  NAND2X0 U3001 ( .IN1(P2_N119), .IN2(n6586), .QN(n2210) );
  NAND2X0 U3005 ( .IN1(n2212), .IN2(n2213), .QN(P2_N5459) );
  NAND2X0 U3006 ( .IN1(n2017), .IN2(n6585), .QN(n2213) );
  NAND2X0 U3007 ( .IN1(P2_N118), .IN2(n6586), .QN(n2212) );
  NAND2X0 U3008 ( .IN1(n2214), .IN2(n2215), .QN(P2_N5458) );
  NAND2X0 U3009 ( .IN1(n2020), .IN2(n6585), .QN(n2215) );
  NAND2X0 U3010 ( .IN1(P2_N117), .IN2(n6586), .QN(n2214) );
  NAND2X0 U3011 ( .IN1(n2216), .IN2(n2217), .QN(P2_N5457) );
  NAND2X0 U3012 ( .IN1(n2023), .IN2(n6585), .QN(n2217) );
  NAND2X0 U3013 ( .IN1(P2_N116), .IN2(n6586), .QN(n2216) );
  NAND2X0 U3014 ( .IN1(n2218), .IN2(n2219), .QN(P2_N5456) );
  NAND2X0 U3015 ( .IN1(n2026), .IN2(n6585), .QN(n2219) );
  NAND2X0 U3016 ( .IN1(P2_N115), .IN2(n6586), .QN(n2218) );
  NAND2X0 U3017 ( .IN1(n2220), .IN2(n2221), .QN(P2_N5454) );
  NAND2X0 U3018 ( .IN1(n2029), .IN2(n6585), .QN(n2221) );
  NAND2X0 U3019 ( .IN1(P2_N114), .IN2(n6586), .QN(n2220) );
  NAND2X0 U3020 ( .IN1(n2222), .IN2(n2223), .QN(P2_N5453) );
  NAND2X0 U3021 ( .IN1(n2032), .IN2(n6585), .QN(n2223) );
  NAND2X0 U3022 ( .IN1(P2_N113), .IN2(n6586), .QN(n2222) );
  NAND2X0 U3023 ( .IN1(n2224), .IN2(n2225), .QN(P2_N5452) );
  NAND2X0 U3024 ( .IN1(n2035), .IN2(n6585), .QN(n2225) );
  NAND2X0 U3025 ( .IN1(P2_N112), .IN2(n6586), .QN(n2224) );
  NAND2X0 U3026 ( .IN1(n2226), .IN2(n2227), .QN(P2_N5451) );
  NAND2X0 U3027 ( .IN1(n2038), .IN2(n6585), .QN(n2227) );
  NAND2X0 U3028 ( .IN1(P2_N111), .IN2(n6586), .QN(n2226) );
  NAND2X0 U3029 ( .IN1(n2228), .IN2(n2229), .QN(P2_N5450) );
  NAND2X0 U3030 ( .IN1(n2041), .IN2(n6585), .QN(n2229) );
  NAND2X0 U3031 ( .IN1(P2_N110), .IN2(n6586), .QN(n2228) );
  NAND2X0 U3032 ( .IN1(n2230), .IN2(n2231), .QN(P2_N5449) );
  NAND2X0 U3033 ( .IN1(n2044), .IN2(n6585), .QN(n2231) );
  NAND2X0 U3034 ( .IN1(P2_N109), .IN2(n6586), .QN(n2230) );
  NAND2X0 U3035 ( .IN1(n2232), .IN2(n2233), .QN(P2_N5448) );
  NAND2X0 U3036 ( .IN1(n2047), .IN2(n6585), .QN(n2233) );
  NAND2X0 U3037 ( .IN1(P2_N108), .IN2(n6586), .QN(n2232) );
  NAND2X0 U3038 ( .IN1(n2234), .IN2(n2235), .QN(P2_N5447) );
  NAND2X0 U3039 ( .IN1(n2050), .IN2(n6585), .QN(n2235) );
  NAND2X0 U3040 ( .IN1(P2_N107), .IN2(n6586), .QN(n2234) );
  NAND2X0 U3041 ( .IN1(n2236), .IN2(n2237), .QN(P2_N5446) );
  NAND2X0 U3042 ( .IN1(n2053), .IN2(n6585), .QN(n2237) );
  NAND2X0 U3043 ( .IN1(P2_N106), .IN2(n6586), .QN(n2236) );
  NAND2X0 U3044 ( .IN1(n2238), .IN2(n2239), .QN(P2_N5445) );
  NAND2X0 U3045 ( .IN1(n2056), .IN2(n6585), .QN(n2239) );
  NAND2X0 U3046 ( .IN1(P2_N105), .IN2(n6586), .QN(n2238) );
  NAND2X0 U3047 ( .IN1(n2240), .IN2(n2241), .QN(P2_N5444) );
  NAND2X0 U3048 ( .IN1(n2059), .IN2(n6585), .QN(n2241) );
  NAND2X0 U3049 ( .IN1(P2_N104), .IN2(n6586), .QN(n2240) );
  NAND2X0 U3050 ( .IN1(n2242), .IN2(n2243), .QN(P2_N5443) );
  NAND2X0 U3051 ( .IN1(n2062), .IN2(n6585), .QN(n2243) );
  NAND2X0 U3052 ( .IN1(P2_N103), .IN2(n6586), .QN(n2242) );
  NAND2X0 U3053 ( .IN1(n2244), .IN2(n2245), .QN(P2_N5442) );
  NAND2X0 U3054 ( .IN1(n2065), .IN2(n6585), .QN(n2245) );
  NAND2X0 U3055 ( .IN1(n6595), .IN2(n6586), .QN(n2244) );
  NAND2X0 U3057 ( .IN1(n2246), .IN2(n2247), .QN(P2_N5439) );
  NOR2X0 U3058 ( .QN(n2247), .IN1(n2248), .IN2(n2249) );
  NAND2X0 U3059 ( .IN1(n2250), .IN2(n2251), .QN(n2249) );
  NAND2X0 U3060 ( .IN1(P2_N4862), .IN2(n2252), .QN(n2251) );
  NAND2X0 U3061 ( .IN1(n2253), .IN2(P2_N344), .QN(n2250) );
  AND2X1 U3062 ( .IN1(P2_N4882), .IN2(n2254), .Q(n2248) );
  NOR2X0 U3063 ( .QN(n2246), .IN1(n2255), .IN2(n2256) );
  NAND2X0 U3064 ( .IN1(n2257), .IN2(n2258), .QN(n2256) );
  NAND2X0 U3065 ( .IN1(n2168), .IN2(P2_N934), .QN(n2258) );
  NAND2X0 U3066 ( .IN1(P2_N4712), .IN2(n2161), .QN(n2257) );
  AND2X1 U3067 ( .IN1(n9501), .IN2(n6589), .Q(n2255) );
  NAND2X0 U3068 ( .IN1(n2259), .IN2(n2260), .QN(P2_N5438) );
  NOR2X0 U3069 ( .QN(n2260), .IN1(n2261), .IN2(n2262) );
  NAND2X0 U3070 ( .IN1(n2263), .IN2(n2264), .QN(n2262) );
  NAND2X0 U3071 ( .IN1(P2_N4861), .IN2(n2252), .QN(n2264) );
  INVX0 U2885 ( .ZN(n2130), .INP(n7395) );
  NOR2X0 U2886 ( .QN(P2_N659), .IN1(n7329), .IN2(n7007) );
  NOR2X0 U2887 ( .QN(P2_N658), .IN1(n7013), .IN2(n7327) );
  NOR2X0 U2888 ( .QN(P2_N657), .IN1(n7015), .IN2(n7325) );
  NOR2X0 U2889 ( .QN(P2_N656), .IN1(n7015), .IN2(n7323) );
  NOR2X0 U2890 ( .QN(P2_N655), .IN1(n7015), .IN2(n7321) );
  NOR2X0 U2891 ( .QN(P2_N654), .IN1(n7015), .IN2(n7319) );
  NOR2X0 U2892 ( .QN(P2_N653), .IN1(n7015), .IN2(n7317) );
  NOR2X0 U2893 ( .QN(P2_N652), .IN1(n7015), .IN2(n7315) );
  NOR2X0 U2894 ( .QN(P2_N651), .IN1(n7013), .IN2(n7313) );
  NOR2X0 U2895 ( .QN(P2_N650), .IN1(n7013), .IN2(n7311) );
  NAND2X0 U2897 ( .IN1(n2006), .IN2(n2133), .QN(P2_N649) );
  NAND2X0 U2898 ( .IN1(P2_N914), .IN2(n2008), .QN(n2133) );
  NAND2X0 U2899 ( .IN1(n2009), .IN2(n2134), .QN(P2_N648) );
  NAND2X0 U2900 ( .IN1(P2_N914), .IN2(n2011), .QN(n2134) );
  NAND2X0 U2901 ( .IN1(n2012), .IN2(n2135), .QN(P2_N647) );
  NAND2X0 U2902 ( .IN1(P2_N914), .IN2(n2014), .QN(n2135) );
  NAND2X0 U2903 ( .IN1(n2015), .IN2(n2136), .QN(P2_N646) );
  NAND2X0 U2904 ( .IN1(P2_N914), .IN2(n2017), .QN(n2136) );
  NAND2X0 U2905 ( .IN1(n2018), .IN2(n2137), .QN(P2_N645) );
  NAND2X0 U2906 ( .IN1(n7009), .IN2(n2020), .QN(n2137) );
  NAND2X0 U2907 ( .IN1(n2021), .IN2(n2138), .QN(P2_N644) );
  NAND2X0 U2908 ( .IN1(n7009), .IN2(n2023), .QN(n2138) );
  NAND2X0 U2909 ( .IN1(n2024), .IN2(n2139), .QN(P2_N643) );
  NAND2X0 U2910 ( .IN1(n7009), .IN2(n2026), .QN(n2139) );
  NAND2X0 U2911 ( .IN1(n2027), .IN2(n2140), .QN(P2_N642) );
  NAND2X0 U2912 ( .IN1(n7010), .IN2(n2029), .QN(n2140) );
  NAND2X0 U2913 ( .IN1(n2030), .IN2(n2141), .QN(P2_N641) );
  NAND2X0 U2914 ( .IN1(n7010), .IN2(n2032), .QN(n2141) );
  NAND2X0 U2915 ( .IN1(n2033), .IN2(n2142), .QN(P2_N640) );
  NAND2X0 U2916 ( .IN1(n7010), .IN2(n2035), .QN(n2142) );
  NAND2X0 U2917 ( .IN1(n2036), .IN2(n2143), .QN(P2_N639) );
  NAND2X0 U2918 ( .IN1(n7010), .IN2(n2038), .QN(n2143) );
  NAND2X0 U2919 ( .IN1(n2039), .IN2(n2144), .QN(P2_N638) );
  NAND2X0 U2920 ( .IN1(n7010), .IN2(n2041), .QN(n2144) );
  NAND2X0 U2921 ( .IN1(n2042), .IN2(n2145), .QN(P2_N637) );
  NAND2X0 U2922 ( .IN1(n7010), .IN2(n2044), .QN(n2145) );
  NAND2X0 U2923 ( .IN1(n2045), .IN2(n2146), .QN(P2_N636) );
  NAND2X0 U2924 ( .IN1(n7006), .IN2(n2047), .QN(n2146) );
  NAND2X0 U2925 ( .IN1(n2048), .IN2(n2147), .QN(P2_N635) );
  NAND2X0 U2926 ( .IN1(n7006), .IN2(n2050), .QN(n2147) );
  NAND2X0 U2927 ( .IN1(n2051), .IN2(n2148), .QN(P2_N634) );
  NAND2X0 U2928 ( .IN1(n7462), .IN2(n2053), .QN(n2148) );
  NAND2X0 U2929 ( .IN1(n2054), .IN2(n2149), .QN(P2_N633) );
  NAND2X0 U2930 ( .IN1(n7462), .IN2(n2056), .QN(n2149) );
  NAND2X0 U2931 ( .IN1(n2057), .IN2(n2150), .QN(P2_N632) );
  NAND2X0 U2932 ( .IN1(n7462), .IN2(n2059), .QN(n2150) );
  NAND2X0 U2933 ( .IN1(n2060), .IN2(n2151), .QN(P2_N631) );
  NAND2X0 U2934 ( .IN1(n7462), .IN2(n2062), .QN(n2151) );
  NAND2X0 U2935 ( .IN1(n2063), .IN2(n2152), .QN(P2_N630) );
  NAND2X0 U2936 ( .IN1(n7462), .IN2(n2065), .QN(n2152) );
  NAND2X0 U2939 ( .IN1(n7332), .IN2(n2153), .QN(P2_N584) );
  AND2X1 U2947 ( .IN1(P2_N4777), .IN2(n2161), .Q(P2_N5486) );
  AND2X1 U2948 ( .IN1(P2_N4744), .IN2(n2161), .Q(P2_N5485) );
  AND2X1 U2949 ( .IN1(P2_N4713), .IN2(n2161), .Q(P2_N5484) );
  NAND2X0 U2950 ( .IN1(n6928), .IN2(n2163), .QN(P2_N5483) );
  NAND2X0 U2951 ( .IN1(n2164), .IN2(n2165), .QN(n2163) );
  AND2X1 U2952 ( .IN1(n7334), .IN2(n7415), .Q(n2165) );
  NOR2X0 U2953 ( .QN(n2164), .IN1(n6589), .IN2(n7421) );
  AND2X1 U2955 ( .IN1(n2161), .IN2(P2_N536), .Q(P2_N5482) );
  AND2X1 U2956 ( .IN1(n2169), .IN2(P2_N4841), .Q(P2_N5476) );
  NAND2X0 U2957 ( .IN1(n2170), .IN2(n2171), .QN(P2_N5475) );
  NAND2X0 U2958 ( .IN1(n2172), .IN2(n6589), .QN(n2171) );
  NAND2X0 U2959 ( .IN1(P2_N133), .IN2(n6588), .QN(n2170) );
  NAND2X0 U2960 ( .IN1(n2173), .IN2(n2174), .QN(P2_N5474) );
  NAND2X0 U2961 ( .IN1(n2175), .IN2(n6589), .QN(n2174) );
  NAND2X0 U2962 ( .IN1(P2_N132), .IN2(n6588), .QN(n2173) );
  NAND2X0 U2963 ( .IN1(n2176), .IN2(n2177), .QN(P2_N5473) );
  NAND2X0 U2964 ( .IN1(n2178), .IN2(n6589), .QN(n2177) );
  NAND2X0 U2965 ( .IN1(P2_N131), .IN2(n6588), .QN(n2176) );
  NAND2X0 U2966 ( .IN1(n2179), .IN2(n2180), .QN(P2_N5472) );
  NAND2X0 U2967 ( .IN1(n2181), .IN2(n6589), .QN(n2180) );
  NAND2X0 U2968 ( .IN1(P2_N130), .IN2(n6588), .QN(n2179) );
  NAND2X0 U2969 ( .IN1(n2182), .IN2(n2183), .QN(P2_N5471) );
  NAND2X0 U2970 ( .IN1(n2184), .IN2(n6589), .QN(n2183) );
  NAND2X0 U2971 ( .IN1(P2_N129), .IN2(n6588), .QN(n2182) );
  NAND2X0 U2972 ( .IN1(n2185), .IN2(n2186), .QN(P2_N5469) );
  NAND2X0 U2973 ( .IN1(n2187), .IN2(n6589), .QN(n2186) );
  NAND2X0 U2974 ( .IN1(P2_N128), .IN2(n6588), .QN(n2185) );
  NAND2X0 U2975 ( .IN1(n2188), .IN2(n2189), .QN(P2_N5468) );
  NAND2X0 U2976 ( .IN1(n2190), .IN2(n6589), .QN(n2189) );
  NAND2X0 U2977 ( .IN1(P2_N127), .IN2(n6588), .QN(n2188) );
  NAND2X0 U2978 ( .IN1(n2191), .IN2(n2192), .QN(P2_N5467) );
  NAND2X0 U2785 ( .IN1(n7462), .IN2(n2065), .QN(n2064) );
  NAND2X0 U2788 ( .IN1(n2067), .IN2(n2068), .QN(P2_N841) );
  NAND2X0 U2789 ( .IN1(P2_N658), .IN2(n2069), .QN(n2068) );
  NAND2X0 U2790 ( .IN1(P2_N392), .IN2(P2_N5494), .QN(n2067) );
  NAND2X0 U2791 ( .IN1(n2071), .IN2(n2072), .QN(P2_N840) );
  NAND2X0 U2792 ( .IN1(P2_N657), .IN2(n2069), .QN(n2072) );
  NAND2X0 U2793 ( .IN1(P2_N391), .IN2(P2_N5494), .QN(n2071) );
  NAND2X0 U2794 ( .IN1(n2073), .IN2(n2074), .QN(P2_N839) );
  NAND2X0 U2795 ( .IN1(P2_N656), .IN2(n2069), .QN(n2074) );
  NAND2X0 U2796 ( .IN1(P2_N390), .IN2(P2_N5494), .QN(n2073) );
  NAND2X0 U2797 ( .IN1(n2075), .IN2(n2076), .QN(P2_N838) );
  NAND2X0 U2798 ( .IN1(P2_N655), .IN2(n2069), .QN(n2076) );
  NAND2X0 U2799 ( .IN1(P2_N389), .IN2(P2_N5494), .QN(n2075) );
  NAND2X0 U2800 ( .IN1(n2077), .IN2(n2078), .QN(P2_N837) );
  NAND2X0 U2801 ( .IN1(P2_N654), .IN2(n2069), .QN(n2078) );
  NAND2X0 U2802 ( .IN1(P2_N388), .IN2(P2_N5494), .QN(n2077) );
  NAND2X0 U2803 ( .IN1(n2079), .IN2(n2080), .QN(P2_N836) );
  NAND2X0 U2804 ( .IN1(P2_N653), .IN2(n2069), .QN(n2080) );
  NAND2X0 U2805 ( .IN1(P2_N387), .IN2(P2_N5494), .QN(n2079) );
  NAND2X0 U2806 ( .IN1(n2081), .IN2(n2082), .QN(P2_N835) );
  NAND2X0 U2807 ( .IN1(P2_N652), .IN2(n2069), .QN(n2082) );
  NAND2X0 U2808 ( .IN1(P2_N386), .IN2(P2_N5494), .QN(n2081) );
  NAND2X0 U2809 ( .IN1(n2083), .IN2(n2084), .QN(P2_N834) );
  NAND2X0 U2810 ( .IN1(P2_N651), .IN2(n2069), .QN(n2084) );
  NAND2X0 U2811 ( .IN1(P2_N385), .IN2(P2_N5494), .QN(n2083) );
  NAND2X0 U2812 ( .IN1(n2085), .IN2(n2086), .QN(P2_N833) );
  NAND2X0 U2813 ( .IN1(P2_N650), .IN2(n2069), .QN(n2086) );
  NAND2X0 U2814 ( .IN1(P2_N384), .IN2(P2_N5494), .QN(n2085) );
  NAND2X0 U2815 ( .IN1(n2087), .IN2(n2088), .QN(P2_N832) );
  NAND2X0 U2816 ( .IN1(n2069), .IN2(P2_N649), .QN(n2088) );
  NAND2X0 U2817 ( .IN1(P2_N383), .IN2(P2_N5494), .QN(n2087) );
  NAND2X0 U2818 ( .IN1(n2089), .IN2(n2090), .QN(P2_N831) );
  NAND2X0 U2819 ( .IN1(n2069), .IN2(P2_N648), .QN(n2090) );
  NAND2X0 U2820 ( .IN1(P2_N382), .IN2(P2_N5494), .QN(n2089) );
  NAND2X0 U2821 ( .IN1(n2091), .IN2(n2092), .QN(P2_N830) );
  NAND2X0 U2822 ( .IN1(n2069), .IN2(P2_N647), .QN(n2092) );
  NAND2X0 U2823 ( .IN1(P2_N381), .IN2(P2_N5494), .QN(n2091) );
  NAND2X0 U2824 ( .IN1(n2093), .IN2(n2094), .QN(P2_N829) );
  NAND2X0 U2825 ( .IN1(n2069), .IN2(P2_N646), .QN(n2094) );
  NAND2X0 U2826 ( .IN1(P2_N380), .IN2(P2_N5494), .QN(n2093) );
  NAND2X0 U2827 ( .IN1(n2095), .IN2(n2096), .QN(P2_N828) );
  NAND2X0 U2828 ( .IN1(n2069), .IN2(P2_N645), .QN(n2096) );
  NAND2X0 U2829 ( .IN1(P2_N379), .IN2(P2_N5494), .QN(n2095) );
  NAND2X0 U2830 ( .IN1(n2097), .IN2(n2098), .QN(P2_N827) );
  NAND2X0 U2831 ( .IN1(n2069), .IN2(P2_N644), .QN(n2098) );
  NAND2X0 U2832 ( .IN1(P2_N378), .IN2(P2_N5494), .QN(n2097) );
  NAND2X0 U2833 ( .IN1(n2099), .IN2(n2100), .QN(P2_N826) );
  NAND2X0 U2834 ( .IN1(n2069), .IN2(P2_N643), .QN(n2100) );
  NAND2X0 U2835 ( .IN1(P2_N377), .IN2(P2_N5494), .QN(n2099) );
  NAND2X0 U2836 ( .IN1(n2101), .IN2(n2102), .QN(P2_N825) );
  NAND2X0 U2837 ( .IN1(n2069), .IN2(P2_N642), .QN(n2102) );
  NAND2X0 U2838 ( .IN1(P2_N376), .IN2(P2_N5494), .QN(n2101) );
  NAND2X0 U2839 ( .IN1(n2103), .IN2(n2104), .QN(P2_N824) );
  NAND2X0 U2840 ( .IN1(n2069), .IN2(P2_N641), .QN(n2104) );
  NAND2X0 U2841 ( .IN1(P2_N375), .IN2(P2_N5494), .QN(n2103) );
  NAND2X0 U2842 ( .IN1(n2105), .IN2(n2106), .QN(P2_N823) );
  NAND2X0 U2843 ( .IN1(n2069), .IN2(P2_N640), .QN(n2106) );
  NAND2X0 U2844 ( .IN1(P2_N374), .IN2(P2_N5494), .QN(n2105) );
  NAND2X0 U2845 ( .IN1(n2107), .IN2(n2108), .QN(P2_N822) );
  NAND2X0 U2846 ( .IN1(n2069), .IN2(P2_N639), .QN(n2108) );
  NAND2X0 U2847 ( .IN1(P2_N373), .IN2(P2_N5494), .QN(n2107) );
  NAND2X0 U2848 ( .IN1(n2109), .IN2(n2110), .QN(P2_N821) );
  NAND2X0 U2849 ( .IN1(n2069), .IN2(P2_N638), .QN(n2110) );
  NAND2X0 U2850 ( .IN1(P2_N372), .IN2(P2_N5494), .QN(n2109) );
  NAND2X0 U2851 ( .IN1(n2111), .IN2(n2112), .QN(P2_N820) );
  NAND2X0 U2852 ( .IN1(n2069), .IN2(P2_N637), .QN(n2112) );
  NAND2X0 U2853 ( .IN1(P2_N371), .IN2(P2_N5494), .QN(n2111) );
  NAND2X0 U2854 ( .IN1(n2113), .IN2(n2114), .QN(P2_N819) );
  NAND2X0 U2855 ( .IN1(n2069), .IN2(P2_N636), .QN(n2114) );
  NAND2X0 U2856 ( .IN1(P2_N370), .IN2(P2_N5494), .QN(n2113) );
  NAND2X0 U2857 ( .IN1(n2115), .IN2(n2116), .QN(P2_N818) );
  NAND2X0 U2858 ( .IN1(n2069), .IN2(P2_N635), .QN(n2116) );
  NAND2X0 U2859 ( .IN1(P2_N369), .IN2(P2_N5494), .QN(n2115) );
  NAND2X0 U2860 ( .IN1(n2117), .IN2(n2118), .QN(P2_N817) );
  NAND2X0 U2861 ( .IN1(n2069), .IN2(P2_N634), .QN(n2118) );
  NAND2X0 U2862 ( .IN1(P2_N368), .IN2(P2_N5494), .QN(n2117) );
  NAND2X0 U2863 ( .IN1(n2119), .IN2(n2120), .QN(P2_N816) );
  NAND2X0 U2864 ( .IN1(n2069), .IN2(P2_N633), .QN(n2120) );
  NAND2X0 U2865 ( .IN1(n18813), .IN2(P2_N5494), .QN(n2119) );
  NAND2X0 U2866 ( .IN1(n2121), .IN2(n2122), .QN(P2_N815) );
  NAND2X0 U2867 ( .IN1(n2069), .IN2(P2_N632), .QN(n2122) );
  NAND2X0 U2868 ( .IN1(n6683), .IN2(P2_N5494), .QN(n2121) );
  NAND2X0 U2869 ( .IN1(n2123), .IN2(n2124), .QN(P2_N814) );
  NAND2X0 U2870 ( .IN1(n2069), .IN2(P2_N631), .QN(n2124) );
  NAND2X0 U2871 ( .IN1(n6682), .IN2(P2_N5494), .QN(n2123) );
  NAND2X0 U2872 ( .IN1(n2125), .IN2(n2126), .QN(P2_N813) );
  NAND2X0 U2873 ( .IN1(n2069), .IN2(P2_N630), .QN(n2126) );
  NAND2X0 U2876 ( .IN1(n6681), .IN2(P2_N5494), .QN(n2125) );
  NAND2X0 U2881 ( .IN1(n7395), .IN2(n2129), .QN(P2_N780) );
  NAND2X0 U2882 ( .IN1(n7396), .IN2(n2130), .QN(P2_N778) );
  NOR2X0 U2883 ( .QN(P2_N842), .IN1(n2130), .IN2(n2129) );
  INVX0 U2884 ( .ZN(n2129), .INP(n7396) );
  OR2X1 U1541 ( .IN2(P2_N342), .IN1(n7401), .Q(n1478) );
  NOR2X0 U1544 ( .QN(n1481), .IN1(n7341), .IN2(n7334) );
  OR2X2 U1545 ( .IN2(n1482), .IN1(P1_N4553), .Q(P1_N5584) );
  NAND2X0 U1546 ( .IN1(P1_N4370), .IN2(P1_N4372), .QN(n1482) );
  OR2X2 U1547 ( .IN2(n1483), .IN1(P1_N4180), .Q(P1_N5583) );
  NAND2X0 U1548 ( .IN1(P1_N3997), .IN2(P1_N3999), .QN(n1483) );
  OR2X2 U1549 ( .IN2(n1484), .IN1(P1_N3807), .Q(P1_N5582) );
  NAND2X0 U1550 ( .IN1(P1_N3624), .IN2(P1_N3626), .QN(n1484) );
  NAND2X0 U1552 ( .IN1(P1_N3251), .IN2(P1_N3253), .QN(n1485) );
  OR2X2 U1553 ( .IN2(n1486), .IN1(P1_N3061), .Q(P1_N5580) );
  NAND2X0 U1554 ( .IN1(P1_N2878), .IN2(P1_N2880), .QN(n1486) );
  OR2X2 U1555 ( .IN2(n1487), .IN1(P1_N2688), .Q(P1_N5579) );
  NAND2X0 U1556 ( .IN1(P1_N2505), .IN2(P1_N2507), .QN(n1487) );
  OR2X2 U1557 ( .IN2(n1488), .IN1(P1_N2315), .Q(P1_N5578) );
  NAND2X0 U1558 ( .IN1(P1_N2132), .IN2(P1_N2134), .QN(n1488) );
  OR2X1 U1559 ( .IN2(n1489), .IN1(P1_N1942), .Q(P1_N5577) );
  NAND2X0 U1560 ( .IN1(P1_N1759), .IN2(P1_N1761), .QN(n1489) );
  OR2X1 U1561 ( .IN2(n1490), .IN1(P1_N968), .Q(P1_N5576) );
  NAND2X0 U1562 ( .IN1(P1_N779), .IN2(P1_N781), .QN(n1490) );
  OR2X1 U1563 ( .IN2(n1491), .IN1(P1_N4816), .Q(P1_N5574) );
  NAND2X0 U1564 ( .IN1(P1_N4752), .IN2(P1_N4754), .QN(n1491) );
  OR2X1 U1565 ( .IN2(n1492), .IN1(P1_N1569), .Q(P1_N5573) );
  NAND2X0 U1566 ( .IN1(P1_N1505), .IN2(P1_N1507), .QN(n1492) );
  OR2X1 U1567 ( .IN2(n1493), .IN1(P1_N1314), .Q(P1_N5572) );
  NAND2X0 U1568 ( .IN1(P1_N1250), .IN2(P1_N1252), .QN(n1493) );
  AND2X1 U1570 ( .IN1(n1494), .IN2(n1495), .Q(P1_N499) );
  NAND2X0 U1571 ( .IN1(P1_N342), .IN2(n7403), .QN(n1495) );
  OR2X1 U1572 ( .IN2(P1_N342), .IN1(n7403), .Q(n1494) );
  NOR2X0 U1574 ( .QN(P1_N4971), .IN1(n1497), .IN2(n1498) );
  NOR2X0 U1575 ( .QN(n1498), .IN1(n1504), .IN2(n6730) );
  NOR2X0 U1576 ( .QN(n1497), .IN1(P1_N363), .IN2(n920) );
  INVX0 U1577 ( .ZN(n920), .INP(n1504) );
  NOR2X0 U1578 ( .QN(P1_N4970), .IN1(n1500), .IN2(n1501) );
  NOR2X0 U1579 ( .QN(n1501), .IN1(n1503), .IN2(n6730) );
  NOR2X0 U1581 ( .QN(n1500), .IN1(P1_N363), .IN2(n981) );
  INVX0 U1582 ( .ZN(n981), .INP(n1503) );
  NOR2X0 U1584 ( .QN(n1502), .IN1(n7340), .IN2(n7337) );
  NOR2X0 U2736 ( .QN(P2_N913), .IN1(n7327), .IN2(n7013) );
  NOR2X0 U2737 ( .QN(P2_N912), .IN1(n7325), .IN2(n7015) );
  NOR2X0 U2738 ( .QN(P2_N911), .IN1(n7323), .IN2(n7015) );
  NOR2X0 U2739 ( .QN(P2_N910), .IN1(n7321), .IN2(n7015) );
  NOR2X0 U2740 ( .QN(P2_N909), .IN1(n7319), .IN2(n7015) );
  NOR2X0 U2741 ( .QN(P2_N908), .IN1(n7317), .IN2(n7015) );
  NOR2X0 U2742 ( .QN(P2_N907), .IN1(n7315), .IN2(n7015) );
  NOR2X0 U2743 ( .QN(P2_N906), .IN1(n7313), .IN2(n7013) );
  NOR2X0 U2744 ( .QN(P2_N905), .IN1(n7311), .IN2(n7013) );
  NAND2X0 U2746 ( .IN1(n2006), .IN2(n2007), .QN(P2_N904) );
  NAND2X0 U2747 ( .IN1(P2_N914), .IN2(n2008), .QN(n2007) );
  NAND2X0 U2748 ( .IN1(n2009), .IN2(n2010), .QN(P2_N903) );
  NAND2X0 U2749 ( .IN1(P2_N914), .IN2(n2011), .QN(n2010) );
  NAND2X0 U2750 ( .IN1(n2012), .IN2(n2013), .QN(P2_N902) );
  NAND2X0 U2751 ( .IN1(P2_N914), .IN2(n2014), .QN(n2013) );
  NAND2X0 U2752 ( .IN1(n2015), .IN2(n2016), .QN(P2_N901) );
  NAND2X0 U2753 ( .IN1(P2_N914), .IN2(n2017), .QN(n2016) );
  NAND2X0 U2754 ( .IN1(n2018), .IN2(n2019), .QN(P2_N900) );
  NAND2X0 U2755 ( .IN1(n7009), .IN2(n2020), .QN(n2019) );
  NAND2X0 U2756 ( .IN1(n2021), .IN2(n2022), .QN(P2_N899) );
  NAND2X0 U2757 ( .IN1(n7009), .IN2(n2023), .QN(n2022) );
  NAND2X0 U2758 ( .IN1(n2024), .IN2(n2025), .QN(P2_N898) );
  NAND2X0 U2759 ( .IN1(n7009), .IN2(n2026), .QN(n2025) );
  NAND2X0 U2760 ( .IN1(n2027), .IN2(n2028), .QN(P2_N897) );
  NAND2X0 U2761 ( .IN1(n7010), .IN2(n2029), .QN(n2028) );
  NAND2X0 U2762 ( .IN1(n2030), .IN2(n2031), .QN(P2_N896) );
  NAND2X0 U2763 ( .IN1(n7010), .IN2(n2032), .QN(n2031) );
  NAND2X0 U2764 ( .IN1(n2033), .IN2(n2034), .QN(P2_N895) );
  NAND2X0 U2765 ( .IN1(n7010), .IN2(n2035), .QN(n2034) );
  NAND2X0 U2766 ( .IN1(n2036), .IN2(n2037), .QN(P2_N894) );
  NAND2X0 U2767 ( .IN1(n7010), .IN2(n2038), .QN(n2037) );
  NAND2X0 U2768 ( .IN1(n2039), .IN2(n2040), .QN(P2_N893) );
  NAND2X0 U2769 ( .IN1(n7010), .IN2(n2041), .QN(n2040) );
  NAND2X0 U2770 ( .IN1(n2042), .IN2(n2043), .QN(P2_N892) );
  NAND2X0 U2771 ( .IN1(n7010), .IN2(n2044), .QN(n2043) );
  NAND2X0 U2772 ( .IN1(n2045), .IN2(n2046), .QN(P2_N891) );
  NAND2X0 U2773 ( .IN1(n7006), .IN2(n2047), .QN(n2046) );
  NAND2X0 U2774 ( .IN1(n2048), .IN2(n2049), .QN(P2_N890) );
  NAND2X0 U2775 ( .IN1(n7006), .IN2(n2050), .QN(n2049) );
  NAND2X0 U2776 ( .IN1(n2051), .IN2(n2052), .QN(P2_N889) );
  NAND2X0 U2777 ( .IN1(n7462), .IN2(n2053), .QN(n2052) );
  NAND2X0 U2778 ( .IN1(n2054), .IN2(n2055), .QN(P2_N888) );
  NAND2X0 U2779 ( .IN1(n7462), .IN2(n2056), .QN(n2055) );
  NAND2X0 U2780 ( .IN1(n2057), .IN2(n2058), .QN(P2_N887) );
  NAND2X0 U2781 ( .IN1(n7462), .IN2(n2059), .QN(n2058) );
  NAND2X0 U2782 ( .IN1(n2060), .IN2(n2061), .QN(P2_N886) );
  NAND2X0 U2783 ( .IN1(n7462), .IN2(n2062), .QN(n2061) );
  NAND2X0 U2784 ( .IN1(n2063), .IN2(n2064), .QN(P2_N885) );
  NAND2X0 U1448 ( .IN1(P2_N5462), .IN2(P2_N5470), .QN(n1423) );
  NAND2X0 U1449 ( .IN1(n6729), .IN2(n6611), .QN(n1422) );
  NAND2X0 U1450 ( .IN1(n1424), .IN2(n1425), .QN(n6298) );
  NAND2X0 U1451 ( .IN1(P2_N5461), .IN2(P2_N5470), .QN(n1425) );
  NAND2X0 U1452 ( .IN1(n6729), .IN2(n6612), .QN(n1424) );
  NAND2X0 U1453 ( .IN1(n1426), .IN2(n1427), .QN(n6299) );
  NAND2X0 U1454 ( .IN1(P2_N5460), .IN2(P2_N5470), .QN(n1427) );
  NAND2X0 U1455 ( .IN1(n6729), .IN2(n6613), .QN(n1426) );
  NAND2X0 U1456 ( .IN1(n1428), .IN2(n1429), .QN(n6300) );
  NAND2X0 U1457 ( .IN1(P2_N5459), .IN2(P2_N5470), .QN(n1429) );
  NAND2X0 U1458 ( .IN1(n6729), .IN2(n6614), .QN(n1428) );
  NAND2X0 U1459 ( .IN1(n1430), .IN2(n1431), .QN(n6301) );
  NAND2X0 U1460 ( .IN1(P2_N5458), .IN2(P2_N5470), .QN(n1431) );
  NAND2X0 U1461 ( .IN1(n6729), .IN2(n6615), .QN(n1430) );
  NAND2X0 U1462 ( .IN1(n1432), .IN2(n1433), .QN(n6302) );
  NAND2X0 U1463 ( .IN1(P2_N5457), .IN2(P2_N5470), .QN(n1433) );
  NAND2X0 U1464 ( .IN1(n6729), .IN2(n6616), .QN(n1432) );
  NAND2X0 U1465 ( .IN1(n1434), .IN2(n1435), .QN(n6303) );
  NAND2X0 U1466 ( .IN1(P2_N5456), .IN2(P2_N5470), .QN(n1435) );
  NAND2X0 U1467 ( .IN1(n6729), .IN2(n6617), .QN(n1434) );
  NAND2X0 U1468 ( .IN1(n1436), .IN2(n1437), .QN(n6304) );
  NAND2X0 U1469 ( .IN1(P2_N5454), .IN2(P2_N5470), .QN(n1437) );
  NAND2X0 U1470 ( .IN1(n6729), .IN2(n6607), .QN(n1436) );
  NAND2X0 U1471 ( .IN1(n1438), .IN2(n1439), .QN(n6305) );
  NAND2X0 U1472 ( .IN1(P2_N5453), .IN2(P2_N5470), .QN(n1439) );
  NAND2X0 U1473 ( .IN1(n6729), .IN2(n6606), .QN(n1438) );
  NAND2X0 U1474 ( .IN1(n1440), .IN2(n1441), .QN(n6306) );
  NAND2X0 U1475 ( .IN1(P2_N5452), .IN2(P2_N5470), .QN(n1441) );
  NAND2X0 U1476 ( .IN1(n6729), .IN2(n6605), .QN(n1440) );
  NAND2X0 U1477 ( .IN1(n1442), .IN2(n1443), .QN(n6307) );
  NAND2X0 U1478 ( .IN1(P2_N5451), .IN2(P2_N5470), .QN(n1443) );
  NAND2X0 U1479 ( .IN1(n6729), .IN2(n6604), .QN(n1442) );
  NAND2X0 U1480 ( .IN1(n1444), .IN2(n1445), .QN(n6308) );
  NAND2X0 U1481 ( .IN1(P2_N5450), .IN2(P2_N5470), .QN(n1445) );
  NAND2X0 U1482 ( .IN1(n6729), .IN2(n6603), .QN(n1444) );
  NAND2X0 U1483 ( .IN1(n1446), .IN2(n1447), .QN(n6309) );
  NAND2X0 U1484 ( .IN1(P2_N5449), .IN2(P2_N5470), .QN(n1447) );
  NAND2X0 U1485 ( .IN1(n6729), .IN2(n6602), .QN(n1446) );
  NAND2X0 U1486 ( .IN1(n1448), .IN2(n1449), .QN(n6310) );
  NAND2X0 U1487 ( .IN1(P2_N5448), .IN2(P2_N5470), .QN(n1449) );
  NAND2X0 U1488 ( .IN1(n6729), .IN2(n6601), .QN(n1448) );
  NAND2X0 U1489 ( .IN1(n1450), .IN2(n1451), .QN(n6311) );
  NAND2X0 U1490 ( .IN1(P2_N5447), .IN2(P2_N5470), .QN(n1451) );
  NAND2X0 U1491 ( .IN1(n6729), .IN2(n6600), .QN(n1450) );
  NAND2X0 U1492 ( .IN1(n1452), .IN2(n1453), .QN(n6312) );
  NAND2X0 U1493 ( .IN1(P2_N5446), .IN2(P2_N5470), .QN(n1453) );
  NAND2X0 U1494 ( .IN1(n6729), .IN2(n6599), .QN(n1452) );
  NAND2X0 U1495 ( .IN1(n1454), .IN2(n1455), .QN(n6313) );
  NAND2X0 U1496 ( .IN1(P2_N5445), .IN2(P2_N5470), .QN(n1455) );
  NAND2X0 U1497 ( .IN1(n6729), .IN2(n6598), .QN(n1454) );
  NAND2X0 U1498 ( .IN1(n1456), .IN2(n1457), .QN(n6314) );
  NAND2X0 U1499 ( .IN1(P2_N5444), .IN2(P2_N5470), .QN(n1457) );
  NAND2X0 U1500 ( .IN1(n6729), .IN2(n6597), .QN(n1456) );
  NAND2X0 U1501 ( .IN1(n1458), .IN2(n1459), .QN(n6315) );
  NAND2X0 U1502 ( .IN1(P2_N5443), .IN2(P2_N5470), .QN(n1459) );
  NAND2X0 U1503 ( .IN1(n6729), .IN2(n6596), .QN(n1458) );
  NAND2X0 U1504 ( .IN1(n1460), .IN2(n1461), .QN(n6316) );
  NAND2X0 U1505 ( .IN1(P2_N5442), .IN2(P2_N5470), .QN(n1461) );
  NAND2X0 U1506 ( .IN1(n6729), .IN2(n6595), .QN(n1460) );
  NAND2X0 U1507 ( .IN1(n1462), .IN2(n1463), .QN(n6317) );
  NAND2X0 U1508 ( .IN1(n6729), .IN2(n10137), .QN(n1463) );
  NAND2X0 U1509 ( .IN1(P2_N5474), .IN2(P2_N5470), .QN(n1462) );
  NAND2X0 U1510 ( .IN1(n1464), .IN2(n1465), .QN(n6318) );
  NAND2X0 U1511 ( .IN1(n6729), .IN2(n6688), .QN(n1465) );
  NAND2X0 U1513 ( .IN1(P2_N5475), .IN2(P2_N5470), .QN(n1464) );
  NOR2X0 U1515 ( .QN(n1466), .IN1(P2_N4398), .IN2(n7397) );
  OR2X1 U1516 ( .IN2(n1467), .IN1(P2_N4054), .Q(P2_N5508) );
  NAND2X0 U1517 ( .IN1(P2_N3871), .IN2(P2_N3873), .QN(n1467) );
  OR2X1 U1518 ( .IN2(n1468), .IN1(P2_N3681), .Q(P2_N5507) );
  NAND2X0 U1519 ( .IN1(P2_N3498), .IN2(P2_N3500), .QN(n1468) );
  OR2X1 U1520 ( .IN2(n1469), .IN1(P2_N3308), .Q(P2_N5506) );
  NAND2X0 U1521 ( .IN1(P2_N3125), .IN2(P2_N3127), .QN(n1469) );
  OR2X1 U1522 ( .IN2(n1470), .IN1(P2_N2935), .Q(P2_N5505) );
  NAND2X0 U1523 ( .IN1(P2_N2752), .IN2(P2_N2754), .QN(n1470) );
  OR2X1 U1524 ( .IN2(n1471), .IN1(P2_N2562), .Q(P2_N5504) );
  NAND2X0 U1525 ( .IN1(P2_N2379), .IN2(P2_N2381), .QN(n1471) );
  OR2X1 U1526 ( .IN2(n1472), .IN1(P2_N2189), .Q(P2_N5503) );
  NAND2X0 U1527 ( .IN1(P2_N2006), .IN2(P2_N2008), .QN(n1472) );
  OR2X1 U1528 ( .IN2(n1473), .IN1(P2_N1816), .Q(P2_N5502) );
  NAND2X0 U1529 ( .IN1(P2_N1633), .IN2(P2_N1635), .QN(n1473) );
  NOR2X0 U1531 ( .QN(n1474), .IN1(P2_N4661), .IN2(n7402) );
  OR2X1 U1532 ( .IN2(n1475), .IN1(P2_N1443), .Q(P2_N5496) );
  NAND2X0 U1533 ( .IN1(P2_N1379), .IN2(P2_N1381), .QN(n1475) );
  OR2X1 U1534 ( .IN2(n1476), .IN1(P2_N1188), .Q(P2_N5495) );
  NAND2X0 U1535 ( .IN1(P2_N1124), .IN2(P2_N1126), .QN(n1476) );
  OR2X1 U1536 ( .IN2(n1477), .IN1(P2_N842), .Q(P2_N5494) );
  NAND2X0 U1537 ( .IN1(P2_N778), .IN2(P2_N780), .QN(n1477) );
  AND2X1 U1539 ( .IN1(n1478), .IN2(n1479), .Q(P2_N499) );
  NAND2X0 U1540 ( .IN1(P2_N342), .IN2(n7401), .QN(n1479) );
  NAND2X0 U1355 ( .IN1(n7291), .IN2(n9126), .QN(n1360) );
  NAND2X0 U1356 ( .IN1(n1362), .IN2(n1363), .QN(n6267) );
  NAND2X0 U1357 ( .IN1(P2_N4767), .IN2(P2_N5484), .QN(n1363) );
  NAND2X0 U1358 ( .IN1(n7291), .IN2(n9130), .QN(n1362) );
  NAND2X0 U1359 ( .IN1(n1364), .IN2(n1365), .QN(n6268) );
  NAND2X0 U1360 ( .IN1(P2_N4766), .IN2(P2_N5484), .QN(n1365) );
  NAND2X0 U1361 ( .IN1(n7291), .IN2(n9134), .QN(n1364) );
  NAND2X0 U1362 ( .IN1(n1366), .IN2(n1367), .QN(n6269) );
  NAND2X0 U1363 ( .IN1(P2_N4765), .IN2(P2_N5484), .QN(n1367) );
  NAND2X0 U1364 ( .IN1(n7291), .IN2(n9138), .QN(n1366) );
  NAND2X0 U1365 ( .IN1(n1368), .IN2(n1369), .QN(n6270) );
  NAND2X0 U1366 ( .IN1(P2_N4764), .IN2(P2_N5484), .QN(n1369) );
  NAND2X0 U1367 ( .IN1(n7291), .IN2(n9142), .QN(n1368) );
  NAND2X0 U1368 ( .IN1(n1370), .IN2(n1371), .QN(n6271) );
  NAND2X0 U1369 ( .IN1(P2_N4763), .IN2(P2_N5484), .QN(n1371) );
  NAND2X0 U1370 ( .IN1(n7291), .IN2(n9146), .QN(n1370) );
  NAND2X0 U1371 ( .IN1(n1372), .IN2(n1373), .QN(n6272) );
  NAND2X0 U1372 ( .IN1(P2_N4762), .IN2(P2_N5484), .QN(n1373) );
  NAND2X0 U1373 ( .IN1(n7291), .IN2(n9150), .QN(n1372) );
  NAND2X0 U1374 ( .IN1(n1374), .IN2(n1375), .QN(n6273) );
  NAND2X0 U1375 ( .IN1(P2_N4761), .IN2(P2_N5484), .QN(n1375) );
  NAND2X0 U1376 ( .IN1(n7291), .IN2(n9154), .QN(n1374) );
  NAND2X0 U1377 ( .IN1(n1376), .IN2(n1377), .QN(n6274) );
  NAND2X0 U1378 ( .IN1(P2_N4760), .IN2(P2_N5484), .QN(n1377) );
  NAND2X0 U1379 ( .IN1(n7291), .IN2(n9158), .QN(n1376) );
  NAND2X0 U1380 ( .IN1(n1378), .IN2(n1379), .QN(n6275) );
  NAND2X0 U1381 ( .IN1(P2_N4759), .IN2(P2_N5484), .QN(n1379) );
  NAND2X0 U1382 ( .IN1(n7291), .IN2(n9162), .QN(n1378) );
  NAND2X0 U1383 ( .IN1(n1380), .IN2(n1381), .QN(n6276) );
  NAND2X0 U1384 ( .IN1(P2_N4758), .IN2(P2_N5484), .QN(n1381) );
  NAND2X0 U1385 ( .IN1(n7291), .IN2(n9166), .QN(n1380) );
  NAND2X0 U1386 ( .IN1(n1382), .IN2(n1383), .QN(n6277) );
  NAND2X0 U1387 ( .IN1(P2_N4757), .IN2(P2_N5484), .QN(n1383) );
  NAND2X0 U1388 ( .IN1(n7291), .IN2(n9170), .QN(n1382) );
  NAND2X0 U1389 ( .IN1(n1384), .IN2(n1385), .QN(n6278) );
  NAND2X0 U1390 ( .IN1(P2_N4756), .IN2(P2_N5484), .QN(n1385) );
  NAND2X0 U1391 ( .IN1(n7291), .IN2(n9174), .QN(n1384) );
  NAND2X0 U1392 ( .IN1(n1386), .IN2(n1387), .QN(n6279) );
  NAND2X0 U1393 ( .IN1(P2_N4755), .IN2(P2_N5484), .QN(n1387) );
  NAND2X0 U1394 ( .IN1(n7291), .IN2(n9178), .QN(n1386) );
  NAND2X0 U1395 ( .IN1(n1388), .IN2(n1389), .QN(n6280) );
  NAND2X0 U1396 ( .IN1(P2_N4754), .IN2(P2_N5484), .QN(n1389) );
  NAND2X0 U1397 ( .IN1(n7291), .IN2(n9182), .QN(n1388) );
  NAND2X0 U1398 ( .IN1(n1390), .IN2(n1391), .QN(n6281) );
  NAND2X0 U1399 ( .IN1(P2_N4753), .IN2(P2_N5484), .QN(n1391) );
  NAND2X0 U1400 ( .IN1(n7291), .IN2(n9186), .QN(n1390) );
  NAND2X0 U1401 ( .IN1(n1392), .IN2(n1393), .QN(n6282) );
  NAND2X0 U1402 ( .IN1(P2_N4752), .IN2(P2_N5484), .QN(n1393) );
  NAND2X0 U1403 ( .IN1(n7291), .IN2(n9190), .QN(n1392) );
  NAND2X0 U1404 ( .IN1(n1394), .IN2(n1395), .QN(n6283) );
  NAND2X0 U1405 ( .IN1(P2_N4751), .IN2(P2_N5484), .QN(n1395) );
  NAND2X0 U1406 ( .IN1(n7291), .IN2(n9194), .QN(n1394) );
  NAND2X0 U1407 ( .IN1(n1396), .IN2(n1397), .QN(n6284) );
  NAND2X0 U1408 ( .IN1(P2_N4750), .IN2(P2_N5484), .QN(n1397) );
  NAND2X0 U1409 ( .IN1(n7291), .IN2(n9198), .QN(n1396) );
  NAND2X0 U1410 ( .IN1(n1398), .IN2(n1399), .QN(n6285) );
  NAND2X0 U1411 ( .IN1(P2_N4749), .IN2(P2_N5484), .QN(n1399) );
  NAND2X0 U1412 ( .IN1(n7291), .IN2(n9202), .QN(n1398) );
  NAND2X0 U1413 ( .IN1(n1400), .IN2(n1401), .QN(n6286) );
  NAND2X0 U1414 ( .IN1(P2_N4748), .IN2(P2_N5484), .QN(n1401) );
  NAND2X0 U1415 ( .IN1(n7291), .IN2(n9206), .QN(n1400) );
  NAND2X0 U1416 ( .IN1(n1402), .IN2(n1403), .QN(n6287) );
  NAND2X0 U1417 ( .IN1(P2_N4747), .IN2(P2_N5484), .QN(n1403) );
  NAND2X0 U1418 ( .IN1(n7291), .IN2(n9210), .QN(n1402) );
  NAND2X0 U1419 ( .IN1(n1404), .IN2(n1405), .QN(n6288) );
  NAND2X0 U1420 ( .IN1(P2_N4746), .IN2(P2_N5484), .QN(n1405) );
  NAND2X0 U1421 ( .IN1(n7291), .IN2(n9214), .QN(n1404) );
  NAND2X0 U1422 ( .IN1(n1406), .IN2(n1407), .QN(n6289) );
  NAND2X0 U1423 ( .IN1(P2_N4745), .IN2(P2_N5484), .QN(n1407) );
  NAND2X0 U1424 ( .IN1(n7291), .IN2(n9218), .QN(n1406) );
  NAND2X0 U1426 ( .IN1(n1408), .IN2(n1409), .QN(n6290) );
  NAND2X0 U1427 ( .IN1(P2_N5469), .IN2(P2_N5470), .QN(n1409) );
  NAND2X0 U1428 ( .IN1(n6729), .IN2(n10183), .QN(n1408) );
  NAND2X0 U1429 ( .IN1(n1410), .IN2(n1411), .QN(n6291) );
  NAND2X0 U1430 ( .IN1(P2_N5468), .IN2(P2_N5470), .QN(n1411) );
  NAND2X0 U1431 ( .IN1(n6729), .IN2(n10377), .QN(n1410) );
  NAND2X0 U1432 ( .IN1(n1412), .IN2(n1413), .QN(n6292) );
  NAND2X0 U1433 ( .IN1(P2_N5467), .IN2(P2_N5470), .QN(n1413) );
  NAND2X0 U1434 ( .IN1(n6729), .IN2(n10191), .QN(n1412) );
  NAND2X0 U1435 ( .IN1(n1414), .IN2(n1415), .QN(n6293) );
  NAND2X0 U1436 ( .IN1(P2_N5466), .IN2(P2_N5470), .QN(n1415) );
  NAND2X0 U1437 ( .IN1(n6729), .IN2(n6719), .QN(n1414) );
  NAND2X0 U1438 ( .IN1(n1416), .IN2(n1417), .QN(n6294) );
  NAND2X0 U1439 ( .IN1(P2_N5465), .IN2(P2_N5470), .QN(n1417) );
  NAND2X0 U1440 ( .IN1(n6729), .IN2(n6608), .QN(n1416) );
  NAND2X0 U1441 ( .IN1(n1418), .IN2(n1419), .QN(n6295) );
  NAND2X0 U1442 ( .IN1(P2_N5464), .IN2(P2_N5470), .QN(n1419) );
  NAND2X0 U1443 ( .IN1(n6729), .IN2(n6609), .QN(n1418) );
  NAND2X0 U1444 ( .IN1(n1420), .IN2(n1421), .QN(n6296) );
  NAND2X0 U1445 ( .IN1(P2_N5463), .IN2(P2_N5470), .QN(n1421) );
  NAND2X0 U1446 ( .IN1(n6729), .IN2(n6610), .QN(n1420) );
  NAND2X0 U1447 ( .IN1(n1422), .IN2(n1423), .QN(n6297) );
  NAND2X0 U1262 ( .IN1(n1300), .IN2(n1301), .QN(n6236) );
  NAND2X0 U1263 ( .IN1(P2_N4768), .IN2(P2_N5485), .QN(n1301) );
  NAND2X0 U1264 ( .IN1(n7309), .IN2(n9250), .QN(n1300) );
  NAND2X0 U1265 ( .IN1(n1302), .IN2(n1303), .QN(n6237) );
  NAND2X0 U1266 ( .IN1(P2_N4767), .IN2(P2_N5485), .QN(n1303) );
  NAND2X0 U1267 ( .IN1(n7309), .IN2(n9254), .QN(n1302) );
  NAND2X0 U1268 ( .IN1(n1304), .IN2(n1305), .QN(n6238) );
  NAND2X0 U1269 ( .IN1(P2_N4766), .IN2(P2_N5485), .QN(n1305) );
  NAND2X0 U1270 ( .IN1(n7309), .IN2(n9258), .QN(n1304) );
  NAND2X0 U1271 ( .IN1(n1306), .IN2(n1307), .QN(n6239) );
  NAND2X0 U1272 ( .IN1(P2_N4765), .IN2(P2_N5485), .QN(n1307) );
  NAND2X0 U1273 ( .IN1(n7309), .IN2(n9262), .QN(n1306) );
  NAND2X0 U1274 ( .IN1(n1308), .IN2(n1309), .QN(n6240) );
  NAND2X0 U1275 ( .IN1(P2_N4764), .IN2(P2_N5485), .QN(n1309) );
  NAND2X0 U1276 ( .IN1(n7309), .IN2(n10112), .QN(n1308) );
  NAND2X0 U1277 ( .IN1(n1310), .IN2(n1311), .QN(n6241) );
  NAND2X0 U1278 ( .IN1(P2_N4763), .IN2(P2_N5485), .QN(n1311) );
  NAND2X0 U1279 ( .IN1(n7309), .IN2(n6680), .QN(n1310) );
  NAND2X0 U1280 ( .IN1(n1312), .IN2(n1313), .QN(n6242) );
  NAND2X0 U1281 ( .IN1(P2_N4762), .IN2(P2_N5485), .QN(n1313) );
  NAND2X0 U1282 ( .IN1(n7309), .IN2(n6679), .QN(n1312) );
  NAND2X0 U1283 ( .IN1(n1314), .IN2(n1315), .QN(n6243) );
  NAND2X0 U1284 ( .IN1(P2_N4761), .IN2(P2_N5485), .QN(n1315) );
  NAND2X0 U1285 ( .IN1(n7309), .IN2(n6678), .QN(n1314) );
  NAND2X0 U1286 ( .IN1(n1316), .IN2(n1317), .QN(n6244) );
  NAND2X0 U1287 ( .IN1(P2_N4760), .IN2(P2_N5485), .QN(n1317) );
  NAND2X0 U1288 ( .IN1(n7309), .IN2(n6677), .QN(n1316) );
  NAND2X0 U1289 ( .IN1(n1318), .IN2(n1319), .QN(n6245) );
  NAND2X0 U1290 ( .IN1(P2_N4759), .IN2(P2_N5485), .QN(n1319) );
  NAND2X0 U1291 ( .IN1(n7309), .IN2(n6676), .QN(n1318) );
  NAND2X0 U1292 ( .IN1(n1320), .IN2(n1321), .QN(n6246) );
  NAND2X0 U1293 ( .IN1(P2_N4758), .IN2(P2_N5485), .QN(n1321) );
  NAND2X0 U1294 ( .IN1(n7309), .IN2(n6675), .QN(n1320) );
  NAND2X0 U1295 ( .IN1(n1322), .IN2(n1323), .QN(n6247) );
  NAND2X0 U1296 ( .IN1(P2_N4757), .IN2(P2_N5485), .QN(n1323) );
  NAND2X0 U1297 ( .IN1(n7309), .IN2(n6674), .QN(n1322) );
  NAND2X0 U1298 ( .IN1(n1324), .IN2(n1325), .QN(n6248) );
  NAND2X0 U1299 ( .IN1(P2_N4756), .IN2(P2_N5485), .QN(n1325) );
  NAND2X0 U1300 ( .IN1(n7309), .IN2(n6673), .QN(n1324) );
  NAND2X0 U1301 ( .IN1(n1326), .IN2(n1327), .QN(n6249) );
  NAND2X0 U1302 ( .IN1(P2_N4755), .IN2(P2_N5485), .QN(n1327) );
  NAND2X0 U1303 ( .IN1(n7309), .IN2(n6672), .QN(n1326) );
  NAND2X0 U1304 ( .IN1(n1328), .IN2(n1329), .QN(n6250) );
  NAND2X0 U1305 ( .IN1(P2_N4754), .IN2(P2_N5485), .QN(n1329) );
  NAND2X0 U1306 ( .IN1(n7309), .IN2(n6671), .QN(n1328) );
  NAND2X0 U1307 ( .IN1(n1330), .IN2(n1331), .QN(n6251) );
  NAND2X0 U1308 ( .IN1(P2_N4753), .IN2(P2_N5485), .QN(n1331) );
  NAND2X0 U1309 ( .IN1(n7309), .IN2(n10250), .QN(n1330) );
  NAND2X0 U1310 ( .IN1(n1332), .IN2(n1333), .QN(n6252) );
  NAND2X0 U1311 ( .IN1(P2_N4752), .IN2(P2_N5485), .QN(n1333) );
  NAND2X0 U1312 ( .IN1(n7309), .IN2(n6670), .QN(n1332) );
  NAND2X0 U1313 ( .IN1(n1334), .IN2(n1335), .QN(n6253) );
  NAND2X0 U1314 ( .IN1(P2_N4751), .IN2(P2_N5485), .QN(n1335) );
  NAND2X0 U1315 ( .IN1(n7309), .IN2(n6669), .QN(n1334) );
  NAND2X0 U1316 ( .IN1(n1336), .IN2(n1337), .QN(n6254) );
  NAND2X0 U1317 ( .IN1(P2_N4750), .IN2(P2_N5485), .QN(n1337) );
  NAND2X0 U1318 ( .IN1(n7309), .IN2(n6668), .QN(n1336) );
  NAND2X0 U1319 ( .IN1(n1338), .IN2(n1339), .QN(n6255) );
  NAND2X0 U1320 ( .IN1(P2_N4749), .IN2(P2_N5485), .QN(n1339) );
  NAND2X0 U1321 ( .IN1(n7309), .IN2(n6667), .QN(n1338) );
  NAND2X0 U1322 ( .IN1(n1340), .IN2(n1341), .QN(n6256) );
  NAND2X0 U1323 ( .IN1(P2_N4748), .IN2(P2_N5485), .QN(n1341) );
  NAND2X0 U1324 ( .IN1(n7309), .IN2(n6666), .QN(n1340) );
  NAND2X0 U1325 ( .IN1(n1342), .IN2(n1343), .QN(n6257) );
  NAND2X0 U1326 ( .IN1(P2_N4747), .IN2(P2_N5485), .QN(n1343) );
  NAND2X0 U1327 ( .IN1(n7309), .IN2(n6665), .QN(n1342) );
  NAND2X0 U1328 ( .IN1(n1344), .IN2(n1345), .QN(n6258) );
  NAND2X0 U1329 ( .IN1(P2_N4746), .IN2(P2_N5485), .QN(n1345) );
  NAND2X0 U1330 ( .IN1(n7309), .IN2(n6664), .QN(n1344) );
  NAND2X0 U1331 ( .IN1(n1346), .IN2(n1347), .QN(n6259) );
  NAND2X0 U1332 ( .IN1(P2_N4745), .IN2(P2_N5485), .QN(n1347) );
  NAND2X0 U1333 ( .IN1(n7309), .IN2(n9838), .QN(n1346) );
  NAND2X0 U1335 ( .IN1(n1348), .IN2(n1349), .QN(n6260) );
  NAND2X0 U1336 ( .IN1(P2_N4774), .IN2(P2_N5484), .QN(n1349) );
  NAND2X0 U1337 ( .IN1(n7291), .IN2(n9102), .QN(n1348) );
  NAND2X0 U1338 ( .IN1(n1350), .IN2(n1351), .QN(n6261) );
  NAND2X0 U1339 ( .IN1(P2_N4773), .IN2(P2_N5484), .QN(n1351) );
  NAND2X0 U1340 ( .IN1(n7291), .IN2(n9106), .QN(n1350) );
  NAND2X0 U1341 ( .IN1(n1352), .IN2(n1353), .QN(n6262) );
  NAND2X0 U1342 ( .IN1(P2_N4772), .IN2(P2_N5484), .QN(n1353) );
  NAND2X0 U1343 ( .IN1(n7291), .IN2(n9110), .QN(n1352) );
  NAND2X0 U1344 ( .IN1(n1354), .IN2(n1355), .QN(n6263) );
  NAND2X0 U1345 ( .IN1(P2_N4771), .IN2(P2_N5484), .QN(n1355) );
  NAND2X0 U1346 ( .IN1(n7291), .IN2(n9114), .QN(n1354) );
  NAND2X0 U1347 ( .IN1(n1356), .IN2(n1357), .QN(n6264) );
  NAND2X0 U1348 ( .IN1(P2_N4770), .IN2(P2_N5484), .QN(n1357) );
  NAND2X0 U1349 ( .IN1(n7291), .IN2(n9118), .QN(n1356) );
  NAND2X0 U1350 ( .IN1(n1358), .IN2(n1359), .QN(n6265) );
  NAND2X0 U1351 ( .IN1(P2_N4769), .IN2(P2_N5484), .QN(n1359) );
  NAND2X0 U1352 ( .IN1(n7291), .IN2(n9122), .QN(n1358) );
  NAND2X0 U1353 ( .IN1(n1360), .IN2(n1361), .QN(n6266) );
  NAND2X0 U1354 ( .IN1(P2_N4768), .IN2(P2_N5484), .QN(n1361) );
  NAND2X0 U1169 ( .IN1(P2_N4802), .IN2(P2_N5486), .QN(n1239) );
  NAND2X0 U1170 ( .IN1(n7303), .IN2(n9286), .QN(n1238) );
  NAND2X0 U1171 ( .IN1(n1240), .IN2(n1241), .QN(n6206) );
  NAND2X0 U1172 ( .IN1(P2_N4801), .IN2(P2_N5486), .QN(n1241) );
  NAND2X0 U1173 ( .IN1(n7303), .IN2(n9290), .QN(n1240) );
  NAND2X0 U1174 ( .IN1(n1242), .IN2(n1243), .QN(n6207) );
  NAND2X0 U1175 ( .IN1(P2_N4800), .IN2(P2_N5486), .QN(n1243) );
  NAND2X0 U1176 ( .IN1(n7303), .IN2(n9294), .QN(n1242) );
  NAND2X0 U1177 ( .IN1(n1244), .IN2(n1245), .QN(n6208) );
  NAND2X0 U1178 ( .IN1(P2_N4799), .IN2(P2_N5486), .QN(n1245) );
  NAND2X0 U1179 ( .IN1(n7303), .IN2(n9298), .QN(n1244) );
  NAND2X0 U1180 ( .IN1(n1246), .IN2(n1247), .QN(n6209) );
  NAND2X0 U1181 ( .IN1(P2_N4798), .IN2(P2_N5486), .QN(n1247) );
  NAND2X0 U1182 ( .IN1(n7303), .IN2(n9302), .QN(n1246) );
  NAND2X0 U1183 ( .IN1(n1248), .IN2(n1249), .QN(n6210) );
  NAND2X0 U1184 ( .IN1(P2_N4797), .IN2(P2_N5486), .QN(n1249) );
  NAND2X0 U1185 ( .IN1(n7303), .IN2(n10117), .QN(n1248) );
  NAND2X0 U1186 ( .IN1(n1250), .IN2(n1251), .QN(n6211) );
  NAND2X0 U1187 ( .IN1(P2_N4796), .IN2(P2_N5486), .QN(n1251) );
  NAND2X0 U1188 ( .IN1(n7303), .IN2(n6663), .QN(n1250) );
  NAND2X0 U1189 ( .IN1(n1252), .IN2(n1253), .QN(n6212) );
  NAND2X0 U1190 ( .IN1(P2_N4795), .IN2(P2_N5486), .QN(n1253) );
  NAND2X0 U1191 ( .IN1(n7303), .IN2(n6662), .QN(n1252) );
  NAND2X0 U1192 ( .IN1(n1254), .IN2(n1255), .QN(n6213) );
  NAND2X0 U1193 ( .IN1(P2_N4794), .IN2(P2_N5486), .QN(n1255) );
  NAND2X0 U1194 ( .IN1(n7303), .IN2(n6661), .QN(n1254) );
  NAND2X0 U1195 ( .IN1(n1256), .IN2(n1257), .QN(n6214) );
  NAND2X0 U1196 ( .IN1(P2_N4793), .IN2(P2_N5486), .QN(n1257) );
  NAND2X0 U1197 ( .IN1(n7303), .IN2(n6660), .QN(n1256) );
  NAND2X0 U1198 ( .IN1(n1258), .IN2(n1259), .QN(n6215) );
  NAND2X0 U1199 ( .IN1(P2_N4792), .IN2(P2_N5486), .QN(n1259) );
  NAND2X0 U1200 ( .IN1(n7303), .IN2(n6659), .QN(n1258) );
  NAND2X0 U1201 ( .IN1(n1260), .IN2(n1261), .QN(n6216) );
  NAND2X0 U1202 ( .IN1(P2_N4791), .IN2(P2_N5486), .QN(n1261) );
  NAND2X0 U1203 ( .IN1(n7303), .IN2(n6658), .QN(n1260) );
  NAND2X0 U1204 ( .IN1(n1262), .IN2(n1263), .QN(n6217) );
  NAND2X0 U1205 ( .IN1(P2_N4790), .IN2(P2_N5486), .QN(n1263) );
  NAND2X0 U1206 ( .IN1(n7303), .IN2(n6657), .QN(n1262) );
  NAND2X0 U1207 ( .IN1(n1264), .IN2(n1265), .QN(n6218) );
  NAND2X0 U1208 ( .IN1(P2_N4789), .IN2(P2_N5486), .QN(n1265) );
  NAND2X0 U1209 ( .IN1(n7303), .IN2(n6656), .QN(n1264) );
  NAND2X0 U1210 ( .IN1(n1266), .IN2(n1267), .QN(n6219) );
  NAND2X0 U1211 ( .IN1(P2_N4788), .IN2(P2_N5486), .QN(n1267) );
  NAND2X0 U1212 ( .IN1(n7303), .IN2(n6655), .QN(n1266) );
  NAND2X0 U1213 ( .IN1(n1268), .IN2(n1269), .QN(n6220) );
  NAND2X0 U1214 ( .IN1(P2_N4787), .IN2(P2_N5486), .QN(n1269) );
  NAND2X0 U1215 ( .IN1(n7303), .IN2(n6654), .QN(n1268) );
  NAND2X0 U1216 ( .IN1(n1270), .IN2(n1271), .QN(n6221) );
  NAND2X0 U1217 ( .IN1(P2_N4786), .IN2(P2_N5486), .QN(n1271) );
  NAND2X0 U1218 ( .IN1(n7303), .IN2(n6653), .QN(n1270) );
  NAND2X0 U1219 ( .IN1(n1272), .IN2(n1273), .QN(n6222) );
  NAND2X0 U1220 ( .IN1(P2_N4785), .IN2(P2_N5486), .QN(n1273) );
  NAND2X0 U1221 ( .IN1(n7303), .IN2(n6652), .QN(n1272) );
  NAND2X0 U1222 ( .IN1(n1274), .IN2(n1275), .QN(n6223) );
  NAND2X0 U1223 ( .IN1(P2_N4784), .IN2(P2_N5486), .QN(n1275) );
  NAND2X0 U1224 ( .IN1(n7303), .IN2(n6651), .QN(n1274) );
  NAND2X0 U1225 ( .IN1(n1276), .IN2(n1277), .QN(n6224) );
  NAND2X0 U1226 ( .IN1(P2_N4783), .IN2(P2_N5486), .QN(n1277) );
  NAND2X0 U1227 ( .IN1(n7303), .IN2(n6650), .QN(n1276) );
  NAND2X0 U1228 ( .IN1(n1278), .IN2(n1279), .QN(n6225) );
  NAND2X0 U1229 ( .IN1(P2_N4782), .IN2(P2_N5486), .QN(n1279) );
  NAND2X0 U1230 ( .IN1(n7303), .IN2(n6649), .QN(n1278) );
  NAND2X0 U1231 ( .IN1(n1280), .IN2(n1281), .QN(n6226) );
  NAND2X0 U1232 ( .IN1(P2_N4781), .IN2(P2_N5486), .QN(n1281) );
  NAND2X0 U1233 ( .IN1(n7303), .IN2(n6648), .QN(n1280) );
  NAND2X0 U1234 ( .IN1(n1282), .IN2(n1283), .QN(n6227) );
  NAND2X0 U1235 ( .IN1(P2_N4780), .IN2(P2_N5486), .QN(n1283) );
  NAND2X0 U1236 ( .IN1(n7303), .IN2(n6721), .QN(n1282) );
  NAND2X0 U1237 ( .IN1(n1284), .IN2(n1285), .QN(n6228) );
  NAND2X0 U1238 ( .IN1(P2_N4779), .IN2(P2_N5486), .QN(n1285) );
  NAND2X0 U1239 ( .IN1(n7303), .IN2(n6720), .QN(n1284) );
  NAND2X0 U1240 ( .IN1(n1286), .IN2(n1287), .QN(n6229) );
  NAND2X0 U1241 ( .IN1(P2_N4778), .IN2(P2_N5486), .QN(n1287) );
  NAND2X0 U1242 ( .IN1(n7303), .IN2(n9843), .QN(n1286) );
  NAND2X0 U1244 ( .IN1(n1288), .IN2(n1289), .QN(n6230) );
  NAND2X0 U1245 ( .IN1(P2_N4774), .IN2(P2_N5485), .QN(n1289) );
  NAND2X0 U1246 ( .IN1(n7309), .IN2(n9226), .QN(n1288) );
  NAND2X0 U1247 ( .IN1(n1290), .IN2(n1291), .QN(n6231) );
  NAND2X0 U1248 ( .IN1(P2_N4773), .IN2(P2_N5485), .QN(n1291) );
  NAND2X0 U1249 ( .IN1(n7309), .IN2(n9230), .QN(n1290) );
  NAND2X0 U1250 ( .IN1(n1292), .IN2(n1293), .QN(n6232) );
  NAND2X0 U1251 ( .IN1(P2_N4772), .IN2(P2_N5485), .QN(n1293) );
  NAND2X0 U1252 ( .IN1(n7309), .IN2(n9234), .QN(n1292) );
  NAND2X0 U1253 ( .IN1(n1294), .IN2(n1295), .QN(n6233) );
  NAND2X0 U1254 ( .IN1(P2_N4771), .IN2(P2_N5485), .QN(n1295) );
  NAND2X0 U1255 ( .IN1(n7309), .IN2(n9238), .QN(n1294) );
  NAND2X0 U1256 ( .IN1(n1296), .IN2(n1297), .QN(n6234) );
  NAND2X0 U1257 ( .IN1(P2_N4770), .IN2(P2_N5485), .QN(n1297) );
  NAND2X0 U1258 ( .IN1(n7309), .IN2(n9242), .QN(n1296) );
  NAND2X0 U1259 ( .IN1(n1298), .IN2(n1299), .QN(n6235) );
  NAND2X0 U1260 ( .IN1(P2_N4769), .IN2(P2_N5485), .QN(n1299) );
  NAND2X0 U1261 ( .IN1(n7309), .IN2(n9246), .QN(n1298) );
  NAND2X0 U1076 ( .IN1(n1176), .IN2(n1177), .QN(n6175) );
  NAND2X0 U1077 ( .IN1(P2_N5072), .IN2(P2_N5476), .QN(n1177) );
  NAND2X0 U1078 ( .IN1(n7270), .IN2(n9337), .QN(n1176) );
  NAND2X0 U1079 ( .IN1(n1178), .IN2(n1179), .QN(n6176) );
  NAND2X0 U1080 ( .IN1(n7270), .IN2(n9389), .QN(n1179) );
  NAND2X0 U1082 ( .IN1(P2_N5476), .IN2(n7035), .QN(n1178) );
  NAND2X0 U1083 ( .IN1(n1180), .IN2(n1181), .QN(n6177) );
  NAND2X0 U1084 ( .IN1(n6729), .IN2(n10133), .QN(n1181) );
  NAND2X0 U1085 ( .IN1(P2_N5473), .IN2(P2_N5470), .QN(n1180) );
  NAND2X0 U1086 ( .IN1(n1183), .IN2(n1184), .QN(n6178) );
  NAND2X0 U1087 ( .IN1(n7285), .IN2(n18209), .QN(n1184) );
  NAND2X0 U1088 ( .IN1(P2_N5439), .IN2(P2_N5419), .QN(n1183) );
  NAND2X0 U1089 ( .IN1(n1186), .IN2(n1187), .QN(n6179) );
  NAND2X0 U1090 ( .IN1(n7285), .IN2(n9417), .QN(n1187) );
  NAND2X0 U1091 ( .IN1(P2_N5438), .IN2(P2_N5419), .QN(n1186) );
  NAND2X0 U1092 ( .IN1(n1188), .IN2(n1189), .QN(n6180) );
  NAND2X0 U1093 ( .IN1(n7285), .IN2(n9421), .QN(n1189) );
  NAND2X0 U1094 ( .IN1(P2_N5437), .IN2(P2_N5419), .QN(n1188) );
  NAND2X0 U1095 ( .IN1(n1190), .IN2(n1191), .QN(n6181) );
  NAND2X0 U1096 ( .IN1(n7285), .IN2(n9425), .QN(n1191) );
  NAND2X0 U1097 ( .IN1(P2_N5436), .IN2(P2_N5419), .QN(n1190) );
  NAND2X0 U1098 ( .IN1(n1192), .IN2(n1193), .QN(n6182) );
  NAND2X0 U1099 ( .IN1(n7285), .IN2(n9429), .QN(n1193) );
  NAND2X0 U1100 ( .IN1(P2_N5435), .IN2(P2_N5419), .QN(n1192) );
  NAND2X0 U1101 ( .IN1(n1194), .IN2(n1195), .QN(n6183) );
  NAND2X0 U1102 ( .IN1(n7285), .IN2(n9433), .QN(n1195) );
  NAND2X0 U1103 ( .IN1(P2_N5434), .IN2(P2_N5419), .QN(n1194) );
  NAND2X0 U1104 ( .IN1(n1196), .IN2(n1197), .QN(n6184) );
  NAND2X0 U1105 ( .IN1(n7285), .IN2(n9437), .QN(n1197) );
  NAND2X0 U1106 ( .IN1(P2_N5433), .IN2(P2_N5419), .QN(n1196) );
  NAND2X0 U1107 ( .IN1(n1198), .IN2(n1199), .QN(n6185) );
  NAND2X0 U1108 ( .IN1(n7285), .IN2(n9441), .QN(n1199) );
  NAND2X0 U1109 ( .IN1(P2_N5432), .IN2(P2_N5419), .QN(n1198) );
  NAND2X0 U1110 ( .IN1(n1200), .IN2(n1201), .QN(n6186) );
  NAND2X0 U1111 ( .IN1(n7285), .IN2(n9445), .QN(n1201) );
  NAND2X0 U1112 ( .IN1(P2_N5431), .IN2(P2_N5419), .QN(n1200) );
  NAND2X0 U1113 ( .IN1(n1202), .IN2(n1203), .QN(n6187) );
  NAND2X0 U1114 ( .IN1(n7285), .IN2(n9449), .QN(n1203) );
  NAND2X0 U1115 ( .IN1(P2_N5430), .IN2(P2_N5419), .QN(n1202) );
  NAND2X0 U1116 ( .IN1(n1204), .IN2(n1205), .QN(n6188) );
  NAND2X0 U1117 ( .IN1(n7285), .IN2(n9453), .QN(n1205) );
  NAND2X0 U1118 ( .IN1(P2_N5429), .IN2(P2_N5419), .QN(n1204) );
  NAND2X0 U1119 ( .IN1(n1206), .IN2(n1207), .QN(n6189) );
  NAND2X0 U1120 ( .IN1(n7285), .IN2(n9457), .QN(n1207) );
  NAND2X0 U1121 ( .IN1(P2_N5428), .IN2(P2_N5419), .QN(n1206) );
  NAND2X0 U1122 ( .IN1(n1208), .IN2(n1209), .QN(n6190) );
  NAND2X0 U1123 ( .IN1(n7285), .IN2(n9461), .QN(n1209) );
  NAND2X0 U1124 ( .IN1(P2_N5427), .IN2(P2_N5419), .QN(n1208) );
  NAND2X0 U1125 ( .IN1(n1210), .IN2(n1211), .QN(n6191) );
  NAND2X0 U1126 ( .IN1(n7285), .IN2(n9465), .QN(n1211) );
  NAND2X0 U1127 ( .IN1(P2_N5426), .IN2(P2_N5419), .QN(n1210) );
  NAND2X0 U1128 ( .IN1(n1212), .IN2(n1213), .QN(n6192) );
  NAND2X0 U1129 ( .IN1(n7285), .IN2(n9469), .QN(n1213) );
  NAND2X0 U1130 ( .IN1(P2_N5425), .IN2(P2_N5419), .QN(n1212) );
  NAND2X0 U1131 ( .IN1(n1214), .IN2(n1215), .QN(n6193) );
  NAND2X0 U1132 ( .IN1(n7285), .IN2(n9473), .QN(n1215) );
  NAND2X0 U1133 ( .IN1(P2_N5424), .IN2(P2_N5419), .QN(n1214) );
  NAND2X0 U1134 ( .IN1(n1216), .IN2(n1217), .QN(n6194) );
  NAND2X0 U1135 ( .IN1(n7285), .IN2(n9477), .QN(n1217) );
  NAND2X0 U1136 ( .IN1(P2_N5423), .IN2(P2_N5419), .QN(n1216) );
  NAND2X0 U1137 ( .IN1(n1218), .IN2(n1219), .QN(n6195) );
  NAND2X0 U1138 ( .IN1(n7285), .IN2(n9481), .QN(n1219) );
  NAND2X0 U1139 ( .IN1(P2_N5422), .IN2(P2_N5419), .QN(n1218) );
  NAND2X0 U1140 ( .IN1(n1220), .IN2(n1221), .QN(n6196) );
  NAND2X0 U1141 ( .IN1(n7285), .IN2(n9485), .QN(n1221) );
  NAND2X0 U1142 ( .IN1(P2_N5421), .IN2(P2_N5419), .QN(n1220) );
  NAND2X0 U1143 ( .IN1(n1222), .IN2(n1223), .QN(n6197) );
  NAND2X0 U1144 ( .IN1(n7285), .IN2(n9489), .QN(n1223) );
  NAND2X0 U1146 ( .IN1(P2_N5420), .IN2(P2_N5419), .QN(n1222) );
  NAND2X0 U1147 ( .IN1(n1224), .IN2(n1225), .QN(n6198) );
  NAND2X0 U1148 ( .IN1(n6729), .IN2(n10141), .QN(n1225) );
  NAND2X0 U1149 ( .IN1(P2_N5472), .IN2(P2_N5470), .QN(n1224) );
  NAND2X0 U1150 ( .IN1(n1226), .IN2(n1227), .QN(n6199) );
  NAND2X0 U1151 ( .IN1(n6729), .IN2(n10369), .QN(n1227) );
  NAND2X0 U1152 ( .IN1(P2_N5471), .IN2(P2_N5470), .QN(n1226) );
  NAND2X0 U1153 ( .IN1(n1228), .IN2(n1229), .QN(n6200) );
  NAND2X0 U1154 ( .IN1(P2_N4807), .IN2(P2_N5486), .QN(n1229) );
  NAND2X0 U1155 ( .IN1(n7303), .IN2(n9266), .QN(n1228) );
  NAND2X0 U1156 ( .IN1(n1230), .IN2(n1231), .QN(n6201) );
  NAND2X0 U1157 ( .IN1(P2_N4806), .IN2(P2_N5486), .QN(n1231) );
  NAND2X0 U1158 ( .IN1(n7303), .IN2(n9270), .QN(n1230) );
  NAND2X0 U1159 ( .IN1(n1232), .IN2(n1233), .QN(n6202) );
  NAND2X0 U1160 ( .IN1(P2_N4805), .IN2(P2_N5486), .QN(n1233) );
  NAND2X0 U1161 ( .IN1(n7303), .IN2(n9274), .QN(n1232) );
  NAND2X0 U1162 ( .IN1(n1234), .IN2(n1235), .QN(n6203) );
  NAND2X0 U1163 ( .IN1(P2_N4804), .IN2(P2_N5486), .QN(n1235) );
  NAND2X0 U1164 ( .IN1(n7303), .IN2(n9278), .QN(n1234) );
  NAND2X0 U1165 ( .IN1(n1236), .IN2(n1237), .QN(n6204) );
  NAND2X0 U1166 ( .IN1(P2_N4803), .IN2(P2_N5486), .QN(n1237) );
  NAND2X0 U1167 ( .IN1(n7303), .IN2(n9282), .QN(n1236) );
  NAND2X0 U1168 ( .IN1(n1238), .IN2(n1239), .QN(n6205) );
  NAND2X0 U983 ( .IN1(n7270), .IN2(n10099), .QN(n1112) );
  NAND2X0 U984 ( .IN1(n1114), .IN2(n1115), .QN(n6145) );
  NAND2X0 U985 ( .IN1(P2_N5482), .IN2(P2_N531), .QN(n1115) );
  NAND2X0 U986 ( .IN1(n1116), .IN2(n6592), .QN(n1114) );
  NAND2X0 U987 ( .IN1(n1117), .IN2(n1118), .QN(n6146) );
  NAND2X0 U988 ( .IN1(P2_N530), .IN2(P2_N5482), .QN(n1118) );
  NAND2X0 U989 ( .IN1(n1116), .IN2(n6593), .QN(n1117) );
  INVX0 U990 ( .ZN(n1116), .INP(P2_N5482) );
  NAND2X0 U991 ( .IN1(n1119), .IN2(n1120), .QN(n6147) );
  NAND2X0 U992 ( .IN1(n6591), .IN2(n1121), .QN(n1120) );
  INVX0 U993 ( .ZN(n1121), .INP(P2_N5483) );
  NAND2X0 U994 ( .IN1(P2_N5483), .IN2(n7442), .QN(n1119) );
  NAND2X0 U995 ( .IN1(n1122), .IN2(n1123), .QN(n6148) );
  NAND2X0 U996 ( .IN1(P2_N5099), .IN2(P2_N5476), .QN(n1123) );
  NAND2X0 U997 ( .IN1(n7270), .IN2(n10019), .QN(n1122) );
  NAND2X0 U998 ( .IN1(n1124), .IN2(n1125), .QN(n6149) );
  NAND2X0 U999 ( .IN1(n7227), .IN2(P2_N5476), .QN(n1125) );
  NAND2X0 U1000 ( .IN1(n7270), .IN2(n10023), .QN(n1124) );
  NAND2X0 U1001 ( .IN1(n1126), .IN2(n1127), .QN(n6150) );
  NAND2X0 U1002 ( .IN1(n7231), .IN2(P2_N5476), .QN(n1127) );
  NAND2X0 U1003 ( .IN1(n7270), .IN2(n10027), .QN(n1126) );
  NAND2X0 U1004 ( .IN1(n1128), .IN2(n1129), .QN(n6151) );
  NAND2X0 U1005 ( .IN1(P2_N5096), .IN2(P2_N5476), .QN(n1129) );
  NAND2X0 U1006 ( .IN1(n7270), .IN2(n10031), .QN(n1128) );
  NAND2X0 U1007 ( .IN1(n1130), .IN2(n1131), .QN(n6152) );
  NAND2X0 U1008 ( .IN1(n7238), .IN2(P2_N5476), .QN(n1131) );
  NAND2X0 U1009 ( .IN1(n7270), .IN2(n10035), .QN(n1130) );
  NAND2X0 U1010 ( .IN1(n1132), .IN2(n1133), .QN(n6153) );
  NAND2X0 U1011 ( .IN1(P2_N5094), .IN2(P2_N5476), .QN(n1133) );
  NAND2X0 U1012 ( .IN1(n7270), .IN2(n10039), .QN(n1132) );
  NAND2X0 U1013 ( .IN1(n1134), .IN2(n1135), .QN(n6154) );
  NAND2X0 U1014 ( .IN1(P2_N5093), .IN2(P2_N5476), .QN(n1135) );
  NAND2X0 U1015 ( .IN1(n7270), .IN2(n10043), .QN(n1134) );
  NAND2X0 U1016 ( .IN1(n1136), .IN2(n1137), .QN(n6155) );
  NAND2X0 U1017 ( .IN1(P2_N5092), .IN2(P2_N5476), .QN(n1137) );
  NAND2X0 U1018 ( .IN1(n7270), .IN2(n10047), .QN(n1136) );
  NAND2X0 U1019 ( .IN1(n1138), .IN2(n1139), .QN(n6156) );
  NAND2X0 U1020 ( .IN1(n7259), .IN2(P2_N5476), .QN(n1139) );
  NAND2X0 U1021 ( .IN1(n7270), .IN2(n10051), .QN(n1138) );
  NAND2X0 U1022 ( .IN1(n1140), .IN2(n1141), .QN(n6157) );
  NAND2X0 U1023 ( .IN1(n7263), .IN2(P2_N5476), .QN(n1141) );
  NAND2X0 U1024 ( .IN1(n7270), .IN2(n10055), .QN(n1140) );
  NAND2X0 U1025 ( .IN1(n1142), .IN2(n1143), .QN(n6158) );
  NAND2X0 U1026 ( .IN1(P2_N5089), .IN2(P2_N5476), .QN(n1143) );
  NAND2X0 U1027 ( .IN1(n7270), .IN2(n10059), .QN(n1142) );
  NAND2X0 U1028 ( .IN1(n1144), .IN2(n1145), .QN(n6159) );
  NAND2X0 U1029 ( .IN1(P2_N5088), .IN2(P2_N5476), .QN(n1145) );
  NAND2X0 U1030 ( .IN1(n7270), .IN2(n10063), .QN(n1144) );
  NAND2X0 U1031 ( .IN1(n1146), .IN2(n1147), .QN(n6160) );
  NAND2X0 U1032 ( .IN1(n7198), .IN2(P2_N5476), .QN(n1147) );
  NAND2X0 U1033 ( .IN1(n7270), .IN2(n10067), .QN(n1146) );
  NAND2X0 U1034 ( .IN1(n1148), .IN2(n1149), .QN(n6161) );
  NAND2X0 U1035 ( .IN1(n7202), .IN2(P2_N5476), .QN(n1149) );
  NAND2X0 U1036 ( .IN1(n7270), .IN2(n10071), .QN(n1148) );
  NAND2X0 U1037 ( .IN1(n1150), .IN2(n1151), .QN(n6162) );
  NAND2X0 U1038 ( .IN1(n7206), .IN2(P2_N5476), .QN(n1151) );
  NAND2X0 U1039 ( .IN1(n7270), .IN2(n10075), .QN(n1150) );
  NAND2X0 U1040 ( .IN1(n1152), .IN2(n1153), .QN(n6163) );
  NAND2X0 U1041 ( .IN1(n7209), .IN2(P2_N5476), .QN(n1153) );
  NAND2X0 U1042 ( .IN1(n7270), .IN2(n10079), .QN(n1152) );
  NAND2X0 U1043 ( .IN1(n1154), .IN2(n1155), .QN(n6164) );
  NAND2X0 U1044 ( .IN1(P2_N5083), .IN2(P2_N5476), .QN(n1155) );
  NAND2X0 U1045 ( .IN1(n7270), .IN2(n10083), .QN(n1154) );
  NAND2X0 U1046 ( .IN1(n1156), .IN2(n1157), .QN(n6165) );
  NAND2X0 U1047 ( .IN1(n7216), .IN2(P2_N5476), .QN(n1157) );
  NAND2X0 U1048 ( .IN1(n7270), .IN2(n10087), .QN(n1156) );
  NAND2X0 U1049 ( .IN1(n1158), .IN2(n1159), .QN(n6166) );
  NAND2X0 U1050 ( .IN1(n7220), .IN2(P2_N5476), .QN(n1159) );
  NAND2X0 U1051 ( .IN1(n7270), .IN2(n10091), .QN(n1158) );
  NAND2X0 U1052 ( .IN1(n1160), .IN2(n1161), .QN(n6167) );
  NAND2X0 U1053 ( .IN1(P2_N5080), .IN2(P2_N5476), .QN(n1161) );
  NAND2X0 U1054 ( .IN1(n7270), .IN2(n9903), .QN(n1160) );
  NAND2X0 U1055 ( .IN1(n1162), .IN2(n1163), .QN(n6168) );
  NAND2X0 U1056 ( .IN1(n7154), .IN2(P2_N5476), .QN(n1163) );
  NAND2X0 U1057 ( .IN1(n7270), .IN2(n9907), .QN(n1162) );
  NAND2X0 U1058 ( .IN1(n1164), .IN2(n1165), .QN(n6169) );
  NAND2X0 U1059 ( .IN1(n7158), .IN2(P2_N5476), .QN(n1165) );
  NAND2X0 U1060 ( .IN1(n7270), .IN2(n9911), .QN(n1164) );
  NAND2X0 U1061 ( .IN1(n1166), .IN2(n1167), .QN(n6170) );
  NAND2X0 U1062 ( .IN1(n7162), .IN2(P2_N5476), .QN(n1167) );
  NAND2X0 U1063 ( .IN1(n7270), .IN2(n9915), .QN(n1166) );
  NAND2X0 U1064 ( .IN1(n1168), .IN2(n1169), .QN(n6171) );
  NAND2X0 U1065 ( .IN1(n7165), .IN2(P2_N5476), .QN(n1169) );
  NAND2X0 U1066 ( .IN1(n7270), .IN2(n9919), .QN(n1168) );
  NAND2X0 U1067 ( .IN1(n1170), .IN2(n1171), .QN(n6172) );
  NAND2X0 U1068 ( .IN1(P2_N5075), .IN2(P2_N5476), .QN(n1171) );
  NAND2X0 U1069 ( .IN1(n7270), .IN2(n9923), .QN(n1170) );
  NAND2X0 U1070 ( .IN1(n1172), .IN2(n1173), .QN(n6173) );
  NAND2X0 U1071 ( .IN1(n7177), .IN2(P2_N5476), .QN(n1173) );
  NAND2X0 U1072 ( .IN1(n7270), .IN2(n9927), .QN(n1172) );
  NAND2X0 U1073 ( .IN1(n1174), .IN2(n1175), .QN(n6174) );
  NAND2X0 U1074 ( .IN1(n7181), .IN2(P2_N5476), .QN(n1175) );
  NAND2X0 U1075 ( .IN1(n7270), .IN2(n9931), .QN(n1174) );
  NAND2X0 U890 ( .IN1(n1051), .IN2(n1052), .QN(n6114) );
  NAND2X0 U891 ( .IN1(P1_N5547), .IN2(P1_N5548), .QN(n1052) );
  NAND2X0 U892 ( .IN1(n6725), .IN2(n10187), .QN(n1051) );
  NAND2X0 U893 ( .IN1(n1053), .IN2(n1054), .QN(n6115) );
  NAND2X0 U894 ( .IN1(P1_N5546), .IN2(P1_N5548), .QN(n1054) );
  NAND2X0 U895 ( .IN1(n6725), .IN2(n10381), .QN(n1053) );
  NAND2X0 U896 ( .IN1(n1055), .IN2(n1056), .QN(n6116) );
  NAND2X0 U897 ( .IN1(P1_N5545), .IN2(P1_N5548), .QN(n1056) );
  NAND2X0 U898 ( .IN1(n6725), .IN2(n10195), .QN(n1055) );
  NAND2X0 U899 ( .IN1(n1057), .IN2(n1058), .QN(n6117) );
  NAND2X0 U900 ( .IN1(P1_N5544), .IN2(P1_N5548), .QN(n1058) );
  NAND2X0 U901 ( .IN1(n6725), .IN2(n6637), .QN(n1057) );
  NAND2X0 U902 ( .IN1(n1059), .IN2(n1060), .QN(n6118) );
  NAND2X0 U903 ( .IN1(P1_N5543), .IN2(P1_N5548), .QN(n1060) );
  NAND2X0 U904 ( .IN1(n6725), .IN2(n6638), .QN(n1059) );
  NAND2X0 U905 ( .IN1(n1061), .IN2(n1062), .QN(n6119) );
  NAND2X0 U906 ( .IN1(P1_N5542), .IN2(P1_N5548), .QN(n1062) );
  NAND2X0 U907 ( .IN1(n6725), .IN2(n6639), .QN(n1061) );
  NAND2X0 U908 ( .IN1(n1063), .IN2(n1064), .QN(n6120) );
  NAND2X0 U909 ( .IN1(P1_N5541), .IN2(P1_N5548), .QN(n1064) );
  NAND2X0 U910 ( .IN1(n6725), .IN2(n6640), .QN(n1063) );
  NAND2X0 U911 ( .IN1(n1065), .IN2(n1066), .QN(n6121) );
  NAND2X0 U912 ( .IN1(P1_N5540), .IN2(P1_N5548), .QN(n1066) );
  NAND2X0 U913 ( .IN1(n6725), .IN2(n6641), .QN(n1065) );
  NAND2X0 U914 ( .IN1(n1067), .IN2(n1068), .QN(n6122) );
  NAND2X0 U915 ( .IN1(P1_N5539), .IN2(P1_N5548), .QN(n1068) );
  NAND2X0 U916 ( .IN1(n6725), .IN2(n6642), .QN(n1067) );
  NAND2X0 U917 ( .IN1(n1069), .IN2(n1070), .QN(n6123) );
  NAND2X0 U918 ( .IN1(P1_N5538), .IN2(P1_N5548), .QN(n1070) );
  NAND2X0 U919 ( .IN1(n6725), .IN2(n6643), .QN(n1069) );
  NAND2X0 U920 ( .IN1(n1071), .IN2(n1072), .QN(n6124) );
  NAND2X0 U921 ( .IN1(P1_N5537), .IN2(P1_N5548), .QN(n1072) );
  NAND2X0 U922 ( .IN1(n6725), .IN2(n6644), .QN(n1071) );
  NAND2X0 U923 ( .IN1(n1073), .IN2(n1074), .QN(n6125) );
  NAND2X0 U924 ( .IN1(P1_N5536), .IN2(P1_N5548), .QN(n1074) );
  NAND2X0 U925 ( .IN1(n6725), .IN2(n6645), .QN(n1073) );
  NAND2X0 U926 ( .IN1(n1075), .IN2(n1076), .QN(n6126) );
  NAND2X0 U927 ( .IN1(P1_N5535), .IN2(P1_N5548), .QN(n1076) );
  NAND2X0 U928 ( .IN1(n6725), .IN2(n6646), .QN(n1075) );
  NAND2X0 U929 ( .IN1(n1077), .IN2(n1078), .QN(n6127) );
  NAND2X0 U930 ( .IN1(P1_N5534), .IN2(P1_N5548), .QN(n1078) );
  NAND2X0 U931 ( .IN1(n6725), .IN2(n6647), .QN(n1077) );
  NAND2X0 U932 ( .IN1(n1079), .IN2(n1080), .QN(n6128) );
  NAND2X0 U933 ( .IN1(P1_N5532), .IN2(P1_N5548), .QN(n1080) );
  NAND2X0 U934 ( .IN1(n6725), .IN2(n6636), .QN(n1079) );
  NAND2X0 U935 ( .IN1(n1081), .IN2(n1082), .QN(n6129) );
  NAND2X0 U936 ( .IN1(P1_N5531), .IN2(P1_N5548), .QN(n1082) );
  NAND2X0 U937 ( .IN1(n6725), .IN2(n6635), .QN(n1081) );
  NAND2X0 U938 ( .IN1(n1083), .IN2(n1084), .QN(n6130) );
  NAND2X0 U939 ( .IN1(P1_N5530), .IN2(P1_N5548), .QN(n1084) );
  NAND2X0 U940 ( .IN1(n6725), .IN2(n6634), .QN(n1083) );
  NAND2X0 U941 ( .IN1(n1085), .IN2(n1086), .QN(n6131) );
  NAND2X0 U942 ( .IN1(P1_N5529), .IN2(P1_N5548), .QN(n1086) );
  NAND2X0 U943 ( .IN1(n6725), .IN2(n6633), .QN(n1085) );
  NAND2X0 U944 ( .IN1(n1087), .IN2(n1088), .QN(n6132) );
  NAND2X0 U945 ( .IN1(P1_N5528), .IN2(P1_N5548), .QN(n1088) );
  NAND2X0 U946 ( .IN1(n6725), .IN2(n6632), .QN(n1087) );
  NAND2X0 U947 ( .IN1(n1089), .IN2(n1090), .QN(n6133) );
  NAND2X0 U948 ( .IN1(P1_N5527), .IN2(P1_N5548), .QN(n1090) );
  NAND2X0 U949 ( .IN1(n6725), .IN2(n6631), .QN(n1089) );
  NAND2X0 U950 ( .IN1(n1091), .IN2(n1092), .QN(n6134) );
  NAND2X0 U951 ( .IN1(P1_N5526), .IN2(P1_N5548), .QN(n1092) );
  NAND2X0 U952 ( .IN1(n6725), .IN2(n6630), .QN(n1091) );
  NAND2X0 U953 ( .IN1(n1093), .IN2(n1094), .QN(n6135) );
  NAND2X0 U954 ( .IN1(P1_N5525), .IN2(P1_N5548), .QN(n1094) );
  NAND2X0 U955 ( .IN1(n6725), .IN2(n6629), .QN(n1093) );
  NAND2X0 U956 ( .IN1(n1095), .IN2(n1096), .QN(n6136) );
  NAND2X0 U957 ( .IN1(P1_N5524), .IN2(P1_N5548), .QN(n1096) );
  NAND2X0 U958 ( .IN1(n6725), .IN2(n6628), .QN(n1095) );
  NAND2X0 U959 ( .IN1(n1097), .IN2(n1098), .QN(n6137) );
  NAND2X0 U960 ( .IN1(P1_N5523), .IN2(P1_N5548), .QN(n1098) );
  NAND2X0 U961 ( .IN1(n6725), .IN2(n6627), .QN(n1097) );
  NAND2X0 U962 ( .IN1(n1099), .IN2(n1100), .QN(n6138) );
  NAND2X0 U963 ( .IN1(P1_N5522), .IN2(P1_N5548), .QN(n1100) );
  NAND2X0 U964 ( .IN1(n6725), .IN2(n6626), .QN(n1099) );
  NAND2X0 U965 ( .IN1(n1101), .IN2(n1102), .QN(n6139) );
  NAND2X0 U966 ( .IN1(P1_N5521), .IN2(P1_N5548), .QN(n1102) );
  NAND2X0 U967 ( .IN1(n6725), .IN2(n6625), .QN(n1101) );
  NAND2X0 U968 ( .IN1(n1103), .IN2(n1104), .QN(n6140) );
  NAND2X0 U969 ( .IN1(P1_N5520), .IN2(P1_N5548), .QN(n1104) );
  NAND2X0 U970 ( .IN1(n6725), .IN2(n6624), .QN(n1103) );
  NAND2X0 U971 ( .IN1(n1105), .IN2(n1106), .QN(n6141) );
  NAND2X0 U972 ( .IN1(n6725), .IN2(n6718), .QN(n1106) );
  NAND2X0 U974 ( .IN1(P1_N5553), .IN2(P1_N5548), .QN(n1105) );
  NAND2X0 U975 ( .IN1(n1107), .IN2(n1108), .QN(n6142) );
  NAND2X0 U976 ( .IN1(n7270), .IN2(n9341), .QN(n1108) );
  NAND2X0 U977 ( .IN1(P2_N5476), .IN2(n7147), .QN(n1107) );
  NAND2X0 U978 ( .IN1(n1110), .IN2(n1111), .QN(n6143) );
  NAND2X0 U979 ( .IN1(P2_N497), .IN2(P2_N5476), .QN(n1111) );
  NAND2X0 U980 ( .IN1(n7270), .IN2(n10107), .QN(n1110) );
  NAND2X0 U981 ( .IN1(n1112), .IN2(n1113), .QN(n6144) );
  NAND2X0 U982 ( .IN1(P2_N5100), .IN2(P2_N5476), .QN(n1113) );
  NAND2X0 U797 ( .IN1(P1_N4899), .IN2(P1_N5562), .QN(n989) );
  NAND2X0 U798 ( .IN1(n7287), .IN2(n8902), .QN(n988) );
  NAND2X0 U799 ( .IN1(n990), .IN2(n991), .QN(n6084) );
  NAND2X0 U800 ( .IN1(P1_N4898), .IN2(P1_N5562), .QN(n991) );
  NAND2X0 U801 ( .IN1(n7287), .IN2(n8906), .QN(n990) );
  NAND2X0 U802 ( .IN1(n992), .IN2(n993), .QN(n6085) );
  NAND2X0 U803 ( .IN1(P1_N4897), .IN2(P1_N5562), .QN(n993) );
  NAND2X0 U804 ( .IN1(n7287), .IN2(n8910), .QN(n992) );
  NAND2X0 U805 ( .IN1(n994), .IN2(n995), .QN(n6086) );
  NAND2X0 U806 ( .IN1(P1_N4896), .IN2(P1_N5562), .QN(n995) );
  NAND2X0 U807 ( .IN1(n7287), .IN2(n8914), .QN(n994) );
  NAND2X0 U808 ( .IN1(n996), .IN2(n997), .QN(n6087) );
  NAND2X0 U809 ( .IN1(P1_N4895), .IN2(P1_N5562), .QN(n997) );
  NAND2X0 U810 ( .IN1(n7287), .IN2(n8918), .QN(n996) );
  NAND2X0 U811 ( .IN1(n998), .IN2(n999), .QN(n6088) );
  NAND2X0 U812 ( .IN1(P1_N4894), .IN2(P1_N5562), .QN(n999) );
  NAND2X0 U813 ( .IN1(n7287), .IN2(n8922), .QN(n998) );
  NAND2X0 U814 ( .IN1(n1000), .IN2(n1001), .QN(n6089) );
  NAND2X0 U815 ( .IN1(P1_N4893), .IN2(P1_N5562), .QN(n1001) );
  NAND2X0 U816 ( .IN1(n7287), .IN2(n8926), .QN(n1000) );
  NAND2X0 U817 ( .IN1(n1002), .IN2(n1003), .QN(n6090) );
  NAND2X0 U818 ( .IN1(P1_N4892), .IN2(P1_N5562), .QN(n1003) );
  NAND2X0 U819 ( .IN1(n7287), .IN2(n8930), .QN(n1002) );
  NAND2X0 U820 ( .IN1(n1004), .IN2(n1005), .QN(n6091) );
  NAND2X0 U821 ( .IN1(P1_N4891), .IN2(P1_N5562), .QN(n1005) );
  NAND2X0 U822 ( .IN1(n7287), .IN2(n8934), .QN(n1004) );
  NAND2X0 U823 ( .IN1(n1006), .IN2(n1007), .QN(n6092) );
  NAND2X0 U824 ( .IN1(P1_N4890), .IN2(P1_N5562), .QN(n1007) );
  NAND2X0 U825 ( .IN1(n7287), .IN2(n8938), .QN(n1006) );
  NAND2X0 U826 ( .IN1(n1008), .IN2(n1009), .QN(n6093) );
  NAND2X0 U827 ( .IN1(P1_N4889), .IN2(P1_N5562), .QN(n1009) );
  NAND2X0 U828 ( .IN1(n7287), .IN2(n8942), .QN(n1008) );
  NAND2X0 U829 ( .IN1(n1010), .IN2(n1011), .QN(n6094) );
  NAND2X0 U830 ( .IN1(P1_N4888), .IN2(P1_N5562), .QN(n1011) );
  NAND2X0 U831 ( .IN1(n7287), .IN2(n8946), .QN(n1010) );
  NAND2X0 U832 ( .IN1(n1012), .IN2(n1013), .QN(n6095) );
  NAND2X0 U833 ( .IN1(P1_N4887), .IN2(P1_N5562), .QN(n1013) );
  NAND2X0 U834 ( .IN1(n7287), .IN2(n8950), .QN(n1012) );
  NAND2X0 U835 ( .IN1(n1014), .IN2(n1015), .QN(n6096) );
  NAND2X0 U836 ( .IN1(P1_N4886), .IN2(P1_N5562), .QN(n1015) );
  NAND2X0 U837 ( .IN1(n7287), .IN2(n8954), .QN(n1014) );
  NAND2X0 U838 ( .IN1(n1016), .IN2(n1017), .QN(n6097) );
  NAND2X0 U839 ( .IN1(P1_N4885), .IN2(P1_N5562), .QN(n1017) );
  NAND2X0 U840 ( .IN1(n7287), .IN2(n8958), .QN(n1016) );
  NAND2X0 U841 ( .IN1(n1018), .IN2(n1019), .QN(n6098) );
  NAND2X0 U842 ( .IN1(P1_N4884), .IN2(P1_N5562), .QN(n1019) );
  NAND2X0 U843 ( .IN1(n7287), .IN2(n8962), .QN(n1018) );
  NAND2X0 U844 ( .IN1(n1020), .IN2(n1021), .QN(n6099) );
  NAND2X0 U845 ( .IN1(P1_N4883), .IN2(P1_N5562), .QN(n1021) );
  NAND2X0 U846 ( .IN1(n7287), .IN2(n8966), .QN(n1020) );
  NAND2X0 U847 ( .IN1(n1022), .IN2(n1023), .QN(n6100) );
  NAND2X0 U848 ( .IN1(P1_N4882), .IN2(P1_N5562), .QN(n1023) );
  NAND2X0 U849 ( .IN1(n7287), .IN2(n8970), .QN(n1022) );
  NAND2X0 U850 ( .IN1(n1024), .IN2(n1025), .QN(n6101) );
  NAND2X0 U851 ( .IN1(P1_N4881), .IN2(P1_N5562), .QN(n1025) );
  NAND2X0 U852 ( .IN1(n7287), .IN2(n8974), .QN(n1024) );
  NAND2X0 U853 ( .IN1(n1026), .IN2(n1027), .QN(n6102) );
  NAND2X0 U854 ( .IN1(P1_N4880), .IN2(P1_N5562), .QN(n1027) );
  NAND2X0 U855 ( .IN1(n7287), .IN2(n8978), .QN(n1026) );
  NAND2X0 U856 ( .IN1(n1028), .IN2(n1029), .QN(n6103) );
  NAND2X0 U857 ( .IN1(P1_N4879), .IN2(P1_N5562), .QN(n1029) );
  NAND2X0 U858 ( .IN1(n7287), .IN2(n8982), .QN(n1028) );
  NAND2X0 U859 ( .IN1(n1030), .IN2(n1031), .QN(n6104) );
  NAND2X0 U860 ( .IN1(P1_N4878), .IN2(P1_N5562), .QN(n1031) );
  NAND2X0 U861 ( .IN1(n7287), .IN2(n8986), .QN(n1030) );
  NAND2X0 U862 ( .IN1(n1032), .IN2(n1033), .QN(n6105) );
  NAND2X0 U863 ( .IN1(P1_N4877), .IN2(P1_N5562), .QN(n1033) );
  NAND2X0 U864 ( .IN1(n7287), .IN2(n8990), .QN(n1032) );
  NAND2X0 U865 ( .IN1(n1034), .IN2(n1035), .QN(n6106) );
  NAND2X0 U866 ( .IN1(P1_N4876), .IN2(P1_N5562), .QN(n1035) );
  NAND2X0 U867 ( .IN1(n7287), .IN2(n8994), .QN(n1034) );
  NAND2X0 U868 ( .IN1(n1036), .IN2(n1037), .QN(n6107) );
  NAND2X0 U869 ( .IN1(P1_N4875), .IN2(P1_N5562), .QN(n1037) );
  NAND2X0 U870 ( .IN1(n7287), .IN2(n8998), .QN(n1036) );
  NAND2X0 U871 ( .IN1(n1038), .IN2(n1039), .QN(n6108) );
  NAND2X0 U872 ( .IN1(P1_N4874), .IN2(P1_N5562), .QN(n1039) );
  NAND2X0 U873 ( .IN1(n7287), .IN2(n9002), .QN(n1038) );
  NAND2X0 U874 ( .IN1(n1040), .IN2(n1041), .QN(n6109) );
  NAND2X0 U875 ( .IN1(P1_N4873), .IN2(P1_N5562), .QN(n1041) );
  NAND2X0 U876 ( .IN1(n7287), .IN2(n9006), .QN(n1040) );
  NAND2X0 U878 ( .IN1(n1042), .IN2(n1043), .QN(n6110) );
  NAND2X0 U879 ( .IN1(n6725), .IN2(n10129), .QN(n1043) );
  NAND2X0 U880 ( .IN1(P1_N5552), .IN2(P1_N5548), .QN(n1042) );
  NAND2X0 U881 ( .IN1(n1045), .IN2(n1046), .QN(n6111) );
  NAND2X0 U882 ( .IN1(n6725), .IN2(n10125), .QN(n1046) );
  NAND2X0 U883 ( .IN1(P1_N5551), .IN2(P1_N5548), .QN(n1045) );
  NAND2X0 U884 ( .IN1(n1047), .IN2(n1048), .QN(n6112) );
  NAND2X0 U885 ( .IN1(n6725), .IN2(n10145), .QN(n1048) );
  NAND2X0 U886 ( .IN1(P1_N5550), .IN2(P1_N5548), .QN(n1047) );
  NAND2X0 U887 ( .IN1(n1049), .IN2(n1050), .QN(n6113) );
  NAND2X0 U888 ( .IN1(n6725), .IN2(n10373), .QN(n1050) );
  NAND2X0 U889 ( .IN1(P1_N5549), .IN2(P1_N5548), .QN(n1049) );
  NAND2X0 U704 ( .IN1(n7299), .IN2(n9026), .QN(n925) );
  NAND2X0 U705 ( .IN1(n927), .IN2(n928), .QN(n6053) );
  NAND2X0 U706 ( .IN1(P1_N4899), .IN2(P1_N5563), .QN(n928) );
  NAND2X0 U707 ( .IN1(n7299), .IN2(n9030), .QN(n927) );
  NAND2X0 U708 ( .IN1(n929), .IN2(n930), .QN(n6054) );
  NAND2X0 U709 ( .IN1(P1_N4898), .IN2(P1_N5563), .QN(n930) );
  NAND2X0 U710 ( .IN1(n7299), .IN2(n9034), .QN(n929) );
  NAND2X0 U711 ( .IN1(n931), .IN2(n932), .QN(n6055) );
  NAND2X0 U712 ( .IN1(P1_N4897), .IN2(P1_N5563), .QN(n932) );
  NAND2X0 U713 ( .IN1(n7299), .IN2(n9038), .QN(n931) );
  NAND2X0 U714 ( .IN1(n933), .IN2(n934), .QN(n6056) );
  NAND2X0 U715 ( .IN1(P1_N4896), .IN2(P1_N5563), .QN(n934) );
  NAND2X0 U716 ( .IN1(n7299), .IN2(n9042), .QN(n933) );
  NAND2X0 U717 ( .IN1(n935), .IN2(n936), .QN(n6057) );
  NAND2X0 U718 ( .IN1(P1_N4895), .IN2(P1_N5563), .QN(n936) );
  NAND2X0 U719 ( .IN1(n7299), .IN2(n9046), .QN(n935) );
  NAND2X0 U720 ( .IN1(n937), .IN2(n938), .QN(n6058) );
  NAND2X0 U721 ( .IN1(P1_N4894), .IN2(P1_N5563), .QN(n938) );
  NAND2X0 U722 ( .IN1(n7299), .IN2(n9050), .QN(n937) );
  NAND2X0 U723 ( .IN1(n939), .IN2(n940), .QN(n6059) );
  NAND2X0 U724 ( .IN1(P1_N4893), .IN2(P1_N5563), .QN(n940) );
  NAND2X0 U725 ( .IN1(n7299), .IN2(n9054), .QN(n939) );
  NAND2X0 U726 ( .IN1(n941), .IN2(n942), .QN(n6060) );
  NAND2X0 U727 ( .IN1(P1_N4892), .IN2(P1_N5563), .QN(n942) );
  NAND2X0 U728 ( .IN1(n7299), .IN2(n9493), .QN(n941) );
  NAND2X0 U729 ( .IN1(n943), .IN2(n944), .QN(n6061) );
  NAND2X0 U730 ( .IN1(P1_N4891), .IN2(P1_N5563), .QN(n944) );
  NAND2X0 U731 ( .IN1(n7299), .IN2(n9693), .QN(n943) );
  NAND2X0 U732 ( .IN1(n945), .IN2(n946), .QN(n6062) );
  NAND2X0 U733 ( .IN1(P1_N4890), .IN2(P1_N5563), .QN(n946) );
  NAND2X0 U734 ( .IN1(n7299), .IN2(n9697), .QN(n945) );
  NAND2X0 U735 ( .IN1(n947), .IN2(n948), .QN(n6063) );
  NAND2X0 U736 ( .IN1(P1_N4889), .IN2(P1_N5563), .QN(n948) );
  NAND2X0 U737 ( .IN1(n7299), .IN2(n9701), .QN(n947) );
  NAND2X0 U738 ( .IN1(n949), .IN2(n950), .QN(n6064) );
  NAND2X0 U739 ( .IN1(P1_N4888), .IN2(P1_N5563), .QN(n950) );
  NAND2X0 U740 ( .IN1(n7299), .IN2(n9705), .QN(n949) );
  NAND2X0 U741 ( .IN1(n951), .IN2(n952), .QN(n6065) );
  NAND2X0 U742 ( .IN1(P1_N4887), .IN2(P1_N5563), .QN(n952) );
  NAND2X0 U743 ( .IN1(n7299), .IN2(n9709), .QN(n951) );
  NAND2X0 U744 ( .IN1(n953), .IN2(n954), .QN(n6066) );
  NAND2X0 U745 ( .IN1(P1_N4886), .IN2(P1_N5563), .QN(n954) );
  NAND2X0 U746 ( .IN1(n7299), .IN2(n9713), .QN(n953) );
  NAND2X0 U747 ( .IN1(n955), .IN2(n956), .QN(n6067) );
  NAND2X0 U748 ( .IN1(P1_N4885), .IN2(P1_N5563), .QN(n956) );
  NAND2X0 U749 ( .IN1(n7299), .IN2(n9717), .QN(n955) );
  NAND2X0 U750 ( .IN1(n957), .IN2(n958), .QN(n6068) );
  NAND2X0 U751 ( .IN1(P1_N4884), .IN2(P1_N5563), .QN(n958) );
  NAND2X0 U752 ( .IN1(n7299), .IN2(n9721), .QN(n957) );
  NAND2X0 U753 ( .IN1(n959), .IN2(n960), .QN(n6069) );
  NAND2X0 U754 ( .IN1(P1_N4883), .IN2(P1_N5563), .QN(n960) );
  NAND2X0 U755 ( .IN1(n7299), .IN2(n9725), .QN(n959) );
  NAND2X0 U756 ( .IN1(n961), .IN2(n962), .QN(n6070) );
  NAND2X0 U757 ( .IN1(P1_N4882), .IN2(P1_N5563), .QN(n962) );
  NAND2X0 U758 ( .IN1(n7299), .IN2(n9729), .QN(n961) );
  NAND2X0 U759 ( .IN1(n963), .IN2(n964), .QN(n6071) );
  NAND2X0 U760 ( .IN1(P1_N4881), .IN2(P1_N5563), .QN(n964) );
  NAND2X0 U761 ( .IN1(n7299), .IN2(n9733), .QN(n963) );
  NAND2X0 U762 ( .IN1(n965), .IN2(n966), .QN(n6072) );
  NAND2X0 U763 ( .IN1(P1_N4880), .IN2(P1_N5563), .QN(n966) );
  NAND2X0 U764 ( .IN1(n7299), .IN2(n9737), .QN(n965) );
  NAND2X0 U765 ( .IN1(n967), .IN2(n968), .QN(n6073) );
  NAND2X0 U766 ( .IN1(P1_N4879), .IN2(P1_N5563), .QN(n968) );
  NAND2X0 U767 ( .IN1(n7299), .IN2(n9741), .QN(n967) );
  NAND2X0 U768 ( .IN1(n969), .IN2(n970), .QN(n6074) );
  NAND2X0 U769 ( .IN1(P1_N4878), .IN2(P1_N5563), .QN(n970) );
  NAND2X0 U770 ( .IN1(n7299), .IN2(n9745), .QN(n969) );
  NAND2X0 U771 ( .IN1(n971), .IN2(n972), .QN(n6075) );
  NAND2X0 U772 ( .IN1(P1_N4877), .IN2(P1_N5563), .QN(n972) );
  NAND2X0 U773 ( .IN1(n7299), .IN2(n9749), .QN(n971) );
  NAND2X0 U774 ( .IN1(n973), .IN2(n974), .QN(n6076) );
  NAND2X0 U775 ( .IN1(P1_N4876), .IN2(P1_N5563), .QN(n974) );
  NAND2X0 U776 ( .IN1(n7299), .IN2(n9753), .QN(n973) );
  NAND2X0 U777 ( .IN1(n975), .IN2(n976), .QN(n6077) );
  NAND2X0 U778 ( .IN1(P1_N4875), .IN2(P1_N5563), .QN(n976) );
  NAND2X0 U779 ( .IN1(n7299), .IN2(n9757), .QN(n975) );
  NAND2X0 U780 ( .IN1(n977), .IN2(n978), .QN(n6078) );
  NAND2X0 U781 ( .IN1(P1_N4874), .IN2(P1_N5563), .QN(n978) );
  NAND2X0 U782 ( .IN1(n7299), .IN2(n9761), .QN(n977) );
  NAND2X0 U783 ( .IN1(n979), .IN2(n980), .QN(n6079) );
  NAND2X0 U784 ( .IN1(P1_N4873), .IN2(P1_N5563), .QN(n980) );
  NAND2X0 U785 ( .IN1(n7299), .IN2(n981), .QN(n979) );
  NAND2X0 U787 ( .IN1(n982), .IN2(n983), .QN(n6080) );
  NAND2X0 U788 ( .IN1(P1_N4902), .IN2(P1_N5562), .QN(n983) );
  NAND2X0 U789 ( .IN1(n7287), .IN2(n8890), .QN(n982) );
  NAND2X0 U790 ( .IN1(n984), .IN2(n985), .QN(n6081) );
  NAND2X0 U791 ( .IN1(P1_N4901), .IN2(P1_N5562), .QN(n985) );
  NAND2X0 U792 ( .IN1(n7287), .IN2(n8894), .QN(n984) );
  NAND2X0 U793 ( .IN1(n986), .IN2(n987), .QN(n6082) );
  NAND2X0 U794 ( .IN1(P1_N4900), .IN2(P1_N5562), .QN(n987) );
  NAND2X0 U795 ( .IN1(n7287), .IN2(n8898), .QN(n986) );
  NAND2X0 U796 ( .IN1(n988), .IN2(n989), .QN(n6083) );
  NAND2X0 U611 ( .IN1(n864), .IN2(n865), .QN(n6022) );
  NAND2X0 U612 ( .IN1(P1_N4933), .IN2(P1_N5564), .QN(n865) );
  NAND2X0 U613 ( .IN1(n7295), .IN2(n9066), .QN(n864) );
  NAND2X0 U614 ( .IN1(n866), .IN2(n867), .QN(n6023) );
  NAND2X0 U615 ( .IN1(P1_N4932), .IN2(P1_N5564), .QN(n867) );
  NAND2X0 U616 ( .IN1(n7295), .IN2(n9070), .QN(n866) );
  NAND2X0 U617 ( .IN1(n868), .IN2(n869), .QN(n6024) );
  NAND2X0 U618 ( .IN1(P1_N4931), .IN2(P1_N5564), .QN(n869) );
  NAND2X0 U619 ( .IN1(n7295), .IN2(n9074), .QN(n868) );
  NAND2X0 U620 ( .IN1(n870), .IN2(n871), .QN(n6025) );
  NAND2X0 U621 ( .IN1(P1_N4930), .IN2(P1_N5564), .QN(n871) );
  NAND2X0 U622 ( .IN1(n7295), .IN2(n9078), .QN(n870) );
  NAND2X0 U623 ( .IN1(n872), .IN2(n873), .QN(n6026) );
  NAND2X0 U624 ( .IN1(P1_N4929), .IN2(P1_N5564), .QN(n873) );
  NAND2X0 U625 ( .IN1(n7295), .IN2(n9082), .QN(n872) );
  NAND2X0 U626 ( .IN1(n874), .IN2(n875), .QN(n6027) );
  NAND2X0 U627 ( .IN1(P1_N4928), .IN2(P1_N5564), .QN(n875) );
  NAND2X0 U628 ( .IN1(n7295), .IN2(n9086), .QN(n874) );
  NAND2X0 U629 ( .IN1(n876), .IN2(n877), .QN(n6028) );
  NAND2X0 U630 ( .IN1(P1_N4927), .IN2(P1_N5564), .QN(n877) );
  NAND2X0 U631 ( .IN1(n7295), .IN2(n9090), .QN(n876) );
  NAND2X0 U632 ( .IN1(n878), .IN2(n879), .QN(n6029) );
  NAND2X0 U633 ( .IN1(P1_N4926), .IN2(P1_N5564), .QN(n879) );
  NAND2X0 U634 ( .IN1(n7295), .IN2(n9094), .QN(n878) );
  NAND2X0 U635 ( .IN1(n880), .IN2(n881), .QN(n6030) );
  NAND2X0 U636 ( .IN1(P1_N4925), .IN2(P1_N5564), .QN(n881) );
  NAND2X0 U637 ( .IN1(n7295), .IN2(n9497), .QN(n880) );
  NAND2X0 U638 ( .IN1(n882), .IN2(n883), .QN(n6031) );
  NAND2X0 U639 ( .IN1(P1_N4924), .IN2(P1_N5564), .QN(n883) );
  NAND2X0 U640 ( .IN1(n7295), .IN2(n9765), .QN(n882) );
  NAND2X0 U641 ( .IN1(n884), .IN2(n885), .QN(n6032) );
  NAND2X0 U642 ( .IN1(P1_N4923), .IN2(P1_N5564), .QN(n885) );
  NAND2X0 U643 ( .IN1(n7295), .IN2(n9769), .QN(n884) );
  NAND2X0 U644 ( .IN1(n886), .IN2(n887), .QN(n6033) );
  NAND2X0 U645 ( .IN1(P1_N4922), .IN2(P1_N5564), .QN(n887) );
  NAND2X0 U646 ( .IN1(n7295), .IN2(n9773), .QN(n886) );
  NAND2X0 U647 ( .IN1(n888), .IN2(n889), .QN(n6034) );
  NAND2X0 U648 ( .IN1(P1_N4921), .IN2(P1_N5564), .QN(n889) );
  NAND2X0 U649 ( .IN1(n7295), .IN2(n9777), .QN(n888) );
  NAND2X0 U650 ( .IN1(n890), .IN2(n891), .QN(n6035) );
  NAND2X0 U651 ( .IN1(P1_N4920), .IN2(P1_N5564), .QN(n891) );
  NAND2X0 U652 ( .IN1(n7295), .IN2(n9781), .QN(n890) );
  NAND2X0 U653 ( .IN1(n892), .IN2(n893), .QN(n6036) );
  NAND2X0 U654 ( .IN1(P1_N4919), .IN2(P1_N5564), .QN(n893) );
  NAND2X0 U655 ( .IN1(n7295), .IN2(n9785), .QN(n892) );
  NAND2X0 U656 ( .IN1(n894), .IN2(n895), .QN(n6037) );
  NAND2X0 U657 ( .IN1(P1_N4918), .IN2(P1_N5564), .QN(n895) );
  NAND2X0 U658 ( .IN1(n7295), .IN2(n9789), .QN(n894) );
  NAND2X0 U659 ( .IN1(n896), .IN2(n897), .QN(n6038) );
  NAND2X0 U660 ( .IN1(P1_N4917), .IN2(P1_N5564), .QN(n897) );
  NAND2X0 U661 ( .IN1(n7295), .IN2(n9793), .QN(n896) );
  NAND2X0 U662 ( .IN1(n898), .IN2(n899), .QN(n6039) );
  NAND2X0 U663 ( .IN1(P1_N4916), .IN2(P1_N5564), .QN(n899) );
  NAND2X0 U664 ( .IN1(n7295), .IN2(n9797), .QN(n898) );
  NAND2X0 U665 ( .IN1(n900), .IN2(n901), .QN(n6040) );
  NAND2X0 U666 ( .IN1(P1_N4915), .IN2(P1_N5564), .QN(n901) );
  NAND2X0 U667 ( .IN1(n7295), .IN2(n9801), .QN(n900) );
  NAND2X0 U668 ( .IN1(n902), .IN2(n903), .QN(n6041) );
  NAND2X0 U669 ( .IN1(P1_N4914), .IN2(P1_N5564), .QN(n903) );
  NAND2X0 U670 ( .IN1(n7295), .IN2(n9805), .QN(n902) );
  NAND2X0 U671 ( .IN1(n904), .IN2(n905), .QN(n6042) );
  NAND2X0 U672 ( .IN1(P1_N4913), .IN2(P1_N5564), .QN(n905) );
  NAND2X0 U673 ( .IN1(n7295), .IN2(n9809), .QN(n904) );
  NAND2X0 U674 ( .IN1(n906), .IN2(n907), .QN(n6043) );
  NAND2X0 U675 ( .IN1(P1_N4912), .IN2(P1_N5564), .QN(n907) );
  NAND2X0 U676 ( .IN1(n7295), .IN2(n9813), .QN(n906) );
  NAND2X0 U677 ( .IN1(n908), .IN2(n909), .QN(n6044) );
  NAND2X0 U678 ( .IN1(P1_N4911), .IN2(P1_N5564), .QN(n909) );
  NAND2X0 U679 ( .IN1(n7295), .IN2(n9817), .QN(n908) );
  NAND2X0 U680 ( .IN1(n910), .IN2(n911), .QN(n6045) );
  NAND2X0 U681 ( .IN1(P1_N4910), .IN2(P1_N5564), .QN(n911) );
  NAND2X0 U682 ( .IN1(n7295), .IN2(n9821), .QN(n910) );
  NAND2X0 U683 ( .IN1(n912), .IN2(n913), .QN(n6046) );
  NAND2X0 U684 ( .IN1(P1_N4909), .IN2(P1_N5564), .QN(n913) );
  NAND2X0 U685 ( .IN1(n7295), .IN2(n9825), .QN(n912) );
  NAND2X0 U686 ( .IN1(n914), .IN2(n915), .QN(n6047) );
  NAND2X0 U687 ( .IN1(P1_N4908), .IN2(P1_N5564), .QN(n915) );
  NAND2X0 U688 ( .IN1(n7295), .IN2(n9829), .QN(n914) );
  NAND2X0 U689 ( .IN1(n916), .IN2(n917), .QN(n6048) );
  NAND2X0 U690 ( .IN1(P1_N4907), .IN2(P1_N5564), .QN(n917) );
  NAND2X0 U691 ( .IN1(n7295), .IN2(n9833), .QN(n916) );
  NAND2X0 U692 ( .IN1(n918), .IN2(n919), .QN(n6049) );
  NAND2X0 U693 ( .IN1(P1_N4906), .IN2(P1_N5564), .QN(n919) );
  NAND2X0 U694 ( .IN1(n7295), .IN2(n920), .QN(n918) );
  NAND2X0 U696 ( .IN1(n921), .IN2(n922), .QN(n6050) );
  NAND2X0 U697 ( .IN1(P1_N4902), .IN2(P1_N5563), .QN(n922) );
  NAND2X0 U698 ( .IN1(n7299), .IN2(n9018), .QN(n921) );
  NAND2X0 U699 ( .IN1(n923), .IN2(n924), .QN(n6051) );
  NAND2X0 U700 ( .IN1(P1_N4901), .IN2(P1_N5563), .QN(n924) );
  NAND2X0 U701 ( .IN1(n7299), .IN2(n9022), .QN(n923) );
  NAND2X0 U702 ( .IN1(n925), .IN2(n926), .QN(n6052) );
  NAND2X0 U703 ( .IN1(P1_N4900), .IN2(P1_N5563), .QN(n926) );
  NAND2X0 U518 ( .IN1(n7031), .IN2(n9875), .QN(n801) );
  NAND2X0 U519 ( .IN1(n803), .IN2(n804), .QN(n5992) );
  NAND2X0 U520 ( .IN1(n7075), .IN2(P1_N5554), .QN(n804) );
  NAND2X0 U521 ( .IN1(n7031), .IN2(n9879), .QN(n803) );
  NAND2X0 U522 ( .IN1(n805), .IN2(n806), .QN(n5993) );
  NAND2X0 U523 ( .IN1(P1_N5155), .IN2(P1_N5554), .QN(n806) );
  NAND2X0 U524 ( .IN1(n7031), .IN2(n9883), .QN(n805) );
  NAND2X0 U525 ( .IN1(n807), .IN2(n808), .QN(n5994) );
  NAND2X0 U526 ( .IN1(P1_N5154), .IN2(P1_N5554), .QN(n808) );
  NAND2X0 U527 ( .IN1(n7031), .IN2(n9887), .QN(n807) );
  NAND2X0 U528 ( .IN1(n809), .IN2(n810), .QN(n5995) );
  NAND2X0 U529 ( .IN1(P1_N5153), .IN2(P1_N5554), .QN(n810) );
  NAND2X0 U530 ( .IN1(n7031), .IN2(n9891), .QN(n809) );
  NAND2X0 U531 ( .IN1(n811), .IN2(n812), .QN(n5996) );
  NAND2X0 U532 ( .IN1(n7041), .IN2(P1_N5554), .QN(n812) );
  NAND2X0 U533 ( .IN1(n7031), .IN2(n9895), .QN(n811) );
  NAND2X0 U534 ( .IN1(n813), .IN2(n814), .QN(n5997) );
  NAND2X0 U535 ( .IN1(n7046), .IN2(P1_N5554), .QN(n814) );
  NAND2X0 U536 ( .IN1(n7031), .IN2(n9899), .QN(n813) );
  NAND2X0 U537 ( .IN1(n815), .IN2(n816), .QN(n5998) );
  NAND2X0 U538 ( .IN1(P1_N5150), .IN2(P1_N5554), .QN(n816) );
  NAND2X0 U539 ( .IN1(n7031), .IN2(n9333), .QN(n815) );
  NAND2X0 U540 ( .IN1(n817), .IN2(n818), .QN(n5999) );
  NAND2X0 U541 ( .IN1(n7031), .IN2(n9385), .QN(n818) );
  NAND2X0 U543 ( .IN1(P1_N5554), .IN2(n7034), .QN(n817) );
  NAND2X0 U544 ( .IN1(n819), .IN2(n820), .QN(n6000) );
  NAND2X0 U545 ( .IN1(n7284), .IN2(n18245), .QN(n820) );
  NAND2X0 U546 ( .IN1(P1_N5517), .IN2(P1_N5497), .QN(n819) );
  NAND2X0 U547 ( .IN1(n822), .IN2(n823), .QN(n6001) );
  NAND2X0 U548 ( .IN1(n7284), .IN2(n9565), .QN(n823) );
  NAND2X0 U549 ( .IN1(P1_N5516), .IN2(P1_N5497), .QN(n822) );
  NAND2X0 U550 ( .IN1(n824), .IN2(n825), .QN(n6002) );
  NAND2X0 U551 ( .IN1(n7284), .IN2(n9569), .QN(n825) );
  NAND2X0 U552 ( .IN1(P1_N5515), .IN2(P1_N5497), .QN(n824) );
  NAND2X0 U553 ( .IN1(n826), .IN2(n827), .QN(n6003) );
  NAND2X0 U554 ( .IN1(n7284), .IN2(n9573), .QN(n827) );
  NAND2X0 U555 ( .IN1(P1_N5514), .IN2(P1_N5497), .QN(n826) );
  NAND2X0 U556 ( .IN1(n828), .IN2(n829), .QN(n6004) );
  NAND2X0 U557 ( .IN1(n7284), .IN2(n9577), .QN(n829) );
  NAND2X0 U558 ( .IN1(P1_N5513), .IN2(P1_N5497), .QN(n828) );
  NAND2X0 U559 ( .IN1(n830), .IN2(n831), .QN(n6005) );
  NAND2X0 U560 ( .IN1(n7284), .IN2(n9581), .QN(n831) );
  NAND2X0 U561 ( .IN1(P1_N5512), .IN2(P1_N5497), .QN(n830) );
  NAND2X0 U562 ( .IN1(n832), .IN2(n833), .QN(n6006) );
  NAND2X0 U563 ( .IN1(n7284), .IN2(n9585), .QN(n833) );
  NAND2X0 U564 ( .IN1(P1_N5511), .IN2(P1_N5497), .QN(n832) );
  NAND2X0 U565 ( .IN1(n834), .IN2(n835), .QN(n6007) );
  NAND2X0 U566 ( .IN1(n7284), .IN2(n9589), .QN(n835) );
  NAND2X0 U567 ( .IN1(P1_N5510), .IN2(P1_N5497), .QN(n834) );
  NAND2X0 U568 ( .IN1(n836), .IN2(n837), .QN(n6008) );
  NAND2X0 U569 ( .IN1(n7284), .IN2(n9593), .QN(n837) );
  NAND2X0 U570 ( .IN1(P1_N5509), .IN2(P1_N5497), .QN(n836) );
  NAND2X0 U571 ( .IN1(n838), .IN2(n839), .QN(n6009) );
  NAND2X0 U572 ( .IN1(n7284), .IN2(n9597), .QN(n839) );
  NAND2X0 U573 ( .IN1(P1_N5508), .IN2(P1_N5497), .QN(n838) );
  NAND2X0 U574 ( .IN1(n840), .IN2(n841), .QN(n6010) );
  NAND2X0 U575 ( .IN1(n7284), .IN2(n9601), .QN(n841) );
  NAND2X0 U576 ( .IN1(P1_N5507), .IN2(P1_N5497), .QN(n840) );
  NAND2X0 U577 ( .IN1(n842), .IN2(n843), .QN(n6011) );
  NAND2X0 U578 ( .IN1(n7284), .IN2(n9605), .QN(n843) );
  NAND2X0 U579 ( .IN1(P1_N5506), .IN2(P1_N5497), .QN(n842) );
  NAND2X0 U580 ( .IN1(n844), .IN2(n845), .QN(n6012) );
  NAND2X0 U581 ( .IN1(n7284), .IN2(n9609), .QN(n845) );
  NAND2X0 U582 ( .IN1(P1_N5505), .IN2(P1_N5497), .QN(n844) );
  NAND2X0 U583 ( .IN1(n846), .IN2(n847), .QN(n6013) );
  NAND2X0 U584 ( .IN1(n7284), .IN2(n9613), .QN(n847) );
  NAND2X0 U585 ( .IN1(P1_N5504), .IN2(P1_N5497), .QN(n846) );
  NAND2X0 U586 ( .IN1(n848), .IN2(n849), .QN(n6014) );
  NAND2X0 U587 ( .IN1(n7284), .IN2(n9617), .QN(n849) );
  NAND2X0 U588 ( .IN1(P1_N5503), .IN2(P1_N5497), .QN(n848) );
  NAND2X0 U589 ( .IN1(n850), .IN2(n851), .QN(n6015) );
  NAND2X0 U590 ( .IN1(n7284), .IN2(n9621), .QN(n851) );
  NAND2X0 U591 ( .IN1(P1_N5502), .IN2(P1_N5497), .QN(n850) );
  NAND2X0 U592 ( .IN1(n852), .IN2(n853), .QN(n6016) );
  NAND2X0 U593 ( .IN1(n7284), .IN2(n9625), .QN(n853) );
  NAND2X0 U594 ( .IN1(P1_N5501), .IN2(P1_N5497), .QN(n852) );
  NAND2X0 U595 ( .IN1(n854), .IN2(n855), .QN(n6017) );
  NAND2X0 U596 ( .IN1(n7284), .IN2(n9629), .QN(n855) );
  NAND2X0 U597 ( .IN1(P1_N5500), .IN2(P1_N5497), .QN(n854) );
  NAND2X0 U598 ( .IN1(n856), .IN2(n857), .QN(n6018) );
  NAND2X0 U599 ( .IN1(n7284), .IN2(n9318), .QN(n857) );
  NAND2X0 U600 ( .IN1(P1_N5499), .IN2(P1_N5497), .QN(n856) );
  NAND2X0 U601 ( .IN1(n858), .IN2(n859), .QN(n6019) );
  NAND2X0 U602 ( .IN1(n7284), .IN2(n9329), .QN(n859) );
  NAND2X0 U604 ( .IN1(P1_N5498), .IN2(P1_N5497), .QN(n858) );
  NAND2X0 U605 ( .IN1(n860), .IN2(n861), .QN(n6020) );
  NAND2X0 U606 ( .IN1(P1_N4935), .IN2(P1_N5564), .QN(n861) );
  NAND2X0 U607 ( .IN1(n7295), .IN2(n9058), .QN(n860) );
  NAND2X0 U608 ( .IN1(n862), .IN2(n863), .QN(n6021) );
  NAND2X0 U609 ( .IN1(P1_N4934), .IN2(P1_N5564), .QN(n863) );
  NAND2X0 U610 ( .IN1(n7295), .IN2(n9062), .QN(n862) );
  NAND2X0 U340 ( .IN1(n738), .IN2(n739), .QN(n5962) );
  NAND2X0 U341 ( .IN1(n7299), .IN2(n9014), .QN(n739) );
  NAND2X0 U342 ( .IN1(P1_N5563), .IN2(n7445), .QN(n738) );
  NAND2X0 U343 ( .IN1(n741), .IN2(n742), .QN(n5963) );
  NAND2X0 U344 ( .IN1(n7287), .IN2(n9310), .QN(n742) );
  NAND2X0 U345 ( .IN1(P1_N5562), .IN2(n7444), .QN(n741) );
  NAND2X0 U347 ( .IN1(n744), .IN2(n745), .QN(n5964) );
  NAND2X0 U348 ( .IN1(n7287), .IN2(n9314), .QN(n745) );
  NAND2X0 U349 ( .IN1(P1_N5562), .IN2(n7445), .QN(n744) );
  NAND2X0 U351 ( .IN1(n746), .IN2(n747), .QN(n5965) );
  NAND2X0 U352 ( .IN1(n7031), .IN2(n9345), .QN(n747) );
  NAND2X0 U353 ( .IN1(P1_N5554), .IN2(n7052), .QN(n746) );
  NAND2X0 U354 ( .IN1(n749), .IN2(n750), .QN(n5966) );
  NAND2X0 U355 ( .IN1(P1_N497), .IN2(P1_N5554), .QN(n750) );
  NAND2X0 U356 ( .IN1(n7031), .IN2(n10103), .QN(n749) );
  NAND2X0 U357 ( .IN1(n751), .IN2(n752), .QN(n5967) );
  NAND2X0 U358 ( .IN1(P1_N5178), .IN2(P1_N5554), .QN(n752) );
  NAND2X0 U359 ( .IN1(n7031), .IN2(n10095), .QN(n751) );
  NAND2X0 U360 ( .IN1(n753), .IN2(n754), .QN(n5968) );
  NAND2X0 U361 ( .IN1(P1_N5560), .IN2(P1_N531), .QN(n754) );
  NAND2X0 U372 ( .IN1(n755), .IN2(n6619), .QN(n753) );
  NAND2X0 U391 ( .IN1(n756), .IN2(n757), .QN(n5969) );
  NAND2X0 U418 ( .IN1(P1_N530), .IN2(P1_N5560), .QN(n757) );
  NAND2X0 U420 ( .IN1(n755), .IN2(n6620), .QN(n756) );
  INVX0 U421 ( .ZN(n755), .INP(P1_N5560) );
  NAND2X0 U422 ( .IN1(n758), .IN2(n759), .QN(n5970) );
  NAND2X0 U423 ( .IN1(n6618), .IN2(n760), .QN(n759) );
  INVX0 U424 ( .ZN(n760), .INP(P1_N5561) );
  NAND2X0 U425 ( .IN1(P1_N5561), .IN2(n7443), .QN(n758) );
  NAND2X0 U428 ( .IN1(n761), .IN2(n762), .QN(n5971) );
  NAND2X0 U429 ( .IN1(P1_N5177), .IN2(P1_N5554), .QN(n762) );
  NAND2X0 U430 ( .IN1(n7031), .IN2(n9935), .QN(n761) );
  NAND2X0 U431 ( .IN1(n763), .IN2(n764), .QN(n5972) );
  NAND2X0 U448 ( .IN1(n7122), .IN2(P1_N5554), .QN(n764) );
  NAND2X0 U456 ( .IN1(n7031), .IN2(n9939), .QN(n763) );
  NAND2X0 U457 ( .IN1(n765), .IN2(n766), .QN(n5973) );
  NAND2X0 U458 ( .IN1(P1_N5175), .IN2(P1_N5554), .QN(n766) );
  NAND2X0 U459 ( .IN1(n7031), .IN2(n9943), .QN(n765) );
  NAND2X0 U460 ( .IN1(n767), .IN2(n768), .QN(n5974) );
  NAND2X0 U461 ( .IN1(P1_N5174), .IN2(P1_N5554), .QN(n768) );
  NAND2X0 U464 ( .IN1(n7031), .IN2(n9947), .QN(n767) );
  NAND2X0 U465 ( .IN1(n769), .IN2(n770), .QN(n5975) );
  NAND2X0 U466 ( .IN1(n7138), .IN2(P1_N5554), .QN(n770) );
  NAND2X0 U467 ( .IN1(n7031), .IN2(n9951), .QN(n769) );
  NAND2X0 U471 ( .IN1(n771), .IN2(n772), .QN(n5976) );
  NAND2X0 U472 ( .IN1(n7141), .IN2(P1_N5554), .QN(n772) );
  NAND2X0 U473 ( .IN1(n7031), .IN2(n9955), .QN(n771) );
  NAND2X0 U474 ( .IN1(n773), .IN2(n774), .QN(n5977) );
  NAND2X0 U475 ( .IN1(P1_N5171), .IN2(P1_N5554), .QN(n774) );
  NAND2X0 U476 ( .IN1(n7031), .IN2(n9959), .QN(n773) );
  NAND2X0 U477 ( .IN1(n775), .IN2(n776), .QN(n5978) );
  NAND2X0 U478 ( .IN1(n7093), .IN2(P1_N5554), .QN(n776) );
  NAND2X0 U479 ( .IN1(n7031), .IN2(n9963), .QN(n775) );
  NAND2X0 U480 ( .IN1(n777), .IN2(n778), .QN(n5979) );
  NAND2X0 U481 ( .IN1(n7096), .IN2(P1_N5554), .QN(n778) );
  NAND2X0 U482 ( .IN1(n7031), .IN2(n9967), .QN(n777) );
  NAND2X0 U483 ( .IN1(n779), .IN2(n780), .QN(n5980) );
  NAND2X0 U484 ( .IN1(n7099), .IN2(P1_N5554), .QN(n780) );
  NAND2X0 U485 ( .IN1(n7031), .IN2(n9971), .QN(n779) );
  NAND2X0 U486 ( .IN1(n781), .IN2(n782), .QN(n5981) );
  NAND2X0 U487 ( .IN1(n7103), .IN2(P1_N5554), .QN(n782) );
  NAND2X0 U488 ( .IN1(n7031), .IN2(n9975), .QN(n781) );
  NAND2X0 U489 ( .IN1(n783), .IN2(n784), .QN(n5982) );
  NAND2X0 U490 ( .IN1(n7106), .IN2(P1_N5554), .QN(n784) );
  NAND2X0 U491 ( .IN1(n7031), .IN2(n9979), .QN(n783) );
  NAND2X0 U492 ( .IN1(n785), .IN2(n786), .QN(n5983) );
  NAND2X0 U493 ( .IN1(n7110), .IN2(P1_N5554), .QN(n786) );
  NAND2X0 U494 ( .IN1(n7031), .IN2(n9983), .QN(n785) );
  NAND2X0 U495 ( .IN1(n787), .IN2(n788), .QN(n5984) );
  NAND2X0 U496 ( .IN1(n7113), .IN2(P1_N5554), .QN(n788) );
  NAND2X0 U497 ( .IN1(n7031), .IN2(n9987), .QN(n787) );
  NAND2X0 U498 ( .IN1(n789), .IN2(n790), .QN(n5985) );
  NAND2X0 U499 ( .IN1(n7116), .IN2(P1_N5554), .QN(n790) );
  NAND2X0 U500 ( .IN1(n7031), .IN2(n9991), .QN(n789) );
  NAND2X0 U501 ( .IN1(n791), .IN2(n792), .QN(n5986) );
  NAND2X0 U502 ( .IN1(P1_N5162), .IN2(P1_N5554), .QN(n792) );
  NAND2X0 U503 ( .IN1(n7031), .IN2(n9995), .QN(n791) );
  NAND2X0 U504 ( .IN1(n793), .IN2(n794), .QN(n5987) );
  NAND2X0 U505 ( .IN1(n7059), .IN2(P1_N5554), .QN(n794) );
  NAND2X0 U506 ( .IN1(n7031), .IN2(n9999), .QN(n793) );
  NAND2X0 U507 ( .IN1(n795), .IN2(n796), .QN(n5988) );
  NAND2X0 U508 ( .IN1(P1_N5160), .IN2(P1_N5554), .QN(n796) );
  NAND2X0 U509 ( .IN1(n7031), .IN2(n10003), .QN(n795) );
  NAND2X0 U510 ( .IN1(n797), .IN2(n798), .QN(n5989) );
  NAND2X0 U511 ( .IN1(n7066), .IN2(P1_N5554), .QN(n798) );
  NAND2X0 U512 ( .IN1(n7031), .IN2(n10007), .QN(n797) );
  NAND2X0 U513 ( .IN1(n799), .IN2(n800), .QN(n5990) );
  NAND2X0 U514 ( .IN1(P1_N5158), .IN2(P1_N5554), .QN(n800) );
  NAND2X0 U515 ( .IN1(n7031), .IN2(n9871), .QN(n799) );
  NAND2X0 U516 ( .IN1(n801), .IN2(n802), .QN(n5991) );
  NAND2X0 U517 ( .IN1(n7072), .IN2(P1_N5554), .QN(n802) );
  AND2X1 U247 ( .IN1(n666), .IN2(n667), .Q(n664) );
  NAND2X0 U248 ( .IN1(P2_N375), .IN2(n598), .QN(n667) );
  NAND2X0 U249 ( .IN1(P2_N4821), .IN2(n599), .QN(n666) );
  NAND2X0 U250 ( .IN1(n668), .IN2(n669), .QN(n1865) );
  NAND2X0 U251 ( .IN1(n2166), .IN2(n9537), .QN(n669) );
  AND2X1 U252 ( .IN1(n670), .IN2(n671), .Q(n668) );
  NAND2X0 U253 ( .IN1(P2_N374), .IN2(n598), .QN(n671) );
  NAND2X0 U254 ( .IN1(P2_N4820), .IN2(n599), .QN(n670) );
  NAND2X0 U255 ( .IN1(n672), .IN2(n673), .QN(n1867) );
  NAND2X0 U256 ( .IN1(n2166), .IN2(n9541), .QN(n673) );
  AND2X1 U257 ( .IN1(n674), .IN2(n675), .Q(n672) );
  NAND2X0 U258 ( .IN1(P2_N373), .IN2(n598), .QN(n675) );
  NAND2X0 U259 ( .IN1(P2_N4819), .IN2(n599), .QN(n674) );
  NAND2X0 U260 ( .IN1(n676), .IN2(n677), .QN(n1869) );
  NAND2X0 U261 ( .IN1(n2166), .IN2(n9545), .QN(n677) );
  AND2X1 U262 ( .IN1(n678), .IN2(n679), .Q(n676) );
  NAND2X0 U263 ( .IN1(P2_N372), .IN2(n598), .QN(n679) );
  NAND2X0 U264 ( .IN1(P2_N4818), .IN2(n599), .QN(n678) );
  NAND2X0 U265 ( .IN1(n680), .IN2(n681), .QN(n1871) );
  NAND2X0 U266 ( .IN1(n2166), .IN2(n9549), .QN(n681) );
  AND2X1 U267 ( .IN1(n682), .IN2(n683), .Q(n680) );
  NAND2X0 U268 ( .IN1(P2_N371), .IN2(n598), .QN(n683) );
  NAND2X0 U269 ( .IN1(P2_N4817), .IN2(n599), .QN(n682) );
  NAND2X0 U270 ( .IN1(n684), .IN2(n685), .QN(n1873) );
  NAND2X0 U271 ( .IN1(n2166), .IN2(n9553), .QN(n685) );
  AND2X1 U272 ( .IN1(n686), .IN2(n687), .Q(n684) );
  NAND2X0 U273 ( .IN1(P2_N370), .IN2(n598), .QN(n687) );
  NAND2X0 U274 ( .IN1(P2_N4816), .IN2(n599), .QN(n686) );
  NAND2X0 U275 ( .IN1(n688), .IN2(n689), .QN(n1875) );
  NAND2X0 U276 ( .IN1(n2166), .IN2(n9557), .QN(n689) );
  AND2X1 U277 ( .IN1(n690), .IN2(n691), .Q(n688) );
  NAND2X0 U278 ( .IN1(P2_N369), .IN2(n598), .QN(n691) );
  NAND2X0 U279 ( .IN1(P2_N4815), .IN2(n599), .QN(n690) );
  NAND2X0 U280 ( .IN1(n692), .IN2(n693), .QN(n1877) );
  NAND2X0 U281 ( .IN1(n2166), .IN2(n9397), .QN(n693) );
  AND2X1 U282 ( .IN1(n694), .IN2(n695), .Q(n692) );
  NAND2X0 U283 ( .IN1(P2_N368), .IN2(n598), .QN(n695) );
  NAND2X0 U284 ( .IN1(P2_N4814), .IN2(n599), .QN(n694) );
  NAND2X0 U285 ( .IN1(n696), .IN2(n697), .QN(n1879) );
  NAND2X0 U286 ( .IN1(n2166), .IN2(n6684), .QN(n697) );
  AND2X1 U287 ( .IN1(n698), .IN2(n699), .Q(n696) );
  NAND2X0 U288 ( .IN1(n18813), .IN2(n598), .QN(n699) );
  NAND2X0 U289 ( .IN1(P2_N4813), .IN2(n599), .QN(n698) );
  NAND2X0 U290 ( .IN1(n700), .IN2(n701), .QN(n1881) );
  NAND2X0 U291 ( .IN1(n2166), .IN2(n6683), .QN(n701) );
  AND2X1 U292 ( .IN1(n702), .IN2(n703), .Q(n700) );
  NAND2X0 U293 ( .IN1(n6683), .IN2(n598), .QN(n703) );
  NAND2X0 U294 ( .IN1(P2_N4812), .IN2(n599), .QN(n702) );
  NAND2X0 U295 ( .IN1(n704), .IN2(n705), .QN(n1883) );
  NAND2X0 U296 ( .IN1(n2166), .IN2(n6682), .QN(n705) );
  AND2X1 U297 ( .IN1(n706), .IN2(n707), .Q(n704) );
  NAND2X0 U298 ( .IN1(n6682), .IN2(n598), .QN(n707) );
  NAND2X0 U299 ( .IN1(P2_N4811), .IN2(n599), .QN(n706) );
  NAND2X0 U300 ( .IN1(n708), .IN2(n709), .QN(n1885) );
  NAND2X0 U301 ( .IN1(n6589), .IN2(n6681), .QN(n709) );
  AND2X1 U302 ( .IN1(n710), .IN2(n711), .Q(n708) );
  NAND2X0 U303 ( .IN1(n6681), .IN2(n598), .QN(n711) );
  NAND2X0 U305 ( .IN1(P2_N4810), .IN2(n599), .QN(n710) );
  INVX0 U307 ( .ZN(n4366), .INP(n4356) );
  NAND2X0 U308 ( .IN1(P1_N499), .IN2(n7414), .QN(n4356) );
  INVX0 U309 ( .ZN(n2459), .INP(n2452) );
  NAND2X0 U310 ( .IN1(P2_N499), .IN2(n7415), .QN(n2452) );
  NAND2X0 U311 ( .IN1(n712), .IN2(n713), .QN(n5953) );
  NAND2X0 U312 ( .IN1(P2_N5486), .IN2(P2_N4809), .QN(n713) );
  NAND2X0 U313 ( .IN1(n7303), .IN2(n9306), .QN(n712) );
  NAND2X0 U314 ( .IN1(n715), .IN2(n716), .QN(n5954) );
  NAND2X0 U315 ( .IN1(P2_N4808), .IN2(P2_N5486), .QN(n716) );
  NAND2X0 U316 ( .IN1(n7303), .IN2(n8870), .QN(n715) );
  NAND2X0 U317 ( .IN1(n717), .IN2(n718), .QN(n5955) );
  NAND2X0 U318 ( .IN1(n7291), .IN2(n9098), .QN(n718) );
  NAND2X0 U319 ( .IN1(P2_N5484), .IN2(n720), .QN(n717) );
  NAND2X0 U320 ( .IN1(n721), .IN2(n722), .QN(n5956) );
  NAND2X0 U321 ( .IN1(n7309), .IN2(n9222), .QN(n722) );
  NAND2X0 U322 ( .IN1(P2_N5485), .IN2(n720), .QN(n721) );
  INVX0 U323 ( .ZN(n720), .INP(n7446) );
  NAND2X0 U324 ( .IN1(n724), .IN2(n725), .QN(n5957) );
  NAND2X0 U325 ( .IN1(n7291), .IN2(n8874), .QN(n725) );
  NAND2X0 U326 ( .IN1(P2_N5484), .IN2(n726), .QN(n724) );
  NAND2X0 U327 ( .IN1(n727), .IN2(n728), .QN(n5958) );
  NAND2X0 U328 ( .IN1(n7309), .IN2(n8878), .QN(n728) );
  NAND2X0 U329 ( .IN1(P2_N5485), .IN2(n726), .QN(n727) );
  INVX0 U330 ( .ZN(n726), .INP(n7447) );
  NAND2X0 U331 ( .IN1(n729), .IN2(n730), .QN(n5959) );
  NAND2X0 U332 ( .IN1(P1_N5564), .IN2(n7444), .QN(n730) );
  NAND2X0 U333 ( .IN1(n7295), .IN2(n8886), .QN(n729) );
  NAND2X0 U334 ( .IN1(n732), .IN2(n733), .QN(n5960) );
  NAND2X0 U335 ( .IN1(n7445), .IN2(P1_N5564), .QN(n733) );
  NAND2X0 U336 ( .IN1(n7295), .IN2(n8882), .QN(n732) );
  NAND2X0 U337 ( .IN1(n734), .IN2(n735), .QN(n5961) );
  NAND2X0 U338 ( .IN1(n7299), .IN2(n9010), .QN(n735) );
  NAND2X0 U339 ( .IN1(P1_N5563), .IN2(n7444), .QN(n734) );
  NAND2X0 U154 ( .IN1(n6580), .IN2(n6621), .QN(n591) );
  AND2X1 U155 ( .IN1(n592), .IN2(n593), .Q(n590) );
  NAND2X0 U156 ( .IN1(n6621), .IN2(n480), .QN(n593) );
  NAND2X0 U158 ( .IN1(P1_N4938), .IN2(n481), .QN(n592) );
  NAND2X0 U160 ( .IN1(n594), .IN2(n595), .QN(n1829) );
  NAND2X0 U161 ( .IN1(n6589), .IN2(n9349), .QN(n595) );
  AND2X1 U162 ( .IN1(n596), .IN2(n597), .Q(n594) );
  NAND2X0 U163 ( .IN1(P2_N392), .IN2(n598), .QN(n597) );
  NAND2X0 U164 ( .IN1(P2_N4838), .IN2(n599), .QN(n596) );
  NAND2X0 U165 ( .IN1(n600), .IN2(n601), .QN(n1831) );
  NAND2X0 U166 ( .IN1(n6589), .IN2(n9353), .QN(n601) );
  AND2X1 U167 ( .IN1(n602), .IN2(n603), .Q(n600) );
  NAND2X0 U168 ( .IN1(P2_N391), .IN2(n598), .QN(n603) );
  NAND2X0 U169 ( .IN1(P2_N4837), .IN2(n599), .QN(n602) );
  NAND2X0 U170 ( .IN1(n604), .IN2(n605), .QN(n1833) );
  NAND2X0 U171 ( .IN1(n6589), .IN2(n9357), .QN(n605) );
  AND2X1 U172 ( .IN1(n606), .IN2(n607), .Q(n604) );
  NAND2X0 U173 ( .IN1(P2_N390), .IN2(n598), .QN(n607) );
  NAND2X0 U174 ( .IN1(P2_N4836), .IN2(n599), .QN(n606) );
  NAND2X0 U175 ( .IN1(n608), .IN2(n609), .QN(n1835) );
  NAND2X0 U176 ( .IN1(n6589), .IN2(n9361), .QN(n609) );
  AND2X1 U177 ( .IN1(n610), .IN2(n611), .Q(n608) );
  NAND2X0 U178 ( .IN1(P2_N389), .IN2(n598), .QN(n611) );
  NAND2X0 U179 ( .IN1(P2_N4835), .IN2(n599), .QN(n610) );
  NAND2X0 U180 ( .IN1(n612), .IN2(n613), .QN(n1837) );
  NAND2X0 U181 ( .IN1(n6589), .IN2(n9365), .QN(n613) );
  AND2X1 U182 ( .IN1(n614), .IN2(n615), .Q(n612) );
  NAND2X0 U183 ( .IN1(P2_N388), .IN2(n598), .QN(n615) );
  NAND2X0 U184 ( .IN1(P2_N4834), .IN2(n599), .QN(n614) );
  NAND2X0 U185 ( .IN1(n616), .IN2(n617), .QN(n1839) );
  NAND2X0 U186 ( .IN1(n6589), .IN2(n9369), .QN(n617) );
  AND2X1 U187 ( .IN1(n618), .IN2(n619), .Q(n616) );
  NAND2X0 U188 ( .IN1(P2_N387), .IN2(n598), .QN(n619) );
  NAND2X0 U189 ( .IN1(P2_N4833), .IN2(n599), .QN(n618) );
  NAND2X0 U190 ( .IN1(n620), .IN2(n621), .QN(n1841) );
  NAND2X0 U191 ( .IN1(n6589), .IN2(n9373), .QN(n621) );
  AND2X1 U192 ( .IN1(n622), .IN2(n623), .Q(n620) );
  NAND2X0 U193 ( .IN1(P2_N386), .IN2(n598), .QN(n623) );
  NAND2X0 U194 ( .IN1(P2_N4832), .IN2(n599), .QN(n622) );
  NAND2X0 U195 ( .IN1(n624), .IN2(n625), .QN(n1843) );
  NAND2X0 U196 ( .IN1(n6589), .IN2(n9377), .QN(n625) );
  AND2X1 U197 ( .IN1(n626), .IN2(n627), .Q(n624) );
  NAND2X0 U198 ( .IN1(P2_N385), .IN2(n598), .QN(n627) );
  NAND2X0 U199 ( .IN1(P2_N4831), .IN2(n599), .QN(n626) );
  NAND2X0 U200 ( .IN1(n628), .IN2(n629), .QN(n1845) );
  NAND2X0 U201 ( .IN1(n6589), .IN2(n9381), .QN(n629) );
  AND2X1 U202 ( .IN1(n630), .IN2(n631), .Q(n628) );
  NAND2X0 U203 ( .IN1(P2_N384), .IN2(n598), .QN(n631) );
  NAND2X0 U204 ( .IN1(P2_N4830), .IN2(n599), .QN(n630) );
  NAND2X0 U205 ( .IN1(n632), .IN2(n633), .QN(n1847) );
  NAND2X0 U206 ( .IN1(n6589), .IN2(n9501), .QN(n633) );
  AND2X1 U207 ( .IN1(n634), .IN2(n635), .Q(n632) );
  NAND2X0 U208 ( .IN1(P2_N383), .IN2(n598), .QN(n635) );
  NAND2X0 U209 ( .IN1(P2_N4829), .IN2(n599), .QN(n634) );
  NAND2X0 U210 ( .IN1(n636), .IN2(n637), .QN(n1849) );
  NAND2X0 U211 ( .IN1(n6589), .IN2(n9505), .QN(n637) );
  AND2X1 U212 ( .IN1(n638), .IN2(n639), .Q(n636) );
  NAND2X0 U213 ( .IN1(P2_N382), .IN2(n598), .QN(n639) );
  NAND2X0 U214 ( .IN1(P2_N4828), .IN2(n599), .QN(n638) );
  NAND2X0 U215 ( .IN1(n640), .IN2(n641), .QN(n1851) );
  NAND2X0 U216 ( .IN1(n2166), .IN2(n9509), .QN(n641) );
  AND2X1 U217 ( .IN1(n642), .IN2(n643), .Q(n640) );
  NAND2X0 U218 ( .IN1(P2_N381), .IN2(n598), .QN(n643) );
  NAND2X0 U219 ( .IN1(P2_N4827), .IN2(n599), .QN(n642) );
  NAND2X0 U220 ( .IN1(n644), .IN2(n645), .QN(n1853) );
  NAND2X0 U221 ( .IN1(n2166), .IN2(n9513), .QN(n645) );
  AND2X1 U222 ( .IN1(n646), .IN2(n647), .Q(n644) );
  NAND2X0 U223 ( .IN1(P2_N380), .IN2(n598), .QN(n647) );
  NAND2X0 U224 ( .IN1(P2_N4826), .IN2(n599), .QN(n646) );
  NAND2X0 U225 ( .IN1(n648), .IN2(n649), .QN(n1855) );
  NAND2X0 U226 ( .IN1(n2166), .IN2(n9517), .QN(n649) );
  AND2X1 U227 ( .IN1(n650), .IN2(n651), .Q(n648) );
  NAND2X0 U228 ( .IN1(P2_N379), .IN2(n598), .QN(n651) );
  NAND2X0 U229 ( .IN1(P2_N4825), .IN2(n599), .QN(n650) );
  NAND2X0 U230 ( .IN1(n652), .IN2(n653), .QN(n1857) );
  NAND2X0 U231 ( .IN1(n2166), .IN2(n9521), .QN(n653) );
  AND2X1 U232 ( .IN1(n654), .IN2(n655), .Q(n652) );
  NAND2X0 U233 ( .IN1(P2_N378), .IN2(n598), .QN(n655) );
  NAND2X0 U234 ( .IN1(P2_N4824), .IN2(n599), .QN(n654) );
  NAND2X0 U235 ( .IN1(n656), .IN2(n657), .QN(n1859) );
  NAND2X0 U236 ( .IN1(n2166), .IN2(n9525), .QN(n657) );
  AND2X1 U237 ( .IN1(n658), .IN2(n659), .Q(n656) );
  NAND2X0 U238 ( .IN1(P2_N377), .IN2(n598), .QN(n659) );
  NAND2X0 U239 ( .IN1(P2_N4823), .IN2(n599), .QN(n658) );
  NAND2X0 U240 ( .IN1(n660), .IN2(n661), .QN(n1861) );
  NAND2X0 U241 ( .IN1(n2166), .IN2(n9529), .QN(n661) );
  AND2X1 U242 ( .IN1(n662), .IN2(n663), .Q(n660) );
  NAND2X0 U243 ( .IN1(P2_N376), .IN2(n598), .QN(n663) );
  NAND2X0 U244 ( .IN1(P2_N4822), .IN2(n599), .QN(n662) );
  NAND2X0 U245 ( .IN1(n664), .IN2(n665), .QN(n1863) );
  NAND2X0 U246 ( .IN1(n2166), .IN2(n9533), .QN(n665) );
  NAND2X0 U61 ( .IN1(P1_N383), .IN2(n480), .QN(n517) );
  NAND2X0 U62 ( .IN1(P1_N4957), .IN2(n481), .QN(n516) );
  NAND2X0 U63 ( .IN1(n518), .IN2(n519), .QN(n1618) );
  NAND2X0 U64 ( .IN1(n6583), .IN2(n9851), .QN(n519) );
  AND2X1 U65 ( .IN1(n520), .IN2(n521), .Q(n518) );
  NAND2X0 U66 ( .IN1(P1_N382), .IN2(n480), .QN(n521) );
  NAND2X0 U67 ( .IN1(P1_N4956), .IN2(n481), .QN(n520) );
  NAND2X0 U68 ( .IN1(n522), .IN2(n523), .QN(n1621) );
  NAND2X0 U69 ( .IN1(n6583), .IN2(n9665), .QN(n523) );
  AND2X1 U70 ( .IN1(n524), .IN2(n525), .Q(n522) );
  NAND2X0 U71 ( .IN1(P1_N381), .IN2(n480), .QN(n525) );
  NAND2X0 U72 ( .IN1(P1_N4955), .IN2(n481), .QN(n524) );
  NAND2X0 U73 ( .IN1(n526), .IN2(n527), .QN(n1624) );
  NAND2X0 U74 ( .IN1(n6583), .IN2(n9855), .QN(n527) );
  AND2X1 U75 ( .IN1(n528), .IN2(n529), .Q(n526) );
  NAND2X0 U76 ( .IN1(P1_N380), .IN2(n480), .QN(n529) );
  NAND2X0 U77 ( .IN1(P1_N4954), .IN2(n481), .QN(n528) );
  NAND2X0 U78 ( .IN1(n530), .IN2(n531), .QN(n1627) );
  NAND2X0 U79 ( .IN1(n6583), .IN2(n9669), .QN(n531) );
  AND2X1 U80 ( .IN1(n532), .IN2(n533), .Q(n530) );
  NAND2X0 U81 ( .IN1(P1_N379), .IN2(n480), .QN(n533) );
  NAND2X0 U82 ( .IN1(P1_N4953), .IN2(n481), .QN(n532) );
  NAND2X0 U83 ( .IN1(n534), .IN2(n535), .QN(n1630) );
  NAND2X0 U84 ( .IN1(n6583), .IN2(n9859), .QN(n535) );
  AND2X1 U85 ( .IN1(n536), .IN2(n537), .Q(n534) );
  NAND2X0 U86 ( .IN1(P1_N378), .IN2(n480), .QN(n537) );
  NAND2X0 U87 ( .IN1(P1_N4952), .IN2(n481), .QN(n536) );
  NAND2X0 U88 ( .IN1(n538), .IN2(n539), .QN(n1633) );
  NAND2X0 U89 ( .IN1(n6583), .IN2(n9673), .QN(n539) );
  AND2X1 U90 ( .IN1(n540), .IN2(n541), .Q(n538) );
  NAND2X0 U91 ( .IN1(P1_N377), .IN2(n480), .QN(n541) );
  NAND2X0 U92 ( .IN1(P1_N4951), .IN2(n481), .QN(n540) );
  NAND2X0 U93 ( .IN1(n542), .IN2(n543), .QN(n1636) );
  NAND2X0 U94 ( .IN1(n6583), .IN2(n9863), .QN(n543) );
  AND2X1 U95 ( .IN1(n544), .IN2(n545), .Q(n542) );
  NAND2X0 U96 ( .IN1(P1_N376), .IN2(n480), .QN(n545) );
  NAND2X0 U97 ( .IN1(P1_N4950), .IN2(n481), .QN(n544) );
  NAND2X0 U98 ( .IN1(n546), .IN2(n547), .QN(n1639) );
  NAND2X0 U99 ( .IN1(n6583), .IN2(n9677), .QN(n547) );
  AND2X1 U100 ( .IN1(n548), .IN2(n549), .Q(n546) );
  NAND2X0 U101 ( .IN1(P1_N375), .IN2(n480), .QN(n549) );
  NAND2X0 U102 ( .IN1(P1_N4949), .IN2(n481), .QN(n548) );
  NAND2X0 U103 ( .IN1(n550), .IN2(n551), .QN(n1642) );
  NAND2X0 U104 ( .IN1(n6583), .IN2(n9867), .QN(n551) );
  AND2X1 U105 ( .IN1(n552), .IN2(n553), .Q(n550) );
  NAND2X0 U106 ( .IN1(P1_N374), .IN2(n480), .QN(n553) );
  NAND2X0 U107 ( .IN1(P1_N4948), .IN2(n481), .QN(n552) );
  NAND2X0 U108 ( .IN1(n554), .IN2(n555), .QN(n1645) );
  NAND2X0 U109 ( .IN1(n6583), .IN2(n9681), .QN(n555) );
  AND2X1 U110 ( .IN1(n556), .IN2(n557), .Q(n554) );
  NAND2X0 U111 ( .IN1(P1_N373), .IN2(n480), .QN(n557) );
  NAND2X0 U112 ( .IN1(P1_N4947), .IN2(n481), .QN(n556) );
  NAND2X0 U113 ( .IN1(n558), .IN2(n559), .QN(n1648) );
  NAND2X0 U114 ( .IN1(n6583), .IN2(n10011), .QN(n559) );
  AND2X1 U115 ( .IN1(n560), .IN2(n561), .Q(n558) );
  NAND2X0 U116 ( .IN1(P1_N372), .IN2(n480), .QN(n561) );
  NAND2X0 U117 ( .IN1(P1_N4946), .IN2(n481), .QN(n560) );
  NAND2X0 U118 ( .IN1(n562), .IN2(n563), .QN(n1651) );
  NAND2X0 U119 ( .IN1(n6583), .IN2(n9685), .QN(n563) );
  AND2X1 U120 ( .IN1(n564), .IN2(n565), .Q(n562) );
  NAND2X0 U121 ( .IN1(P1_N371), .IN2(n480), .QN(n565) );
  NAND2X0 U122 ( .IN1(P1_N4945), .IN2(n481), .QN(n564) );
  NAND2X0 U123 ( .IN1(n566), .IN2(n567), .QN(n1654) );
  NAND2X0 U124 ( .IN1(n6580), .IN2(n10015), .QN(n567) );
  AND2X1 U125 ( .IN1(n568), .IN2(n569), .Q(n566) );
  NAND2X0 U126 ( .IN1(P1_N370), .IN2(n480), .QN(n569) );
  NAND2X0 U127 ( .IN1(P1_N4944), .IN2(n481), .QN(n568) );
  NAND2X0 U128 ( .IN1(n570), .IN2(n571), .QN(n1657) );
  NAND2X0 U129 ( .IN1(n6580), .IN2(n9689), .QN(n571) );
  AND2X1 U130 ( .IN1(n572), .IN2(n573), .Q(n570) );
  NAND2X0 U131 ( .IN1(P1_N369), .IN2(n480), .QN(n573) );
  NAND2X0 U132 ( .IN1(P1_N4943), .IN2(n481), .QN(n572) );
  NAND2X0 U133 ( .IN1(n574), .IN2(n575), .QN(n1660) );
  NAND2X0 U134 ( .IN1(n6580), .IN2(n9657), .QN(n575) );
  AND2X1 U135 ( .IN1(n576), .IN2(n577), .Q(n574) );
  NAND2X0 U136 ( .IN1(P1_N368), .IN2(n480), .QN(n577) );
  NAND2X0 U137 ( .IN1(P1_N4942), .IN2(n481), .QN(n576) );
  NAND2X0 U138 ( .IN1(n578), .IN2(n579), .QN(n1663) );
  NAND2X0 U139 ( .IN1(n6580), .IN2(n6594), .QN(n579) );
  AND2X1 U140 ( .IN1(n580), .IN2(n581), .Q(n578) );
  NAND2X0 U141 ( .IN1(n18451), .IN2(n480), .QN(n581) );
  NAND2X0 U142 ( .IN1(P1_N4941), .IN2(n481), .QN(n580) );
  NAND2X0 U143 ( .IN1(n582), .IN2(n583), .QN(n1666) );
  NAND2X0 U144 ( .IN1(n6580), .IN2(n6623), .QN(n583) );
  AND2X1 U145 ( .IN1(n584), .IN2(n585), .Q(n582) );
  NAND2X0 U146 ( .IN1(n6623), .IN2(n480), .QN(n585) );
  NAND2X0 U147 ( .IN1(P1_N4940), .IN2(n481), .QN(n584) );
  NAND2X0 U148 ( .IN1(n586), .IN2(n587), .QN(n1669) );
  NAND2X0 U149 ( .IN1(n6580), .IN2(n6622), .QN(n587) );
  AND2X1 U150 ( .IN1(n588), .IN2(n589), .Q(n586) );
  NAND2X0 U151 ( .IN1(n6622), .IN2(n480), .QN(n589) );
  NAND2X0 U152 ( .IN1(P1_N4939), .IN2(n481), .QN(n588) );
  NAND2X0 U153 ( .IN1(n590), .IN2(n591), .QN(n1673) );
  SDFFARX1 P1_addr_reg_7_ ( .QN(n18268), .CLK(clock_G1B2I27_1), .RSTB(n7545), 
        .SE(n7553), .SI(n18269), .D(n6012) );
  SDFFARX1 P1_addr_reg_8_ ( .QN(n18266), .CLK(clock_G1B2I27_1), .RSTB(n7546), 
        .SE(n7553), .SI(n18267), .D(n6011) );
  SDFFARX1 P1_addr_reg_9_ ( .QN(n18186), .CLK(clock_G1B2I27_1), .RSTB(n7546), 
        .SE(n7553), .SI(n18265), .D(n6010), .Q(Scan_Out) );
  SDFFARX1 P1_addr_reg_10_ ( .QN(n18264), .CLK(clock_G1B2I23_1), .RSTB(n6564), 
        .SE(n6576), .SI(test_si2), .D(n6009) );
  SDFFARX1 P1_addr_reg_11_ ( .QN(n18262), .CLK(clock_G1B2I10_1), .RSTB(n7534), 
        .SE(n7536), .SI(n18263), .D(n6008) );
  SDFFARX1 P1_addr_reg_12_ ( .QN(n18260), .CLK(clock_G1B2I10_1), .RSTB(n7532), 
        .SE(n7536), .SI(n18261), .D(n6007) );
  SDFFARX1 P1_addr_reg_13_ ( .QN(n18258), .CLK(clock_G1B2I10_1), .RSTB(n7532), 
        .SE(n7535), .SI(n18259), .D(n6006) );
  SDFFARX1 P1_addr_reg_14_ ( .QN(n18256), .CLK(clock_G1B2I10_1), .RSTB(n7533), 
        .SE(n7535), .SI(n18257), .D(n6005) );
  SDFFARX1 P1_addr_reg_15_ ( .QN(n18254), .CLK(clock_G1B2I10_1), .RSTB(n7533), 
        .SE(n7535), .SI(n18255), .D(n6004) );
  SDFFARX1 P1_addr_reg_16_ ( .QN(n18252), .CLK(clock_G1B2I10_1), .RSTB(n7533), 
        .SE(n7536), .SI(n18253), .D(n6003) );
  SDFFARX1 P1_addr_reg_17_ ( .QN(n18250), .CLK(clock_G1B2I10_1), .RSTB(n7531), 
        .SE(n7536), .SI(n18251), .D(n6002) );
  SDFFARX1 P1_addr_reg_18_ ( .QN(n18248), .CLK(clock_G1B2I10_1), .RSTB(n6564), 
        .SE(n6576), .SI(n18249), .D(n6001) );
  SDFFARX1 P1_addr_reg_19_ ( .QN(n18246), .CLK(clock_G1B2I10_1), .RSTB(n7534), 
        .SE(n7536), .SI(n18247), .D(n6000) );
  SDFFARX1 P2_addr_reg_1_ ( .QN(n18244), .CLK(clock_G1B2I26_1), .RSTB(n7544), 
        .SE(n7452), .SI(n19002), .D(n6196) );
  SDFFARX1 P2_addr_reg_2_ ( .QN(n18242), .CLK(clock_G1B2I26_1), .RSTB(n7544), 
        .SE(n7452), .SI(n18243), .D(n6195) );
  SDFFARX1 P2_addr_reg_3_ ( .QN(n18240), .CLK(clock_G1B2I26_1), .RSTB(n7543), 
        .SE(n7452), .SI(n18241), .D(n6194) );
  SDFFARX1 P2_addr_reg_4_ ( .QN(n18238), .CLK(clock_G1B2I26_1), .RSTB(n7543), 
        .SE(n7452), .SI(n18239), .D(n6193) );
  SDFFARX1 P2_addr_reg_5_ ( .QN(n18236), .CLK(clock_G1B2I26_1), .RSTB(n7542), 
        .SE(n7554), .SI(n18237), .D(n6192) );
  SDFFARX1 P2_addr_reg_6_ ( .QN(n18234), .CLK(clock_G1B2I26_1), .RSTB(n7543), 
        .SE(n7554), .SI(n18235), .D(n6191) );
  SDFFARX1 P2_addr_reg_7_ ( .QN(n18232), .CLK(clock_G1B2I26_1), .RSTB(n7542), 
        .SE(n7552), .SI(n18233), .D(n6190) );
  SDFFARX1 P2_addr_reg_8_ ( .QN(n18230), .CLK(clock_G1B2I3_1), .RSTB(n7542), 
        .SE(n7555), .SI(n18231), .D(n6189) );
  SDFFARX1 P2_addr_reg_9_ ( .QN(n18185), .CLK(clock_G1B2I3_1), .RSTB(n7541), 
        .SE(n7555), .SI(n18229), .D(n6188), .Q(test_so6) );
  SDFFARX1 P2_addr_reg_10_ ( .QN(n18228), .CLK(clock_G1B2I3_1), .RSTB(n7541), 
        .SE(n7555), .SI(test_si7), .D(n6187) );
  SDFFARX1 P2_addr_reg_11_ ( .QN(n18226), .CLK(clock_G1B2I3_1), .RSTB(n7542), 
        .SE(n7554), .SI(n18227), .D(n6186) );
  SDFFARX1 P2_addr_reg_12_ ( .QN(n18224), .CLK(clock_G1B2I26_1), .RSTB(n7543), 
        .SE(n7549), .SI(n18225), .D(n6185) );
  SDFFARX1 P2_addr_reg_13_ ( .QN(n18222), .CLK(clock_G1B2I27_1), .RSTB(n7544), 
        .SE(n7549), .SI(n18223), .D(n6184) );
  SDFFARX1 P2_addr_reg_14_ ( .QN(n18220), .CLK(clock_G1B2I27_1), .RSTB(n7544), 
        .SE(n7549), .SI(n18221), .D(n6183) );
  SDFFARX1 P2_addr_reg_15_ ( .QN(n18218), .CLK(clock_G1B2I27_1), .RSTB(n7543), 
        .SE(n7553), .SI(n18219), .D(n6182) );
  SDFFARX1 P2_addr_reg_16_ ( .QN(n18216), .CLK(clock_G1B2I26_1), .RSTB(n7542), 
        .SE(n7554), .SI(n18217), .D(n6181) );
  SDFFARX1 P2_addr_reg_17_ ( .QN(n18214), .CLK(clock_G1B2I26_1), .RSTB(n7542), 
        .SE(n7552), .SI(n18215), .D(n6180) );
  SDFFARX1 P2_addr_reg_18_ ( .QN(n18212), .CLK(clock_G1B2I26_1), .RSTB(n7543), 
        .SE(n7554), .SI(n18213), .D(n6179) );
  SDFFARX1 P2_addr_reg_19_ ( .QN(n18210), .CLK(clock_G1B2I26_1), .RSTB(n7544), 
        .SE(n7452), .SI(n18211), .D(n6178) );
  SDFFARX1 P2_B_reg ( .QN(P2_N506), .CLK(clock_G1B2I25_1), .RSTB(n7501), 
        .SE(n6573), .SI(test_si6), .D(n6147) );
  SDFFARX1 P2_d_reg_1_ ( .QN(n18207), .CLK(clock_G1B2I25_1), .RSTB(n7501), 
        .SE(n6573), .SI(n6593), .D(n6145) );
  SDFFARX1 P2_d_reg_0_ ( .QN(n18205), .CLK(clock_G1B2I25_1), .RSTB(n7501), 
        .SE(n6573), .SI(n18209), .D(n6146) );
  SDFFARX1 P2_reg1_reg_30_ ( .QN(n18203), .CLK(clock_G1B2I6_1), .RSTB(n7605), 
        .SE(n7496), .SI(n18884), .D(n5958) );
  SDFFARX1 P2_reg0_reg_30_ ( .QN(n18201), .CLK(clock_G1B2I6_1), .RSTB(n7604), 
        .SE(n7450), .SI(n18822), .D(n5957) );
  SDFFARX1 P2_reg2_reg_30_ ( .QN(n18199), .CLK(clock_G1B2I6_1), .RSTB(n7605), 
        .SE(n7495), .SI(n18942), .D(n5954) );
  NOR2X0 U3 ( .QN(wr), .IN1(n470), .IN2(n471) );
  NOR2X0 U6 ( .QN(n471), .IN1(n9325), .IN2(n18189) );
  AND2X1 U7 ( .IN1(n18189), .IN2(n9325), .Q(n470) );
  NOR2X0 U9 ( .QN(rd), .IN1(n473), .IN2(n474) );
  NOR2X0 U10 ( .QN(n474), .IN1(n9322), .IN2(N71) );
  AND2X1 U11 ( .IN1(N71), .IN2(n9322), .Q(n473) );
  NAND2X0 U13 ( .IN1(n476), .IN2(n477), .QN(n1559) );
  NAND2X0 U14 ( .IN1(n6580), .IN2(n9633), .QN(n477) );
  AND2X1 U15 ( .IN1(n478), .IN2(n479), .Q(n476) );
  NAND2X0 U16 ( .IN1(P1_N392), .IN2(n480), .QN(n479) );
  NAND2X0 U17 ( .IN1(P1_N4966), .IN2(n481), .QN(n478) );
  NAND2X0 U18 ( .IN1(n482), .IN2(n483), .QN(n1591) );
  NAND2X0 U19 ( .IN1(n6580), .IN2(n9401), .QN(n483) );
  AND2X1 U20 ( .IN1(n484), .IN2(n485), .Q(n482) );
  NAND2X0 U21 ( .IN1(P1_N391), .IN2(n480), .QN(n485) );
  NAND2X0 U22 ( .IN1(P1_N4965), .IN2(n481), .QN(n484) );
  NAND2X0 U23 ( .IN1(n486), .IN2(n487), .QN(n1594) );
  NAND2X0 U24 ( .IN1(n6580), .IN2(n9637), .QN(n487) );
  AND2X1 U25 ( .IN1(n488), .IN2(n489), .Q(n486) );
  NAND2X0 U26 ( .IN1(P1_N390), .IN2(n480), .QN(n489) );
  NAND2X0 U27 ( .IN1(P1_N4964), .IN2(n481), .QN(n488) );
  NAND2X0 U28 ( .IN1(n490), .IN2(n491), .QN(n1597) );
  NAND2X0 U29 ( .IN1(n6580), .IN2(n9405), .QN(n491) );
  AND2X1 U30 ( .IN1(n492), .IN2(n493), .Q(n490) );
  NAND2X0 U31 ( .IN1(P1_N389), .IN2(n480), .QN(n493) );
  NAND2X0 U32 ( .IN1(P1_N4963), .IN2(n481), .QN(n492) );
  NAND2X0 U33 ( .IN1(n494), .IN2(n495), .QN(n1600) );
  NAND2X0 U34 ( .IN1(n6580), .IN2(n9641), .QN(n495) );
  AND2X1 U35 ( .IN1(n496), .IN2(n497), .Q(n494) );
  NAND2X0 U36 ( .IN1(P1_N388), .IN2(n480), .QN(n497) );
  NAND2X0 U37 ( .IN1(P1_N4962), .IN2(n481), .QN(n496) );
  NAND2X0 U38 ( .IN1(n498), .IN2(n499), .QN(n1603) );
  NAND2X0 U39 ( .IN1(n6580), .IN2(n9409), .QN(n499) );
  AND2X1 U40 ( .IN1(n500), .IN2(n501), .Q(n498) );
  NAND2X0 U41 ( .IN1(P1_N387), .IN2(n480), .QN(n501) );
  NAND2X0 U42 ( .IN1(P1_N4961), .IN2(n481), .QN(n500) );
  NAND2X0 U43 ( .IN1(n502), .IN2(n503), .QN(n1606) );
  NAND2X0 U44 ( .IN1(n6580), .IN2(n9645), .QN(n503) );
  AND2X1 U45 ( .IN1(n504), .IN2(n505), .Q(n502) );
  NAND2X0 U46 ( .IN1(P1_N386), .IN2(n480), .QN(n505) );
  NAND2X0 U47 ( .IN1(P1_N4960), .IN2(n481), .QN(n504) );
  NAND2X0 U48 ( .IN1(n506), .IN2(n507), .QN(n1609) );
  NAND2X0 U49 ( .IN1(n6580), .IN2(n9413), .QN(n507) );
  AND2X1 U50 ( .IN1(n508), .IN2(n509), .Q(n506) );
  NAND2X0 U51 ( .IN1(P1_N385), .IN2(n480), .QN(n509) );
  NAND2X0 U52 ( .IN1(P1_N4959), .IN2(n481), .QN(n508) );
  NAND2X0 U53 ( .IN1(n510), .IN2(n511), .QN(n1612) );
  NAND2X0 U54 ( .IN1(n6580), .IN2(n9649), .QN(n511) );
  AND2X1 U55 ( .IN1(n512), .IN2(n513), .Q(n510) );
  NAND2X0 U56 ( .IN1(P1_N384), .IN2(n480), .QN(n513) );
  NAND2X0 U57 ( .IN1(P1_N4958), .IN2(n481), .QN(n512) );
  NAND2X0 U58 ( .IN1(n514), .IN2(n515), .QN(n1615) );
  NAND2X0 U59 ( .IN1(n6583), .IN2(n9661), .QN(n515) );
  AND2X1 U60 ( .IN1(n516), .IN2(n517), .Q(n514) );
  SDFFARX1 P1_reg3_reg_3_ ( .QN(n18451), .CLK(clock_G1B2I2_1), .RSTB(n7575), 
        .SE(n7584), .SI(n6623), .D(n1663) );
  SDFFARX1 P1_datao_reg_4_ ( .QN(n18449), .CLK(clock_G1B2I30_1), .RSTB(n7590), 
        .SE(n7573), .SI(n18452), .D(n5995) );
  SDFFARX1 P1_reg3_reg_4_ ( .QN(n18447), .CLK(clock_G1B2I28_1), .RSTB(n7532), 
        .SE(n7530), .SI(n6594), .D(n1660) );
  SDFFARX1 P1_datao_reg_5_ ( .QN(n18445), .CLK(clock_G1B2I35_1), .RSTB(n7593), 
        .SE(n7598), .SI(n18448), .D(n5994) );
  SDFFARX1 P1_reg3_reg_5_ ( .QN(n18443), .CLK(clock_G1B2I10_1), .RSTB(n7532), 
        .SE(n7530), .SI(n18446), .D(n1657) );
  SDFFARX1 P1_datao_reg_6_ ( .QN(n18441), .CLK(clock_G1B2I35_1), .RSTB(n7593), 
        .SE(n7598), .SI(n18444), .D(n5993) );
  SDFFARX1 P1_reg3_reg_6_ ( .QN(n18439), .CLK(clock_G1B2I10_1), .RSTB(n6564), 
        .SE(n6576), .SI(n18442), .D(n1654) );
  SDFFARX1 P1_datao_reg_7_ ( .QN(n18437), .CLK(clock_G1B2I35_1), .RSTB(n7593), 
        .SE(n7598), .SI(n18440), .D(n5992) );
  SDFFARX1 P1_reg3_reg_7_ ( .QN(n18435), .CLK(clock_G1B2I23_1), .RSTB(n6564), 
        .SE(n7518), .SI(n18438), .D(n1651) );
  SDFFARX1 P1_datao_reg_8_ ( .QN(n18433), .CLK(clock_G1B2I35_1), .RSTB(n7593), 
        .SE(n7598), .SI(n18436), .D(n5991) );
  SDFFARX1 P1_reg3_reg_8_ ( .QN(n18431), .CLK(clock_G1B2I23_1), .RSTB(n7531), 
        .SE(n7530), .SI(n18434), .D(n1648) );
  SDFFARX1 P1_datao_reg_9_ ( .QN(n18429), .CLK(clock_G1B2I35_1), .RSTB(n7593), 
        .SE(n7598), .SI(n18432), .D(n5990) );
  SDFFARX1 P1_reg3_reg_9_ ( .QN(n18427), .CLK(clock_G1B2I29_1), .RSTB(n7507), 
        .SE(n7517), .SI(n18430), .D(n1645) );
  SDFFARX1 P1_datao_reg_10_ ( .QN(n18425), .CLK(clock_G1B2I35_1), .RSTB(n6560), 
        .SE(n7467), .SI(n18428), .D(n5989) );
  SDFFARX1 P1_reg3_reg_10_ ( .QN(n18423), .CLK(clock_G1B2I29_1), .RSTB(n7508), 
        .SE(n7451), .SI(n18426), .D(n1642) );
  SDFFARX1 P1_datao_reg_11_ ( .QN(n18421), .CLK(clock_G1B2I19_1), .RSTB(n7502), 
        .SE(n7465), .SI(n18424), .D(n5988) );
  SDFFARX1 P1_reg3_reg_11_ ( .QN(n18419), .CLK(clock_G1B2I29_1), .RSTB(n7508), 
        .SE(n7451), .SI(n18422), .D(n1639) );
  SDFFARX1 P1_datao_reg_12_ ( .QN(n18417), .CLK(clock_G1B2I19_1), .RSTB(n7537), 
        .SE(n7467), .SI(n18420), .D(n5987) );
  SDFFARX1 P1_reg3_reg_12_ ( .QN(n18415), .CLK(clock_G1B2I29_1), .RSTB(n7508), 
        .SE(n7451), .SI(n18418), .D(n1636) );
  SDFFARX1 P1_datao_reg_13_ ( .QN(n18413), .CLK(clock_G1B2I19_1), .RSTB(n7537), 
        .SE(n7467), .SI(n18416), .D(n5986) );
  SDFFARX1 P1_reg3_reg_13_ ( .QN(n18411), .CLK(clock_G1B2I29_1), .RSTB(n7507), 
        .SE(n7516), .SI(n18414), .D(n1633) );
  SDFFARX1 P1_datao_reg_14_ ( .QN(n18409), .CLK(clock_G1B2I19_1), .RSTB(n7537), 
        .SE(n7467), .SI(n18412), .D(n5985) );
  SDFFARX1 P1_reg3_reg_14_ ( .QN(n18407), .CLK(clock_G1B2I37_1), .RSTB(n7507), 
        .SE(n7516), .SI(n18410), .D(n1630) );
  SDFFARX1 P1_datao_reg_15_ ( .QN(n18405), .CLK(clock_G1B2I19_1), .RSTB(n7524), 
        .SE(n7465), .SI(n18408), .D(n5984) );
  SDFFARX1 P1_reg3_reg_15_ ( .QN(n18403), .CLK(clock_G1B2I37_1), .RSTB(n7509), 
        .SE(n7516), .SI(n18406), .D(n1627) );
  SDFFARX1 P1_datao_reg_16_ ( .QN(n18401), .CLK(clock_G1B2I35_1), .RSTB(n7524), 
        .SE(n7467), .SI(n18404), .D(n5983) );
  SDFFARX1 P1_reg3_reg_16_ ( .QN(n18399), .CLK(clock_G1B2I37_1), .RSTB(n7523), 
        .SE(n7528), .SI(n18402), .D(n1624) );
  SDFFARX1 P1_datao_reg_17_ ( .QN(n18397), .CLK(clock_G1B2I35_1), .RSTB(n7593), 
        .SE(n7598), .SI(n18400), .D(n5982) );
  SDFFARX1 P1_reg3_reg_17_ ( .QN(n18395), .CLK(clock_G1B2I31_1), .RSTB(n7523), 
        .SE(n7527), .SI(n18398), .D(n1621) );
  SDFFARX1 P1_datao_reg_18_ ( .QN(n18393), .CLK(clock_G1B2I30_1), .RSTB(n7592), 
        .SE(n7573), .SI(n18396), .D(n5981) );
  SDFFARX1 P1_reg3_reg_18_ ( .QN(n18391), .CLK(clock_G1B2I31_1), .RSTB(n7523), 
        .SE(n7526), .SI(n18394), .D(n1618) );
  SDFFARX1 P1_datao_reg_19_ ( .QN(n18389), .CLK(clock_G1B2I30_1), .RSTB(n7590), 
        .SE(n7573), .SI(n18392), .D(n5980) );
  SDFFARX1 P1_reg3_reg_19_ ( .QN(n18387), .CLK(clock_G1B2I31_1), .RSTB(n7523), 
        .SE(n7526), .SI(n18390), .D(n1615) );
  SDFFARX1 P1_datao_reg_20_ ( .QN(n18385), .CLK(clock_G1B2I22_1), .RSTB(n7545), 
        .SE(n6574), .SI(n18388), .D(n5979) );
  SDFFARX1 P1_reg3_reg_20_ ( .QN(n18383), .CLK(clock_G1B2I11_1), .RSTB(n7476), 
        .SE(n6578), .SI(n18386), .D(n1612) );
  SDFFARX1 P1_datao_reg_21_ ( .QN(n18381), .CLK(clock_G1B2I22_1), .RSTB(n7546), 
        .SE(n6574), .SI(n18384), .D(n5978) );
  SDFFARX1 P1_reg3_reg_21_ ( .QN(n18379), .CLK(clock_G1B2I11_1), .RSTB(n7476), 
        .SE(n6578), .SI(n18382), .D(n1609) );
  SDFFARX1 P1_datao_reg_22_ ( .QN(n18377), .CLK(clock_G1B2I22_1), .RSTB(n7548), 
        .SE(n7549), .SI(n18380), .D(n5977) );
  SDFFARX1 P1_reg3_reg_22_ ( .QN(n18375), .CLK(clock_G1B2I11_1), .RSTB(n6566), 
        .SE(n6575), .SI(n18378), .D(n1606) );
  SDFFARX1 P1_datao_reg_23_ ( .QN(n18373), .CLK(clock_G1B2I24_1), .RSTB(n7606), 
        .SE(n7489), .SI(n18376), .D(n5976) );
  SDFFARX1 P1_reg3_reg_23_ ( .QN(n18371), .CLK(clock_G1B2I20_1), .RSTB(n6566), 
        .SE(n7478), .SI(n18374), .D(n1603) );
  SDFFARX1 P1_datao_reg_24_ ( .QN(n18369), .CLK(clock_G1B2I24_1), .RSTB(n7606), 
        .SE(n7489), .SI(n18372), .D(n5975) );
  SDFFARX1 P1_reg3_reg_24_ ( .QN(n18367), .CLK(clock_G1B2I1_1), .RSTB(n7576), 
        .SE(n7585), .SI(n18370), .D(n1600) );
  SDFFARX1 P1_datao_reg_25_ ( .QN(n18365), .CLK(clock_G1B2I24_1), .RSTB(n7606), 
        .SE(n7490), .SI(n18368), .D(n5974) );
  SDFFARX1 P1_reg3_reg_25_ ( .QN(n18363), .CLK(clock_G1B2I1_1), .RSTB(n7576), 
        .SE(n7586), .SI(n18366), .D(n1597) );
  SDFFARX1 P1_datao_reg_26_ ( .QN(n18361), .CLK(clock_G1B2I24_1), .RSTB(n7594), 
        .SE(n7490), .SI(n18364), .D(n5973) );
  SDFFARX1 P1_reg3_reg_26_ ( .QN(n18359), .CLK(clock_G1B2I1_1), .RSTB(n7576), 
        .SE(n7586), .SI(n18362), .D(n1594) );
  SDFFARX1 P1_datao_reg_27_ ( .QN(n18357), .CLK(clock_G1B2I24_1), .RSTB(n7594), 
        .SE(n7490), .SI(n18360), .D(n5972) );
  SDFFARX1 P1_reg3_reg_27_ ( .QN(n18355), .CLK(clock_G1B2I1_1), .RSTB(n7576), 
        .SE(n7586), .SI(n18358), .D(n1591) );
  SDFFARX1 P1_datao_reg_28_ ( .QN(n18353), .CLK(clock_G1B2I24_1), .RSTB(n7606), 
        .SE(n7489), .SI(n18356), .D(n5971) );
  SDFFARX1 P2_IR_reg_28_ ( .QN(n18351), .CLK(clock_G1B2I3_1), .RSTB(n6562), 
        .SE(n7555), .SI(n18348), .D(n6198) );
  SDFFARX1 P2_IR_reg_27_ ( .QN(n18349), .CLK(clock_G1B2I3_1), .RSTB(n6562), 
        .SE(n7556), .SI(n18320), .D(n6199) );
  SDFFARX1 P2_IR_reg_0_ ( .QN(n18347), .CLK(clock_G1B2I13_1), .RSTB(n7589), 
        .SE(n7599), .SI(n6591), .D(n6316) );
  SDFFARX1 P2_IR_reg_1_ ( .QN(n18345), .CLK(clock_G1B2I13_1), .RSTB(n7589), 
        .SE(n7600), .SI(n6595), .D(n6315) );
  SDFFARX1 P2_IR_reg_2_ ( .QN(n18343), .CLK(clock_G1B2I13_1), .RSTB(n7591), 
        .SE(n7600), .SI(n6596), .D(n6314) );
  SDFFARX1 P2_IR_reg_3_ ( .QN(n18341), .CLK(clock_G1B2I14_1), .RSTB(n6565), 
        .SE(n7596), .SI(n6597), .D(n6313) );
  SDFFARX1 P2_IR_reg_4_ ( .QN(n18339), .CLK(clock_G1B2I19_1), .RSTB(n7537), 
        .SE(n7467), .SI(n6598), .D(n6312) );
  SDFFARX1 P2_IR_reg_5_ ( .QN(n18337), .CLK(clock_G1B2I19_1), .RSTB(n7537), 
        .SE(n7466), .SI(n6599), .D(n6311) );
  SDFFARX1 P2_IR_reg_6_ ( .QN(n18335), .CLK(clock_G1B2I19_1), .RSTB(n7537), 
        .SE(n7466), .SI(n6600), .D(n6310) );
  SDFFARX1 P2_IR_reg_7_ ( .QN(n18333), .CLK(clock_G1B2I19_1), .RSTB(n6560), 
        .SE(n7466), .SI(n6601), .D(n6309) );
  SDFFARX1 P2_IR_reg_8_ ( .QN(n18331), .CLK(clock_G1B2I19_1), .RSTB(n7524), 
        .SE(n7466), .SI(n6602), .D(n6308) );
  SDFFARX1 P2_IR_reg_9_ ( .QN(n18329), .CLK(clock_G1B2I18_1), .RSTB(n7534), 
        .SE(n7466), .SI(n6603), .D(n6307) );
  SDFFARX1 P2_IR_reg_10_ ( .QN(n18327), .CLK(clock_G1B2I18_1), .RSTB(n7538), 
        .SE(n6572), .SI(n6604), .D(n6306) );
  SDFFARX1 P2_IR_reg_11_ ( .QN(n18325), .CLK(clock_G1B2I18_1), .RSTB(n7538), 
        .SE(n7464), .SI(n6605), .D(n6305) );
  SDFFARX1 P2_IR_reg_12_ ( .QN(n18323), .CLK(clock_G1B2I18_1), .RSTB(n7538), 
        .SE(n7464), .SI(n6606), .D(n6304) );
  SDFFARX1 P2_IR_reg_26_ ( .QN(n18321), .CLK(clock_G1B2I3_1), .RSTB(n7541), 
        .SE(n7556), .SI(n18318), .D(n6290) );
  SDFFARX1 P2_IR_reg_25_ ( .QN(n18319), .CLK(clock_G1B2I3_1), .RSTB(n7541), 
        .SE(n7556), .SI(n18316), .D(n6291) );
  SDFFARX1 P2_IR_reg_24_ ( .QN(n18317), .CLK(clock_G1B2I30_1), .RSTB(n7590), 
        .SE(n7550), .SI(n6719), .D(n6292) );
  SDFFARX1 P2_IR_reg_22_ ( .QN(n18315), .CLK(clock_G1B2I30_1), .RSTB(n7592), 
        .SE(Scan_Enable), .SI(n6609), .D(n6294) );
  SDFFARX1 P2_IR_reg_21_ ( .QN(n18313), .CLK(clock_G1B2I13_1), .RSTB(n7591), 
        .SE(n7600), .SI(n6610), .D(n6295) );
  SDFFARX1 P2_IR_reg_20_ ( .QN(n18311), .CLK(clock_G1B2I36_1), .RSTB(n7588), 
        .SE(n7597), .SI(n6611), .D(n6296) );
  SDFFARX1 P2_IR_reg_19_ ( .QN(n18309), .CLK(clock_G1B2I36_1), .RSTB(n7592), 
        .SE(n7597), .SI(n6612), .D(n6297) );
  SDFFARX1 P2_IR_reg_18_ ( .QN(n18307), .CLK(clock_G1B2I14_1), .RSTB(n6565), 
        .SE(n7596), .SI(n6613), .D(n6298) );
  SDFFARX1 P2_IR_reg_17_ ( .QN(n18305), .CLK(clock_G1B2I18_1), .RSTB(n7534), 
        .SE(n7465), .SI(n6614), .D(n6299) );
  SDFFARX1 P2_IR_reg_16_ ( .QN(n18303), .CLK(clock_G1B2I18_1), .RSTB(n7534), 
        .SE(n7465), .SI(n6615), .D(n6300) );
  SDFFARX1 P2_IR_reg_15_ ( .QN(n18301), .CLK(clock_G1B2I18_1), .RSTB(n6560), 
        .SE(n7464), .SI(n6616), .D(n6301) );
  SDFFARX1 P2_IR_reg_14_ ( .QN(n18299), .CLK(clock_G1B2I18_1), .RSTB(n7538), 
        .SE(n7464), .SI(n6617), .D(n6302) );
  SDFFARX1 P2_IR_reg_13_ ( .QN(n18297), .CLK(clock_G1B2I18_1), .RSTB(n7538), 
        .SE(n7464), .SI(n6607), .D(n6303) );
  SDFFARX1 P2_rd_reg ( .QN(N71), .CLK(clock_G1B2I22_1), .RSTB(n7546), 
        .SE(n6574), .SI(n19010), .D(P2_N5440) );
  SDFFARX1 P1_reg3_reg_28_ ( .QN(n18294), .CLK(clock_G1B2I1_1), .RSTB(n7578), 
        .SE(n7582), .SI(n18354), .D(n1559) );
  SDFFARX1 P1_reg2_reg_31_ ( .QN(n18292), .CLK(clock_G1B2I2_1), .RSTB(n7575), 
        .SE(n7581), .SI(n18289), .D(n5959) );
  SDFFARX1 P1_reg2_reg_30_ ( .QN(n18290), .CLK(clock_G1B2I1_1), .RSTB(n7580), 
        .SE(n7583), .SI(n18586), .D(n5960) );
  SDFFARX1 P1_B_reg ( .QN(P1_N506), .CLK(clock_G1B2I11_1), .RSTB(n7476), 
        .SE(n6578), .SI(Scan_In), .D(n5970) );
  SDFFARX1 P1_d_reg_1_ ( .QN(n18287), .CLK(clock_G1B2I2_1), .RSTB(n7580), 
        .SE(n7583), .SI(n6620), .D(n5968) );
  SDFFARX1 P1_d_reg_0_ ( .QN(n18285), .CLK(clock_G1B2I2_1), .RSTB(n7575), 
        .SE(n7584), .SI(n18245), .D(n5969) );
  SDFFARX1 P1_rd_reg ( .QN(N74), .CLK(clock_G1B2I10_1), .RSTB(n6564), 
        .SE(n6576), .SI(n19014), .D(P1_N5518) );
  SDFFARX1 P1_addr_reg_0_ ( .QN(n18282), .CLK(clock_G1B2I27_1), .RSTB(n7533), 
        .SE(n7535), .SI(n6708), .D(n6019) );
  SDFFARX1 P1_addr_reg_1_ ( .QN(n18280), .CLK(clock_G1B2I27_1), .RSTB(n7533), 
        .SE(n7535), .SI(n18281), .D(n6018) );
  SDFFARX1 P1_addr_reg_2_ ( .QN(n18278), .CLK(clock_G1B2I27_1), .RSTB(n7533), 
        .SE(n7535), .SI(n18279), .D(n6017) );
  SDFFARX1 P1_addr_reg_3_ ( .QN(n18276), .CLK(clock_G1B2I27_1), .RSTB(n7545), 
        .SE(n7554), .SI(n18277), .D(n6016) );
  SDFFARX1 P1_addr_reg_4_ ( .QN(n18274), .CLK(clock_G1B2I27_1), .RSTB(n7545), 
        .SE(n7549), .SI(n18275), .D(n6015) );
  SDFFARX1 P1_addr_reg_5_ ( .QN(n18272), .CLK(clock_G1B2I27_1), .RSTB(n7545), 
        .SE(n7553), .SI(n18273), .D(n6014) );
  SDFFARX1 P1_addr_reg_6_ ( .QN(n18270), .CLK(clock_G1B2I27_1), .RSTB(n7545), 
        .SE(n7553), .SI(n18271), .D(n6013) );
  SDFFARX1 P1_reg2_reg_6_ ( .QN(n18631), .CLK(clock_G1B2I23_1), .RSTB(n7531), 
        .SE(n7451), .SI(n18632), .D(n6043) );
  SDFFARX1 P1_reg2_reg_7_ ( .QN(n18629), .CLK(clock_G1B2I23_1), .RSTB(n7509), 
        .SE(n7517), .SI(n18630), .D(n6042) );
  SDFFARX1 P1_reg2_reg_8_ ( .QN(n18627), .CLK(clock_G1B2I29_1), .RSTB(n7509), 
        .SE(n7517), .SI(n18628), .D(n6041) );
  SDFFARX1 P1_reg2_reg_9_ ( .QN(n18625), .CLK(clock_G1B2I29_1), .RSTB(n7507), 
        .SE(n7516), .SI(n18626), .D(n6040) );
  SDFFARX1 P1_reg2_reg_10_ ( .QN(n18623), .CLK(clock_G1B2I21_1), .RSTB(n7508), 
        .SE(n7515), .SI(n18624), .D(n6039) );
  SDFFARX1 P1_reg2_reg_11_ ( .QN(n18621), .CLK(clock_G1B2I21_1), .RSTB(n7508), 
        .SE(n7515), .SI(n18622), .D(n6038) );
  SDFFARX1 P1_reg2_reg_12_ ( .QN(n18619), .CLK(clock_G1B2I21_1), .RSTB(n7510), 
        .SE(n7514), .SI(n18620), .D(n6037) );
  SDFFARX1 P1_reg2_reg_13_ ( .QN(n18617), .CLK(clock_G1B2I21_1), .RSTB(n7512), 
        .SE(n7514), .SI(n18618), .D(n6036) );
  SDFFARX1 P1_reg2_reg_14_ ( .QN(n18615), .CLK(clock_G1B2I34_1), .RSTB(n7511), 
        .SE(n7513), .SI(n18616), .D(n6035) );
  SDFFARX1 P1_reg2_reg_15_ ( .QN(n18613), .CLK(clock_G1B2I34_1), .RSTB(n7512), 
        .SE(n7513), .SI(n18614), .D(n6034) );
  SDFFARX1 P1_reg2_reg_16_ ( .QN(n18611), .CLK(clock_G1B2I34_1), .RSTB(n7522), 
        .SE(n7525), .SI(n18612), .D(n6033) );
  SDFFARX1 P1_reg2_reg_17_ ( .QN(n18609), .CLK(clock_G1B2I34_1), .RSTB(n7522), 
        .SE(n7525), .SI(n18610), .D(n6032) );
  SDFFARX1 P1_reg2_reg_18_ ( .QN(n18607), .CLK(clock_G1B2I37_1), .RSTB(n7519), 
        .SE(n7527), .SI(n18608), .D(n6031) );
  SDFFARX1 P1_reg2_reg_19_ ( .QN(n18188), .CLK(clock_G1B2I31_1), .RSTB(n7521), 
        .SE(n7527), .SI(n18606), .D(n6030), .Q(test_so4) );
  SDFFARX1 P1_reg2_reg_20_ ( .QN(n18605), .CLK(clock_G1B2I31_1), .RSTB(n7524), 
        .SE(n7526), .SI(test_si5), .D(n6029) );
  SDFFARX1 P1_reg2_reg_21_ ( .QN(n18603), .CLK(clock_G1B2I11_1), .RSTB(n7476), 
        .SE(n7475), .SI(n18604), .D(n6028) );
  SDFFARX1 P1_reg2_reg_22_ ( .QN(n18601), .CLK(clock_G1B2I11_1), .RSTB(n7476), 
        .SE(n7475), .SI(n18602), .D(n6027) );
  SDFFARX1 P1_reg2_reg_23_ ( .QN(n18599), .CLK(clock_G1B2I20_1), .RSTB(n6566), 
        .SE(n7478), .SI(n18600), .D(n6026) );
  SDFFARX1 P1_reg2_reg_24_ ( .QN(n18597), .CLK(clock_G1B2I20_1), .RSTB(n7577), 
        .SE(n7585), .SI(n18598), .D(n6025) );
  SDFFARX1 P1_reg2_reg_25_ ( .QN(n18595), .CLK(clock_G1B2I1_1), .RSTB(n7576), 
        .SE(n7585), .SI(n18596), .D(n6024) );
  SDFFARX1 P1_reg2_reg_26_ ( .QN(n18593), .CLK(clock_G1B2I1_1), .RSTB(n7576), 
        .SE(n7586), .SI(n18594), .D(n6023) );
  SDFFARX1 P1_reg2_reg_27_ ( .QN(n18591), .CLK(clock_G1B2I1_1), .RSTB(n7578), 
        .SE(n7586), .SI(n18592), .D(n6022) );
  SDFFARX1 P1_reg2_reg_28_ ( .QN(n18589), .CLK(clock_G1B2I1_1), .RSTB(n7578), 
        .SE(n7582), .SI(n18590), .D(n6021) );
  SDFFARX1 P1_reg2_reg_29_ ( .QN(n18587), .CLK(clock_G1B2I1_1), .RSTB(n7578), 
        .SE(n7582), .SI(n18588), .D(n6020) );
  SDFFARX1 P1_reg1_reg_0_ ( .QN(n1503), .CLK(clock_G1B2I20_1), .RSTB(n7477), 
        .SE(n7475), .SI(n19016), .D(n6079) );
  SDFFARX1 P1_reg1_reg_1_ ( .QN(n18585), .CLK(clock_G1B2I28_1), .RSTB(n7574), 
        .SE(n6569), .SI(n18194), .D(n6078) );
  SDFFARX1 P1_reg1_reg_2_ ( .QN(n18583), .CLK(clock_G1B2I28_1), .RSTB(n7574), 
        .SE(n6569), .SI(n18584), .D(n6077) );
  SDFFARX1 P1_reg1_reg_3_ ( .QN(n18581), .CLK(clock_G1B2I28_1), .RSTB(n7574), 
        .SE(n7587), .SI(n18582), .D(n6076) );
  SDFFARX1 P1_reg1_reg_4_ ( .QN(n18579), .CLK(clock_G1B2I28_1), .RSTB(n7574), 
        .SE(n7587), .SI(n18580), .D(n6075) );
  SDFFARX1 P1_reg1_reg_5_ ( .QN(n18577), .CLK(clock_G1B2I10_1), .RSTB(n7532), 
        .SE(n7530), .SI(n18578), .D(n6074) );
  SDFFARX1 P1_reg1_reg_6_ ( .QN(n18575), .CLK(clock_G1B2I23_1), .RSTB(n7531), 
        .SE(n7451), .SI(n18576), .D(n6073) );
  SDFFARX1 P1_reg1_reg_7_ ( .QN(n18573), .CLK(clock_G1B2I23_1), .RSTB(n7509), 
        .SE(n7517), .SI(n18574), .D(n6072) );
  SDFFARX1 P1_reg1_reg_8_ ( .QN(n18187), .CLK(clock_G1B2I29_1), .RSTB(n7507), 
        .SE(n7516), .SI(n18572), .D(n6071), .Q(test_so3) );
  SDFFARX1 P1_reg1_reg_9_ ( .QN(n18571), .CLK(clock_G1B2I21_1), .RSTB(n7510), 
        .SE(n7515), .SI(test_si4), .D(n6070) );
  SDFFARX1 P1_reg1_reg_10_ ( .QN(n18569), .CLK(clock_G1B2I21_1), .RSTB(n7510), 
        .SE(n7515), .SI(n18570), .D(n6069) );
  SDFFARX1 P1_reg1_reg_11_ ( .QN(n18567), .CLK(clock_G1B2I21_1), .RSTB(n7510), 
        .SE(n7514), .SI(n18568), .D(n6068) );
  SDFFARX1 P1_reg1_reg_12_ ( .QN(n18565), .CLK(clock_G1B2I21_1), .RSTB(n7510), 
        .SE(n7514), .SI(n18566), .D(n6067) );
  SDFFARX1 P1_reg1_reg_13_ ( .QN(n18563), .CLK(clock_G1B2I21_1), .RSTB(n7511), 
        .SE(n7513), .SI(n18564), .D(n6066) );
  SDFFARX1 P1_reg1_reg_14_ ( .QN(n18561), .CLK(clock_G1B2I34_1), .RSTB(n7511), 
        .SE(n7513), .SI(n18562), .D(n6065) );
  SDFFARX1 P1_reg1_reg_15_ ( .QN(n18559), .CLK(clock_G1B2I34_1), .RSTB(n7522), 
        .SE(n7525), .SI(n18560), .D(n6064) );
  SDFFARX1 P1_reg1_reg_16_ ( .QN(n18557), .CLK(clock_G1B2I34_1), .RSTB(n7522), 
        .SE(n7525), .SI(n18558), .D(n6063) );
  SDFFARX1 P1_reg1_reg_17_ ( .QN(n18555), .CLK(clock_G1B2I37_1), .RSTB(n7522), 
        .SE(n7525), .SI(n18556), .D(n6062) );
  SDFFARX1 P1_reg1_reg_18_ ( .QN(n18553), .CLK(clock_G1B2I31_1), .RSTB(n7519), 
        .SE(n7527), .SI(n18554), .D(n6061) );
  SDFFARX1 P1_reg1_reg_19_ ( .QN(n18551), .CLK(clock_G1B2I31_1), .RSTB(n7521), 
        .SE(n7526), .SI(n18552), .D(n6060) );
  SDFFARX1 P1_reg1_reg_20_ ( .QN(n18549), .CLK(clock_G1B2I31_1), .RSTB(n7523), 
        .SE(n7526), .SI(n18550), .D(n6059) );
  SDFFARX1 P1_reg1_reg_21_ ( .QN(n18547), .CLK(clock_G1B2I11_1), .RSTB(n7477), 
        .SE(n6578), .SI(n18548), .D(n6058) );
  SDFFARX1 P1_reg1_reg_22_ ( .QN(n18545), .CLK(clock_G1B2I11_1), .RSTB(n7477), 
        .SE(n7475), .SI(n18546), .D(n6057) );
  SDFFARX1 P1_reg1_reg_23_ ( .QN(n18543), .CLK(clock_G1B2I20_1), .RSTB(n7477), 
        .SE(n7478), .SI(n18544), .D(n6056) );
  SDFFARX1 P1_reg1_reg_24_ ( .QN(n18541), .CLK(clock_G1B2I20_1), .RSTB(n7471), 
        .SE(n7478), .SI(n18542), .D(n6055) );
  SDFFARX1 P1_reg1_reg_25_ ( .QN(n18539), .CLK(clock_G1B2I20_1), .RSTB(n7579), 
        .SE(n7586), .SI(n18540), .D(n6054) );
  SDFFARX1 P1_reg1_reg_26_ ( .QN(n18537), .CLK(clock_G1B2I20_1), .RSTB(n7577), 
        .SE(n7585), .SI(n18538), .D(n6053) );
  SDFFARX1 P1_reg1_reg_27_ ( .QN(n18535), .CLK(clock_G1B2I1_1), .RSTB(n7577), 
        .SE(n7584), .SI(n18536), .D(n6052) );
  SDFFARX1 P1_reg1_reg_28_ ( .QN(n18533), .CLK(clock_G1B2I2_1), .RSTB(n7579), 
        .SE(n7583), .SI(n18534), .D(n6051) );
  SDFFARX1 P1_reg1_reg_29_ ( .QN(n18531), .CLK(clock_G1B2I2_1), .RSTB(n7579), 
        .SE(n7583), .SI(n18532), .D(n6050) );
  SDFFARX1 P1_reg1_reg_30_ ( .QN(n18529), .CLK(clock_G1B2I2_1), .RSTB(n7579), 
        .SE(n7581), .SI(n18530), .D(n5962) );
  SDFFARX1 P1_reg1_reg_31_ ( .QN(n18527), .CLK(clock_G1B2I20_1), .RSTB(n7575), 
        .SE(n6569), .SI(n18528), .D(n5961) );
  SDFFARX1 P1_reg0_reg_0_ ( .QN(n18525), .CLK(clock_G1B2I28_1), .RSTB(n7574), 
        .SE(n7587), .SI(n18283), .D(n6109) );
  SDFFARX1 P1_reg0_reg_1_ ( .QN(n18523), .CLK(clock_G1B2I2_1), .RSTB(n6557), 
        .SE(n7581), .SI(n18524), .D(n6108) );
  SDFFARX1 P1_reg0_reg_2_ ( .QN(n18521), .CLK(clock_G1B2I2_1), .RSTB(n6557), 
        .SE(n7584), .SI(n18522), .D(n6107) );
  SDFFARX1 P1_reg0_reg_3_ ( .QN(n18519), .CLK(clock_G1B2I28_1), .RSTB(n6557), 
        .SE(n7587), .SI(n18520), .D(n6106) );
  SDFFARX1 P1_reg0_reg_4_ ( .QN(n18517), .CLK(clock_G1B2I28_1), .RSTB(n7532), 
        .SE(n7530), .SI(n18518), .D(n6105) );
  SDFFARX1 P1_reg0_reg_5_ ( .QN(n18515), .CLK(clock_G1B2I10_1), .RSTB(n7531), 
        .SE(n6576), .SI(n18516), .D(n6104) );
  SDFFARX1 P1_reg0_reg_6_ ( .QN(n18513), .CLK(clock_G1B2I10_1), .RSTB(n6564), 
        .SE(n6576), .SI(n18514), .D(n6103) );
  SDFFARX1 P1_reg0_reg_7_ ( .QN(n18511), .CLK(clock_G1B2I23_1), .RSTB(n7509), 
        .SE(n7517), .SI(n18512), .D(n6102) );
  SDFFARX1 P1_reg0_reg_8_ ( .QN(n18509), .CLK(clock_G1B2I23_1), .RSTB(n7509), 
        .SE(n7517), .SI(n18510), .D(n6101) );
  SDFFARX1 P1_reg0_reg_9_ ( .QN(n18507), .CLK(clock_G1B2I29_1), .RSTB(n7507), 
        .SE(n7516), .SI(n18508), .D(n6100) );
  SDFFARX1 P1_reg0_reg_10_ ( .QN(n18505), .CLK(clock_G1B2I29_1), .RSTB(n7508), 
        .SE(n7451), .SI(n18506), .D(n6099) );
  SDFFARX1 P1_reg0_reg_11_ ( .QN(n18503), .CLK(clock_G1B2I21_1), .RSTB(n7510), 
        .SE(n7515), .SI(n18504), .D(n6098) );
  SDFFARX1 P1_reg0_reg_12_ ( .QN(n18501), .CLK(clock_G1B2I21_1), .RSTB(n7512), 
        .SE(n7515), .SI(n18502), .D(n6097) );
  SDFFARX1 P1_reg0_reg_13_ ( .QN(n18499), .CLK(clock_G1B2I21_1), .RSTB(n7512), 
        .SE(n7514), .SI(n18500), .D(n6096) );
  SDFFARX1 P1_reg0_reg_14_ ( .QN(n18497), .CLK(clock_G1B2I21_1), .RSTB(n7511), 
        .SE(n7514), .SI(n18498), .D(n6095) );
  SDFFARX1 P1_reg0_reg_15_ ( .QN(n18495), .CLK(clock_G1B2I34_1), .RSTB(n7511), 
        .SE(n7513), .SI(n18496), .D(n6094) );
  SDFFARX1 P1_reg0_reg_16_ ( .QN(n18493), .CLK(clock_G1B2I34_1), .RSTB(n7511), 
        .SE(n7513), .SI(n18494), .D(n6093) );
  SDFFARX1 P1_reg0_reg_17_ ( .QN(n18491), .CLK(clock_G1B2I37_1), .RSTB(n7522), 
        .SE(n7525), .SI(n18492), .D(n6092) );
  SDFFARX1 P1_reg0_reg_18_ ( .QN(n18489), .CLK(clock_G1B2I37_1), .RSTB(n7521), 
        .SE(n7527), .SI(n18490), .D(n6091) );
  SDFFARX1 P1_reg0_reg_19_ ( .QN(n18487), .CLK(clock_G1B2I31_1), .RSTB(n7521), 
        .SE(n7527), .SI(n18488), .D(n6090) );
  SDFFARX1 P1_reg0_reg_20_ ( .QN(n18485), .CLK(clock_G1B2I31_1), .RSTB(n7523), 
        .SE(n7526), .SI(n18486), .D(n6089) );
  SDFFARX1 P1_reg0_reg_21_ ( .QN(n18483), .CLK(clock_G1B2I11_1), .RSTB(n7476), 
        .SE(n6578), .SI(n18484), .D(n6088) );
  SDFFARX1 P1_reg0_reg_22_ ( .QN(n18481), .CLK(clock_G1B2I11_1), .RSTB(n7477), 
        .SE(n6575), .SI(n18482), .D(n6087) );
  SDFFARX1 P1_reg0_reg_23_ ( .QN(n18479), .CLK(clock_G1B2I20_1), .RSTB(n7477), 
        .SE(n7478), .SI(n18480), .D(n6086) );
  SDFFARX1 P1_reg0_reg_24_ ( .QN(n18477), .CLK(clock_G1B2I20_1), .RSTB(n7471), 
        .SE(n7478), .SI(n18478), .D(n6085) );
  SDFFARX1 P1_reg0_reg_25_ ( .QN(n18475), .CLK(clock_G1B2I20_1), .RSTB(n7577), 
        .SE(n7585), .SI(n18476), .D(n6084) );
  SDFFARX1 P1_reg0_reg_26_ ( .QN(n18473), .CLK(clock_G1B2I1_1), .RSTB(n7577), 
        .SE(n7585), .SI(n18474), .D(n6083) );
  SDFFARX1 P1_reg0_reg_27_ ( .QN(n18471), .CLK(clock_G1B2I1_1), .RSTB(n7577), 
        .SE(n7584), .SI(n18472), .D(n6082) );
  SDFFARX1 P1_reg0_reg_28_ ( .QN(n18469), .CLK(clock_G1B2I1_1), .RSTB(n7578), 
        .SE(n7583), .SI(n18470), .D(n6081) );
  SDFFARX1 P1_reg0_reg_29_ ( .QN(n18467), .CLK(clock_G1B2I1_1), .RSTB(n7578), 
        .SE(n7582), .SI(n18468), .D(n6080) );
  SDFFARX1 P1_reg3_reg_0_ ( .QN(n18465), .CLK(clock_G1B2I2_1), .RSTB(n7580), 
        .SE(n7584), .SI(n18291), .D(n1673) );
  SDFFARX1 P1_datao_reg_0_ ( .QN(n18463), .CLK(clock_G1B2I3_1), .RSTB(n7541), 
        .SE(n7556), .SI(n6619), .D(n5999) );
  SDFFARX1 P1_datao_reg_1_ ( .QN(n18461), .CLK(clock_G1B2I3_1), .RSTB(n6562), 
        .SE(n7556), .SI(n18462), .D(n5998) );
  SDFFARX1 P1_reg3_reg_1_ ( .QN(n18459), .CLK(clock_G1B2I2_1), .RSTB(n7580), 
        .SE(n7582), .SI(n6621), .D(n1669) );
  SDFFARX1 P1_datao_reg_2_ ( .QN(n18457), .CLK(clock_G1B2I3_1), .RSTB(n6562), 
        .SE(n7555), .SI(n18460), .D(n5997) );
  SDFFARX1 P1_reg3_reg_2_ ( .QN(n18455), .CLK(clock_G1B2I2_1), .RSTB(n7575), 
        .SE(n7583), .SI(n6622), .D(n1666) );
  SDFFARX1 P1_datao_reg_3_ ( .QN(n18453), .CLK(clock_G1B2I30_1), .RSTB(n7590), 
        .SE(n7573), .SI(n18456), .D(n5996) );
  SDFFARX1 P2_reg3_reg_4_ ( .QN(n18811), .CLK(clock_G1B2I17_1), .RSTB(n7558), 
        .SE(n7571), .SI(n6684), .D(n1877) );
  SDFFARX1 P2_reg3_reg_5_ ( .QN(n18809), .CLK(clock_G1B2I17_1), .RSTB(n7558), 
        .SE(n7566), .SI(n18810), .D(n1875) );
  SDFFARX1 P2_reg3_reg_6_ ( .QN(n18807), .CLK(clock_G1B2I17_1), .RSTB(n7560), 
        .SE(n7570), .SI(n18808), .D(n1873) );
  SDFFARX1 P2_reg3_reg_7_ ( .QN(n18805), .CLK(clock_G1B2I17_1), .RSTB(n7563), 
        .SE(n7570), .SI(n18806), .D(n1871) );
  SDFFARX1 P2_reg3_reg_8_ ( .QN(n18803), .CLK(clock_G1B2I17_1), .RSTB(n7563), 
        .SE(n7570), .SI(n18804), .D(n1869) );
  SDFFARX1 P2_reg3_reg_9_ ( .QN(n18801), .CLK(clock_G1B2I7_1), .RSTB(n7563), 
        .SE(n7569), .SI(n18802), .D(n1867) );
  SDFFARX1 P2_reg3_reg_10_ ( .QN(n18799), .CLK(clock_G1B2I7_1), .RSTB(n7563), 
        .SE(n7569), .SI(n18800), .D(n1865) );
  SDFFARX1 P2_reg3_reg_11_ ( .QN(n18797), .CLK(clock_G1B2I7_1), .RSTB(n7562), 
        .SE(n7568), .SI(n18798), .D(n1863) );
  SDFFARX1 P2_reg3_reg_12_ ( .QN(n18795), .CLK(clock_G1B2I7_1), .RSTB(n7562), 
        .SE(n7571), .SI(n18796), .D(n1861) );
  SDFFARX1 P2_reg3_reg_13_ ( .QN(n18793), .CLK(clock_G1B2I9_1), .RSTB(n7562), 
        .SE(n7567), .SI(n18794), .D(n1859) );
  SDFFARX1 P2_reg3_reg_14_ ( .QN(n18791), .CLK(clock_G1B2I9_1), .RSTB(n7561), 
        .SE(n7572), .SI(n18792), .D(n1857) );
  SDFFARX1 P2_reg3_reg_15_ ( .QN(n18789), .CLK(clock_G1B2I9_1), .RSTB(n7561), 
        .SE(n7572), .SI(n18790), .D(n1855) );
  SDFFARX1 P2_reg3_reg_16_ ( .QN(n18787), .CLK(clock_G1B2I16_1), .RSTB(n7561), 
        .SE(n7565), .SI(n18788), .D(n1853) );
  SDFFARX1 P2_reg3_reg_17_ ( .QN(n18785), .CLK(clock_G1B2I16_1), .RSTB(n7502), 
        .SE(n7504), .SI(n18786), .D(n1851) );
  SDFFARX1 P2_reg3_reg_18_ ( .QN(n18783), .CLK(clock_G1B2I16_1), .RSTB(n7499), 
        .SE(n7504), .SI(n18784), .D(n1849) );
  SDFFARX1 P2_reg3_reg_19_ ( .QN(n18781), .CLK(clock_G1B2I25_1), .RSTB(n7498), 
        .SE(n7504), .SI(n18782), .D(n1847) );
  SDFFARX1 P2_reg3_reg_20_ ( .QN(n18779), .CLK(clock_G1B2I15_1), .RSTB(n7497), 
        .SE(n7506), .SI(n18780), .D(n1845) );
  SDFFARX1 P2_reg3_reg_21_ ( .QN(n18777), .CLK(clock_G1B2I15_1), .RSTB(n7497), 
        .SE(n7506), .SI(n18778), .D(n1843) );
  SDFFARX1 P2_reg3_reg_22_ ( .QN(n18775), .CLK(clock_G1B2I15_1), .RSTB(n7497), 
        .SE(n7506), .SI(n18776), .D(n1841) );
  SDFFARX1 P2_reg3_reg_23_ ( .QN(n18773), .CLK(clock_G1B2I33_1), .RSTB(n7500), 
        .SE(n7492), .SI(n18774), .D(n1839) );
  SDFFARX1 P2_reg3_reg_24_ ( .QN(n18771), .CLK(clock_G1B2I33_1), .RSTB(n7500), 
        .SE(n7496), .SI(n18772), .D(n1837) );
  SDFFARX1 P2_reg3_reg_25_ ( .QN(n18769), .CLK(clock_G1B2I33_1), .RSTB(n7500), 
        .SE(n7496), .SI(n18770), .D(n1835) );
  SDFFARX1 P2_reg3_reg_26_ ( .QN(n18767), .CLK(clock_G1B2I33_1), .RSTB(n7497), 
        .SE(n7496), .SI(n18768), .D(n1833) );
  SDFFARX1 P2_reg3_reg_27_ ( .QN(n18765), .CLK(clock_G1B2I33_1), .RSTB(n7497), 
        .SE(n7496), .SI(n18766), .D(n1831) );
  SDFFARX1 P2_reg3_reg_28_ ( .QN(n18763), .CLK(clock_G1B2I33_1), .RSTB(n7497), 
        .SE(n7506), .SI(n18764), .D(n1829) );
  SDFFARX1 P2_wr_reg ( .QN(n18189), .CLK(clock_G1B2I18_1), .RSTB(n7538), 
        .SE(n7464), .SI(n6586), .D(P2_N5476), .Q(test_so10) );
  SDFFARX1 P2_datao_reg_0_ ( .QN(n18761), .CLK(clock_G1B2I13_1), .RSTB(n7591), 
        .SE(n7599), .SI(n6592), .D(n6176) );
  SDFFARX1 P2_datao_reg_1_ ( .QN(n18759), .CLK(clock_G1B2I13_1), .RSTB(n7588), 
        .SE(n7597), .SI(n18760), .D(n6175) );
  SDFFARX1 P2_datao_reg_2_ ( .QN(n18757), .CLK(clock_G1B2I36_1), .RSTB(n7588), 
        .SE(n7597), .SI(n18758), .D(n6174) );
  SDFFARX1 P2_datao_reg_3_ ( .QN(n18755), .CLK(clock_G1B2I36_1), .RSTB(n7588), 
        .SE(n7597), .SI(n18756), .D(n6173) );
  SDFFARX1 P2_datao_reg_4_ ( .QN(n18753), .CLK(clock_G1B2I36_1), .RSTB(n7588), 
        .SE(n7595), .SI(n18754), .D(n6172) );
  SDFFARX1 P2_datao_reg_5_ ( .QN(n18751), .CLK(clock_G1B2I36_1), .RSTB(n7594), 
        .SE(n7595), .SI(n18752), .D(n6171) );
  SDFFARX1 P2_datao_reg_6_ ( .QN(n18749), .CLK(clock_G1B2I14_1), .RSTB(n6565), 
        .SE(n7596), .SI(n18750), .D(n6170) );
  SDFFARX1 P2_datao_reg_7_ ( .QN(n18747), .CLK(clock_G1B2I14_1), .RSTB(n7512), 
        .SE(n7465), .SI(n18748), .D(n6169) );
  SDFFARX1 P2_datao_reg_8_ ( .QN(n18745), .CLK(clock_G1B2I14_1), .RSTB(n7594), 
        .SE(n7595), .SI(n18746), .D(n6168) );
  SDFFARX1 P2_datao_reg_9_ ( .QN(n18743), .CLK(clock_G1B2I14_1), .RSTB(n6565), 
        .SE(n7596), .SI(n18744), .D(n6167) );
  SDFFARX1 P2_datao_reg_10_ ( .QN(n18741), .CLK(clock_G1B2I14_1), .RSTB(n6565), 
        .SE(n7596), .SI(n18742), .D(n6166) );
  SDFFARX1 P2_datao_reg_11_ ( .QN(n18739), .CLK(clock_G1B2I14_1), .RSTB(n7512), 
        .SE(n7465), .SI(n18740), .D(n6165) );
  SDFFARX1 P2_datao_reg_12_ ( .QN(n18737), .CLK(clock_G1B2I14_1), .RSTB(n6565), 
        .SE(n7596), .SI(n18738), .D(n6164) );
  SDFFARX1 P2_datao_reg_13_ ( .QN(n18735), .CLK(clock_G1B2I14_1), .RSTB(n7594), 
        .SE(n7595), .SI(n18736), .D(n6163) );
  SDFFARX1 P2_datao_reg_14_ ( .QN(n18733), .CLK(clock_G1B2I36_1), .RSTB(n7594), 
        .SE(n7595), .SI(n18734), .D(n6162) );
  SDFFARX1 P2_datao_reg_15_ ( .QN(n18731), .CLK(clock_G1B2I36_1), .RSTB(n7592), 
        .SE(n7595), .SI(n18732), .D(n6161) );
  SDFFARX1 P2_datao_reg_16_ ( .QN(n18729), .CLK(clock_G1B2I36_1), .RSTB(n7588), 
        .SE(n7597), .SI(n18730), .D(n6160) );
  SDFFARX1 P2_datao_reg_17_ ( .QN(n18727), .CLK(clock_G1B2I13_1), .RSTB(n7591), 
        .SE(n7600), .SI(n18728), .D(n6159) );
  SDFFARX1 P2_datao_reg_18_ ( .QN(n18725), .CLK(clock_G1B2I13_1), .RSTB(n7591), 
        .SE(n7600), .SI(n18726), .D(n6158) );
  SDFFARX1 P2_datao_reg_19_ ( .QN(n18723), .CLK(clock_G1B2I3_1), .RSTB(n6562), 
        .SE(n7551), .SI(n18724), .D(n6157) );
  SDFFARX1 P2_datao_reg_20_ ( .QN(n18721), .CLK(clock_G1B2I22_1), .RSTB(n7546), 
        .SE(n6574), .SI(n18722), .D(n6156) );
  SDFFARX1 P2_datao_reg_21_ ( .QN(n18719), .CLK(clock_G1B2I22_1), .RSTB(n7548), 
        .SE(n7549), .SI(n18720), .D(n6155) );
  SDFFARX1 P2_datao_reg_22_ ( .QN(n18717), .CLK(clock_G1B2I24_1), .RSTB(n7605), 
        .SE(n7489), .SI(n18718), .D(n6154) );
  SDFFARX1 P2_datao_reg_23_ ( .QN(n18715), .CLK(clock_G1B2I32_1), .RSTB(n7601), 
        .SE(n7490), .SI(n18716), .D(n6153) );
  SDFFARX1 P2_datao_reg_24_ ( .QN(n18713), .CLK(clock_G1B2I32_1), .RSTB(n7601), 
        .SE(n7490), .SI(n18714), .D(n6152) );
  SDFFARX1 P2_datao_reg_25_ ( .QN(n18711), .CLK(clock_G1B2I32_1), .RSTB(n7601), 
        .SE(n7491), .SI(n18712), .D(n6151) );
  SDFFARX1 P2_datao_reg_26_ ( .QN(n18709), .CLK(clock_G1B2I32_1), .RSTB(n7602), 
        .SE(n7491), .SI(n18710), .D(n6150) );
  SDFFARX1 P2_datao_reg_27_ ( .QN(n18707), .CLK(clock_G1B2I32_1), .RSTB(n7602), 
        .SE(n7491), .SI(n18708), .D(n6149) );
  SDFFARX1 P2_datao_reg_28_ ( .QN(n18705), .CLK(clock_G1B2I32_1), .RSTB(n7602), 
        .SE(n7491), .SI(n18706), .D(n6148) );
  SDFFARX1 P1_IR_reg_28_ ( .QN(n18703), .CLK(clock_G1B2I38_1), .RSTB(n7519), 
        .SE(n7528), .SI(n18698), .D(n6112) );
  SDFFARX1 P1_IR_reg_30_ ( .QN(n18701), .CLK(clock_G1B2I38_1), .RSTB(n7519), 
        .SE(n7528), .SI(n18696), .D(n6110) );
  SDFFARX1 P1_IR_reg_27_ ( .QN(n18699), .CLK(clock_G1B2I38_1), .RSTB(n7519), 
        .SE(n7528), .SI(n18668), .D(n6113) );
  SDFFARX1 P1_IR_reg_29_ ( .QN(n18697), .CLK(clock_G1B2I38_1), .RSTB(n7519), 
        .SE(n7528), .SI(n18702), .D(n6111) );
  SDFFARX1 P1_IR_reg_0_ ( .QN(n18695), .CLK(clock_G1B2I8_1), .RSTB(n7520), 
        .SE(n7529), .SI(n6618), .D(n6140) );
  SDFFARX1 P1_IR_reg_1_ ( .QN(n18693), .CLK(clock_G1B2I4_1), .RSTB(n7469), 
        .SE(n7474), .SI(n6624), .D(n6139) );
  SDFFARX1 P1_IR_reg_2_ ( .QN(n18691), .CLK(clock_G1B2I4_1), .RSTB(n7468), 
        .SE(n7474), .SI(n6625), .D(n6138) );
  SDFFARX1 P1_IR_reg_3_ ( .QN(n18689), .CLK(clock_G1B2I4_1), .RSTB(n7468), 
        .SE(n7472), .SI(n6626), .D(n6137) );
  SDFFARX1 P1_IR_reg_4_ ( .QN(n18687), .CLK(clock_G1B2I4_1), .RSTB(n7468), 
        .SE(n7472), .SI(n6627), .D(n6136) );
  SDFFARX1 P1_IR_reg_5_ ( .QN(n18685), .CLK(clock_G1B2I4_1), .RSTB(n7471), 
        .SE(n7472), .SI(n6628), .D(n6135) );
  SDFFARX1 P1_IR_reg_6_ ( .QN(n18683), .CLK(clock_G1B2I4_1), .RSTB(n7470), 
        .SE(n7473), .SI(n6629), .D(n6134) );
  SDFFARX1 P1_IR_reg_7_ ( .QN(n18681), .CLK(clock_G1B2I4_1), .RSTB(n7470), 
        .SE(n7473), .SI(n6630), .D(n6133) );
  SDFFARX1 P1_IR_reg_8_ ( .QN(n18679), .CLK(clock_G1B2I4_1), .RSTB(n7471), 
        .SE(n7474), .SI(n6631), .D(n6132) );
  SDFFARX1 P1_IR_reg_9_ ( .QN(n18677), .CLK(clock_G1B2I4_1), .RSTB(n7470), 
        .SE(n7473), .SI(n6632), .D(n6131) );
  SDFFARX1 P1_IR_reg_10_ ( .QN(n18675), .CLK(clock_G1B2I4_1), .RSTB(n7470), 
        .SE(n7473), .SI(n6633), .D(n6130) );
  SDFFARX1 P1_IR_reg_11_ ( .QN(n18673), .CLK(clock_G1B2I4_1), .RSTB(n7470), 
        .SE(n7473), .SI(n6634), .D(n6129) );
  SDFFARX1 P1_IR_reg_12_ ( .QN(n18671), .CLK(clock_G1B2I4_1), .RSTB(n7470), 
        .SE(n7473), .SI(n6635), .D(n6128) );
  SDFFARX1 P1_IR_reg_26_ ( .QN(n18669), .CLK(clock_G1B2I38_1), .RSTB(n7521), 
        .SE(n7528), .SI(n18666), .D(n6114) );
  SDFFARX1 P1_IR_reg_25_ ( .QN(n18667), .CLK(clock_G1B2I38_1), .RSTB(n7521), 
        .SE(n7529), .SI(n18664), .D(n6115) );
  SDFFARX1 P1_IR_reg_24_ ( .QN(n18665), .CLK(clock_G1B2I8_1), .RSTB(n7520), 
        .SE(n7529), .SI(n6637), .D(n6116) );
  SDFFARX1 P1_IR_reg_23_ ( .QN(n18663), .CLK(clock_G1B2I8_1), .RSTB(n7520), 
        .SE(n7529), .SI(n6638), .D(n6117) );
  SDFFARX1 P1_IR_reg_22_ ( .QN(n18661), .CLK(clock_G1B2I8_1), .RSTB(n7520), 
        .SE(n7529), .SI(n6639), .D(n6118) );
  SDFFARX1 P1_IR_reg_21_ ( .QN(n18659), .CLK(clock_G1B2I8_1), .RSTB(n7520), 
        .SE(n7530), .SI(n6640), .D(n6119) );
  SDFFARX1 P1_IR_reg_20_ ( .QN(n18657), .CLK(clock_G1B2I8_1), .RSTB(n7469), 
        .SE(n7475), .SI(n6641), .D(n6120) );
  SDFFARX1 P1_IR_reg_19_ ( .QN(n18655), .CLK(clock_G1B2I8_1), .RSTB(n7469), 
        .SE(n7475), .SI(n6642), .D(n6121) );
  SDFFARX1 P1_IR_reg_18_ ( .QN(n18653), .CLK(clock_G1B2I8_1), .RSTB(n7469), 
        .SE(n7474), .SI(n6643), .D(n6122) );
  SDFFARX1 P1_IR_reg_17_ ( .QN(n18651), .CLK(clock_G1B2I8_1), .RSTB(n7469), 
        .SE(n7474), .SI(n6644), .D(n6123) );
  SDFFARX1 P1_IR_reg_16_ ( .QN(n18649), .CLK(clock_G1B2I4_1), .RSTB(n7469), 
        .SE(n7474), .SI(n6645), .D(n6124) );
  SDFFARX1 P1_IR_reg_15_ ( .QN(n18647), .CLK(clock_G1B2I4_1), .RSTB(n7468), 
        .SE(n7472), .SI(n6646), .D(n6125) );
  SDFFARX1 P1_IR_reg_14_ ( .QN(n18645), .CLK(clock_G1B2I4_1), .RSTB(n7468), 
        .SE(n7472), .SI(n6647), .D(n6126) );
  SDFFARX1 P1_IR_reg_13_ ( .QN(n18643), .CLK(clock_G1B2I4_1), .RSTB(n7468), 
        .SE(n7472), .SI(n6636), .D(n6127) );
  SDFFARX1 P1_wr_reg ( .QN(n18183), .CLK(clock_G1B2I19_1), .RSTB(n6560), 
        .SE(n7466), .SI(n6582), .D(P1_N5554), .Q(test_so5) );
  SDFFARX1 P1_reg2_reg_0_ ( .QN(n1504), .CLK(clock_G1B2I20_1), .RSTB(n7579), 
        .SE(n6569), .SI(n18526), .D(n6049) );
  SDFFARX1 P1_reg2_reg_1_ ( .QN(n18641), .CLK(clock_G1B2I28_1), .RSTB(n6557), 
        .SE(n6569), .SI(n18195), .D(n6048) );
  SDFFARX1 P1_reg2_reg_2_ ( .QN(n18639), .CLK(clock_G1B2I2_1), .RSTB(n6557), 
        .SE(n7581), .SI(n18640), .D(n6047) );
  SDFFARX1 P1_reg2_reg_3_ ( .QN(n18637), .CLK(clock_G1B2I2_1), .RSTB(n6557), 
        .SE(n7581), .SI(n18638), .D(n6046) );
  SDFFARX1 P1_reg2_reg_4_ ( .QN(n18635), .CLK(clock_G1B2I28_1), .RSTB(n7574), 
        .SE(n7587), .SI(n18636), .D(n6045) );
  SDFFARX1 P1_reg2_reg_5_ ( .QN(n18633), .CLK(clock_G1B2I10_1), .RSTB(n7531), 
        .SE(n7536), .SI(n18634), .D(n6044) );
  SDFFARX1 P2_reg2_reg_3_ ( .QN(n18993), .CLK(clock_G1B2I12_1), .RSTB(n7548), 
        .SE(n7551), .SI(n6721), .D(n6226) );
  SDFFARX1 P2_reg2_reg_4_ ( .QN(n18991), .CLK(clock_G1B2I12_1), .RSTB(n7548), 
        .SE(n7551), .SI(n6648), .D(n6225) );
  SDFFARX1 P2_reg2_reg_5_ ( .QN(n18989), .CLK(clock_G1B2I13_1), .RSTB(n7589), 
        .SE(n7600), .SI(n6649), .D(n6224) );
  SDFFARX1 P2_reg2_reg_6_ ( .QN(n18987), .CLK(clock_G1B2I13_1), .RSTB(n7589), 
        .SE(n7599), .SI(n6650), .D(n6223) );
  SDFFARX1 P2_reg2_reg_7_ ( .QN(n18985), .CLK(clock_G1B2I13_1), .RSTB(n7589), 
        .SE(n7599), .SI(n6651), .D(n6222) );
  SDFFARX1 P2_reg2_reg_8_ ( .QN(n18983), .CLK(clock_G1B2I13_1), .RSTB(n7589), 
        .SE(n7599), .SI(n6652), .D(n6221) );
  SDFFARX1 P2_reg2_reg_9_ ( .QN(n18981), .CLK(clock_G1B2I17_1), .RSTB(n7558), 
        .SE(n7566), .SI(n6653), .D(n6220) );
  SDFFARX1 P2_reg2_reg_10_ ( .QN(n18979), .CLK(clock_G1B2I17_1), .RSTB(n7557), 
        .SE(n7566), .SI(n6654), .D(n6219) );
  SDFFARX1 P2_reg2_reg_11_ ( .QN(n18977), .CLK(clock_G1B2I7_1), .RSTB(n7557), 
        .SE(n7569), .SI(n6655), .D(n6218) );
  SDFFARX1 P2_reg2_reg_12_ ( .QN(n18975), .CLK(clock_G1B2I9_1), .RSTB(n6559), 
        .SE(n7568), .SI(n6656), .D(n6217) );
  SDFFARX1 P2_reg2_reg_13_ ( .QN(n18973), .CLK(clock_G1B2I9_1), .RSTB(n6559), 
        .SE(n7567), .SI(n6657), .D(n6216) );
  SDFFARX1 P2_reg2_reg_14_ ( .QN(n18971), .CLK(clock_G1B2I9_1), .RSTB(n6559), 
        .SE(n7572), .SI(n6658), .D(n6215) );
  SDFFARX1 P2_reg2_reg_15_ ( .QN(n18969), .CLK(clock_G1B2I16_1), .RSTB(n7564), 
        .SE(n7565), .SI(n6659), .D(n6214) );
  SDFFARX1 P2_reg2_reg_16_ ( .QN(n18967), .CLK(clock_G1B2I16_1), .RSTB(n7502), 
        .SE(n7504), .SI(n6660), .D(n6213) );
  SDFFARX1 P2_reg2_reg_17_ ( .QN(n18965), .CLK(clock_G1B2I16_1), .RSTB(n7502), 
        .SE(n7503), .SI(n6661), .D(n6212) );
  SDFFARX1 P2_reg2_reg_18_ ( .QN(n18963), .CLK(clock_G1B2I16_1), .RSTB(n7499), 
        .SE(n7503), .SI(n6662), .D(n6211) );
  SDFFARX1 P2_reg2_reg_19_ ( .QN(n18191), .CLK(clock_G1B2I25_1), .RSTB(n7498), 
        .SE(n7503), .SI(n6663), .D(n6210), .Q(test_so9) );
  SDFFARX1 P2_reg2_reg_20_ ( .QN(n18961), .CLK(clock_G1B2I22_1), .RSTB(n7548), 
        .SE(n6574), .SI(test_si10), .D(n6209) );
  SDFFARX1 P2_reg2_reg_21_ ( .QN(n18959), .CLK(clock_G1B2I25_1), .RSTB(n7501), 
        .SE(n7505), .SI(n18960), .D(n6208) );
  SDFFARX1 P2_reg2_reg_22_ ( .QN(n18957), .CLK(clock_G1B2I15_1), .RSTB(n7502), 
        .SE(n7505), .SI(n18958), .D(n6207) );
  SDFFARX1 P2_reg2_reg_23_ ( .QN(n18955), .CLK(clock_G1B2I33_1), .RSTB(n6558), 
        .SE(n7450), .SI(n18956), .D(n6206) );
  SDFFARX1 P2_reg2_reg_24_ ( .QN(n18953), .CLK(clock_G1B2I6_1), .RSTB(n7605), 
        .SE(n7494), .SI(n18954), .D(n6205) );
  SDFFARX1 P2_reg2_reg_25_ ( .QN(n18951), .CLK(clock_G1B2I5_1), .RSTB(n7603), 
        .SE(n7494), .SI(n18952), .D(n6204) );
  SDFFARX1 P2_reg2_reg_26_ ( .QN(n18949), .CLK(clock_G1B2I5_1), .RSTB(n7603), 
        .SE(n7494), .SI(n18950), .D(n6203) );
  SDFFARX1 P2_reg2_reg_27_ ( .QN(n18947), .CLK(clock_G1B2I5_1), .RSTB(n7603), 
        .SE(n7493), .SI(n18948), .D(n6202) );
  SDFFARX1 P2_reg2_reg_28_ ( .QN(n18945), .CLK(clock_G1B2I5_1), .RSTB(n7602), 
        .SE(n7493), .SI(n18946), .D(n6201) );
  SDFFARX1 P2_reg2_reg_29_ ( .QN(n18943), .CLK(clock_G1B2I5_1), .RSTB(n7602), 
        .SE(n7491), .SI(n18944), .D(n6200) );
  SDFFARX1 P2_reg1_reg_0_ ( .QN(n18941), .CLK(clock_G1B2I12_1), .RSTB(n7547), 
        .SE(n7552), .SI(n18820), .D(n6259) );
  SDFFARX1 P2_reg1_reg_1_ ( .QN(n18939), .CLK(clock_G1B2I12_1), .RSTB(n7547), 
        .SE(n7552), .SI(n18940), .D(n6258) );
  SDFFARX1 P2_reg1_reg_2_ ( .QN(n18937), .CLK(clock_G1B2I12_1), .RSTB(n7547), 
        .SE(n7551), .SI(n6664), .D(n6257) );
  SDFFARX1 P2_reg1_reg_3_ ( .QN(n18935), .CLK(clock_G1B2I12_1), .RSTB(n7548), 
        .SE(n7551), .SI(n6665), .D(n6256) );
  SDFFARX1 P2_reg1_reg_4_ ( .QN(n18933), .CLK(clock_G1B2I12_1), .RSTB(n7559), 
        .SE(n7573), .SI(n6666), .D(n6255) );
  SDFFARX1 P2_reg1_reg_5_ ( .QN(n18931), .CLK(clock_G1B2I12_1), .RSTB(n7559), 
        .SE(n7573), .SI(n6667), .D(n6254) );
  SDFFARX1 P2_reg1_reg_6_ ( .QN(n18929), .CLK(clock_G1B2I30_1), .RSTB(n7592), 
        .SE(n7449), .SI(n6668), .D(n6253) );
  SDFFARX1 P2_reg1_reg_7_ ( .QN(n18927), .CLK(clock_G1B2I30_1), .RSTB(n7592), 
        .SE(n7587), .SI(n6669), .D(n6252) );
  SDFFARX1 P2_reg1_reg_8_ ( .QN(n18190), .CLK(clock_G1B2I17_1), .RSTB(n7558), 
        .SE(n7566), .SI(n6670), .D(n6251), .Q(test_so8) );
  SDFFARX1 P2_reg1_reg_9_ ( .QN(n18925), .CLK(clock_G1B2I13_1), .RSTB(n7591), 
        .SE(n7599), .SI(test_si9), .D(n6250) );
  SDFFARX1 P2_reg1_reg_10_ ( .QN(n18923), .CLK(clock_G1B2I17_1), .RSTB(n7557), 
        .SE(n7566), .SI(n6671), .D(n6249) );
  SDFFARX1 P2_reg1_reg_11_ ( .QN(n18921), .CLK(clock_G1B2I7_1), .RSTB(n7557), 
        .SE(n7569), .SI(n6672), .D(n6248) );
  SDFFARX1 P2_reg1_reg_12_ ( .QN(n18919), .CLK(clock_G1B2I7_1), .RSTB(n7559), 
        .SE(n7568), .SI(n6673), .D(n6247) );
  SDFFARX1 P2_reg1_reg_13_ ( .QN(n18917), .CLK(clock_G1B2I9_1), .RSTB(n6559), 
        .SE(n7567), .SI(n6674), .D(n6246) );
  SDFFARX1 P2_reg1_reg_14_ ( .QN(n18915), .CLK(clock_G1B2I9_1), .RSTB(n7563), 
        .SE(n7565), .SI(n6675), .D(n6245) );
  SDFFARX1 P2_reg1_reg_15_ ( .QN(n18913), .CLK(clock_G1B2I16_1), .RSTB(n7561), 
        .SE(n7565), .SI(n6676), .D(n6244) );
  SDFFARX1 P2_reg1_reg_16_ ( .QN(n18911), .CLK(clock_G1B2I16_1), .RSTB(n7564), 
        .SE(n7565), .SI(n6677), .D(n6243) );
  SDFFARX1 P2_reg1_reg_17_ ( .QN(n18909), .CLK(clock_G1B2I16_1), .RSTB(n7499), 
        .SE(n7503), .SI(n6678), .D(n6242) );
  SDFFARX1 P2_reg1_reg_18_ ( .QN(n18907), .CLK(clock_G1B2I25_1), .RSTB(n7499), 
        .SE(n7503), .SI(n6679), .D(n6241) );
  SDFFARX1 P2_reg1_reg_19_ ( .QN(n18905), .CLK(clock_G1B2I25_1), .RSTB(n7498), 
        .SE(n7506), .SI(n6680), .D(n6240) );
  SDFFARX1 P2_reg1_reg_20_ ( .QN(n18903), .CLK(clock_G1B2I25_1), .RSTB(n7498), 
        .SE(n6573), .SI(n18904), .D(n6239) );
  SDFFARX1 P2_reg1_reg_21_ ( .QN(n18901), .CLK(clock_G1B2I15_1), .RSTB(n7500), 
        .SE(n7505), .SI(n18902), .D(n6238) );
  SDFFARX1 P2_reg1_reg_22_ ( .QN(n18899), .CLK(clock_G1B2I15_1), .RSTB(n7502), 
        .SE(n7505), .SI(n18900), .D(n6237) );
  SDFFARX1 P2_reg1_reg_23_ ( .QN(n18897), .CLK(clock_G1B2I6_1), .RSTB(n6558), 
        .SE(n7450), .SI(n18898), .D(n6236) );
  SDFFARX1 P2_reg1_reg_24_ ( .QN(n18895), .CLK(clock_G1B2I6_1), .RSTB(n7604), 
        .SE(n7495), .SI(n18896), .D(n6235) );
  SDFFARX1 P2_reg1_reg_25_ ( .QN(n18893), .CLK(clock_G1B2I6_1), .RSTB(n7604), 
        .SE(n7495), .SI(n18894), .D(n6234) );
  SDFFARX1 P2_reg1_reg_26_ ( .QN(n18891), .CLK(clock_G1B2I6_1), .RSTB(n7604), 
        .SE(n7495), .SI(n18892), .D(n6233) );
  SDFFARX1 P2_reg1_reg_27_ ( .QN(n18889), .CLK(clock_G1B2I5_1), .RSTB(n7605), 
        .SE(n7493), .SI(n18890), .D(n6232) );
  SDFFARX1 P2_reg1_reg_28_ ( .QN(n18887), .CLK(clock_G1B2I5_1), .RSTB(n7602), 
        .SE(n7493), .SI(n18888), .D(n6231) );
  SDFFARX1 P2_reg1_reg_29_ ( .QN(n18885), .CLK(clock_G1B2I5_1), .RSTB(n7601), 
        .SE(n7495), .SI(n18886), .D(n6230) );
  SDFFARX1 P2_reg1_reg_31_ ( .QN(n18883), .CLK(clock_G1B2I6_1), .RSTB(n6558), 
        .SE(n7450), .SI(n18202), .D(n5956) );
  SDFFARX1 P2_reg0_reg_0_ ( .QN(n18881), .CLK(clock_G1B2I9_1), .RSTB(n6559), 
        .SE(n7572), .SI(n18295), .D(n6289) );
  SDFFARX1 P2_reg0_reg_1_ ( .QN(n18879), .CLK(clock_G1B2I9_1), .RSTB(n6559), 
        .SE(n7567), .SI(n18880), .D(n6288) );
  SDFFARX1 P2_reg0_reg_2_ ( .QN(n18877), .CLK(clock_G1B2I7_1), .RSTB(n7559), 
        .SE(n7568), .SI(n18878), .D(n6287) );
  SDFFARX1 P2_reg0_reg_3_ ( .QN(n18875), .CLK(clock_G1B2I7_1), .RSTB(n7557), 
        .SE(n7568), .SI(n18876), .D(n6286) );
  SDFFARX1 P2_reg0_reg_4_ ( .QN(n18873), .CLK(clock_G1B2I7_1), .RSTB(n7557), 
        .SE(n7569), .SI(n18874), .D(n6285) );
  SDFFARX1 P2_reg0_reg_5_ ( .QN(n18871), .CLK(clock_G1B2I17_1), .RSTB(n7558), 
        .SE(n7569), .SI(n18872), .D(n6284) );
  SDFFARX1 P2_reg0_reg_6_ ( .QN(n18869), .CLK(clock_G1B2I17_1), .RSTB(n7558), 
        .SE(n7566), .SI(n18870), .D(n6283) );
  SDFFARX1 P2_reg0_reg_7_ ( .QN(n18867), .CLK(clock_G1B2I17_1), .RSTB(n7560), 
        .SE(n7571), .SI(n18868), .D(n6282) );
  SDFFARX1 P2_reg0_reg_8_ ( .QN(n18865), .CLK(clock_G1B2I17_1), .RSTB(n7560), 
        .SE(n7570), .SI(n18866), .D(n6281) );
  SDFFARX1 P2_reg0_reg_9_ ( .QN(n18863), .CLK(clock_G1B2I17_1), .RSTB(n7560), 
        .SE(n7570), .SI(n18864), .D(n6280) );
  SDFFARX1 P2_reg0_reg_10_ ( .QN(n18861), .CLK(clock_G1B2I17_1), .RSTB(n7560), 
        .SE(n7570), .SI(n18862), .D(n6279) );
  SDFFARX1 P2_reg0_reg_11_ ( .QN(n18859), .CLK(clock_G1B2I7_1), .RSTB(n7563), 
        .SE(n7571), .SI(n18860), .D(n6278) );
  SDFFARX1 P2_reg0_reg_12_ ( .QN(n18857), .CLK(clock_G1B2I7_1), .RSTB(n7562), 
        .SE(n7571), .SI(n18858), .D(n6277) );
  SDFFARX1 P2_reg0_reg_13_ ( .QN(n18855), .CLK(clock_G1B2I9_1), .RSTB(n7562), 
        .SE(n7572), .SI(n18856), .D(n6276) );
  SDFFARX1 P2_reg0_reg_14_ ( .QN(n18853), .CLK(clock_G1B2I9_1), .RSTB(n7562), 
        .SE(n7567), .SI(n18854), .D(n6275) );
  SDFFARX1 P2_reg0_reg_15_ ( .QN(n18851), .CLK(clock_G1B2I9_1), .RSTB(n7561), 
        .SE(n7572), .SI(n18852), .D(n6274) );
  SDFFARX1 P2_reg0_reg_16_ ( .QN(n18849), .CLK(clock_G1B2I16_1), .RSTB(n7561), 
        .SE(n7565), .SI(n18850), .D(n6273) );
  SDFFARX1 P2_reg0_reg_17_ ( .QN(n18847), .CLK(clock_G1B2I16_1), .RSTB(n7499), 
        .SE(n7504), .SI(n18848), .D(n6272) );
  SDFFARX1 P2_reg0_reg_18_ ( .QN(n18845), .CLK(clock_G1B2I16_1), .RSTB(n7499), 
        .SE(n7503), .SI(n18846), .D(n6271) );
  SDFFARX1 P2_reg0_reg_19_ ( .QN(n18843), .CLK(clock_G1B2I25_1), .RSTB(n7498), 
        .SE(n7504), .SI(n18844), .D(n6270) );
  SDFFARX1 P2_reg0_reg_20_ ( .QN(n18841), .CLK(clock_G1B2I25_1), .RSTB(n7498), 
        .SE(n7506), .SI(n18842), .D(n6269) );
  SDFFARX1 P2_reg0_reg_21_ ( .QN(n18839), .CLK(clock_G1B2I15_1), .RSTB(n7500), 
        .SE(n7505), .SI(n18840), .D(n6268) );
  SDFFARX1 P2_reg0_reg_22_ ( .QN(n18837), .CLK(clock_G1B2I15_1), .RSTB(n7500), 
        .SE(n7505), .SI(n18838), .D(n6267) );
  SDFFARX1 P2_reg0_reg_23_ ( .QN(n18835), .CLK(clock_G1B2I6_1), .RSTB(n6558), 
        .SE(n7450), .SI(n18836), .D(n6266) );
  SDFFARX1 P2_reg0_reg_24_ ( .QN(n18833), .CLK(clock_G1B2I6_1), .RSTB(n7604), 
        .SE(n7495), .SI(n18834), .D(n6265) );
  SDFFARX1 P2_reg0_reg_25_ ( .QN(n18831), .CLK(clock_G1B2I6_1), .RSTB(n7603), 
        .SE(n7494), .SI(n18832), .D(n6264) );
  SDFFARX1 P2_reg0_reg_26_ ( .QN(n18829), .CLK(clock_G1B2I6_1), .RSTB(n7603), 
        .SE(n7494), .SI(n18830), .D(n6263) );
  SDFFARX1 P2_reg0_reg_27_ ( .QN(n18827), .CLK(clock_G1B2I5_1), .RSTB(n7603), 
        .SE(n7494), .SI(n18828), .D(n6262) );
  SDFFARX1 P2_reg0_reg_28_ ( .QN(n18825), .CLK(clock_G1B2I5_1), .RSTB(n7604), 
        .SE(n7493), .SI(n18826), .D(n6261) );
  SDFFARX1 P2_reg0_reg_29_ ( .QN(n18823), .CLK(clock_G1B2I5_1), .RSTB(n7605), 
        .SE(n7493), .SI(n18824), .D(n6260) );
  SDFFARX1 P2_reg0_reg_31_ ( .QN(n18821), .CLK(clock_G1B2I6_1), .RSTB(n6558), 
        .SE(n7450), .SI(n18200), .D(n5955) );
  SDFFARX1 P2_reg3_reg_0_ ( .QN(n18819), .CLK(clock_G1B2I25_1), .RSTB(n7501), 
        .SE(n6573), .SI(n19012), .D(n1885) );
  SDFFARX1 P2_reg3_reg_1_ ( .QN(n18817), .CLK(clock_G1B2I7_1), .RSTB(n7559), 
        .SE(n7567), .SI(n6681), .D(n1883) );
  SDFFARX1 P2_reg3_reg_2_ ( .QN(n18815), .CLK(clock_G1B2I7_1), .RSTB(n7559), 
        .SE(n7568), .SI(n6682), .D(n1881) );
  SDFFARX1 P2_reg3_reg_3_ ( .QN(n18813), .CLK(clock_G1B2I17_1), .RSTB(n7560), 
        .SE(n7571), .SI(n6683), .D(n1879) );
  AND2X1 P1_C21519 ( .IN1(P1_N536), .IN2(P1_N530), .Q(P1_N6363) );
  AND2X1 P1_C21520 ( .IN1(n7271), .IN2(n6620), .Q(P1_N6364) );
  AND2X1 P1_C21692 ( .IN1(P1_N536), .IN2(P1_N531), .Q(P1_N6425) );
  AND2X1 P1_C21693 ( .IN1(n7271), .IN2(n6619), .Q(P1_N6426) );
  AND2X1 P1_C21696 ( .IN1(P1_N536), .IN2(P1_N530), .Q(P1_N6427) );
  AND2X1 P1_C21697 ( .IN1(n7271), .IN2(n6620), .Q(P1_N6428) );
  AND2X1 P1_C21872 ( .IN1(P1_N536), .IN2(P1_N531), .Q(P1_N6489) );
  AND2X1 P1_C21873 ( .IN1(n7271), .IN2(n6619), .Q(P1_N6490) );
  AND2X1 P1_C21876 ( .IN1(P1_N536), .IN2(P1_N530), .Q(P1_N6491) );
  AND2X1 P1_C21877 ( .IN1(n7271), .IN2(n6620), .Q(P1_N6492) );
  AND2X1 P1_C22049 ( .IN1(P1_N536), .IN2(P1_N531), .Q(P1_N6553) );
  AND2X1 P1_C22050 ( .IN1(n7271), .IN2(n6619), .Q(P1_N6554) );
  AND2X1 P1_C22053 ( .IN1(P1_N536), .IN2(P1_N530), .Q(P1_N6555) );
  AND2X1 P1_C22054 ( .IN1(n7271), .IN2(n6620), .Q(P1_N6556) );
  AND2X1 P1_C22226 ( .IN1(P1_N536), .IN2(P1_N531), .Q(P1_N6617) );
  AND2X1 P1_C22227 ( .IN1(n7271), .IN2(n6619), .Q(P1_N6618) );
  AND2X1 P1_C22230 ( .IN1(P1_N536), .IN2(P1_N530), .Q(P1_N6619) );
  AND2X1 P1_C22231 ( .IN1(n7271), .IN2(n6620), .Q(P1_N6620) );
  AND2X1 P1_C22410 ( .IN1(P1_N536), .IN2(P1_N531), .Q(P1_N6681) );
  AND2X1 P1_C22411 ( .IN1(n7271), .IN2(n6619), .Q(P1_N6682) );
  AND2X1 P1_C22414 ( .IN1(P1_N536), .IN2(P1_N530), .Q(P1_N6683) );
  AND2X1 P1_C22415 ( .IN1(n7271), .IN2(n6620), .Q(P1_N6684) );
  OR2X1 P1_C22512 ( .IN2(n6618), .IN1(P1_N5137), .Q(P1_N5284) );
  OR2X1 P1_C22515 ( .IN2(n6618), .IN1(P1_N6685), .Q(P1_N5286) );
  OR2X1 P1_C22519 ( .IN2(n6618), .IN1(P1_N5140), .Q(P1_N5288) );
  OR2X1 P1_C22522 ( .IN2(n6618), .IN1(P1_N6686), .Q(P1_N5290) );
  OR2X1 P1_C22526 ( .IN2(n6618), .IN1(n14521), .Q(P1_N5292) );
  OR2X1 P1_C22530 ( .IN2(n6618), .IN1(P1_N5143), .Q(P1_N5294) );
  OR2X1 P1_C22536 ( .IN2(n6618), .IN1(P1_N5362), .Q(P1_N5363) );
  OR2X1 P1_C22542 ( .IN2(n6618), .IN1(P1_N6688), .Q(P1_N5432) );
  AND2X1 C109 ( .IN1(n18245), .IN2(n18209), .Q(N76) );
  AND2X1 C108 ( .IN1(N76), .IN2(N71), .Q(N77) );
  AND2X1 C106 ( .IN1(n18246), .IN2(n18210), .Q(N73) );
  AND2X1 C105 ( .IN1(N73), .IN2(N74), .Q(N75) );
  OR2X1 C104 ( .IN2(N77), .IN1(N75), .Q(N5) );
  SDFFARX1 P2_IR_reg_31_ ( .QN(n19025), .CLK(clock_G1B2I30_1), .RSTB(n7590), 
        .SE(Scan_Enable), .SI(n19020), .D(n6318) );
  SDFFARX1 P2_datao_reg_30_ ( .QN(n18193), .CLK(clock_G1B2I32_1), .RSTB(n7601), 
        .SE(n7490), .SI(n19018), .D(n6143), .Q(test_so7) );
  SDFFARX1 P1_reg0_reg_30_ ( .QN(n19023), .CLK(clock_G1B2I2_1), .RSTB(n7575), 
        .SE(n7581), .SI(n18466), .D(n5964) );
  SDFFARX1 P1_datao_reg_30_ ( .QN(n18192), .CLK(clock_G1B2I24_1), .RSTB(n7606), 
        .SE(n7489), .SI(n19006), .D(n5966), .Q(test_so2) );
  SDFFARX1 P2_IR_reg_30_ ( .QN(n19021), .CLK(clock_G1B2I3_1), .RSTB(n7541), 
        .SE(n7556), .SI(n19004), .D(n6317) );
  SDFFARX1 P2_datao_reg_29_ ( .QN(n19019), .CLK(clock_G1B2I32_1), .RSTB(n7601), 
        .SE(n7491), .SI(n18704), .D(n6144) );
  SDFFARX1 P1_reg0_reg_31_ ( .QN(n19017), .CLK(clock_G1B2I20_1), .RSTB(n7579), 
        .SE(n6569), .SI(n19022), .D(n5963) );
  SDFFARX1 P1_datao_reg_31_ ( .QN(n19015), .CLK(clock_G1B2I11_1), .RSTB(n7471), 
        .SE(n6578), .SI(test_si3), .D(n5965) );
  SDFFARX1 P2_reg2_reg_31_ ( .QN(n19013), .CLK(clock_G1B2I6_1), .RSTB(n6558), 
        .SE(n7496), .SI(n18198), .D(n5953) );
  SDFFARX1 P2_datao_reg_31_ ( .QN(n19011), .CLK(clock_G1B2I22_1), .RSTB(n7546), 
        .SE(n6574), .SI(test_si8), .D(n6142) );
  SDFFARX1 P1_IR_reg_31_ ( .QN(n19009), .CLK(clock_G1B2I8_1), .RSTB(n7520), 
        .SE(n7529), .SI(n18700), .D(n6141) );
  SDFFARX1 P1_datao_reg_29_ ( .QN(n19007), .CLK(clock_G1B2I24_1), .RSTB(n7606), 
        .SE(n7489), .SI(n18352), .D(n5967) );
  SDFFARX1 P2_IR_reg_29_ ( .QN(n19005), .CLK(clock_G1B2I3_1), .RSTB(n6562), 
        .SE(n7555), .SI(n18350), .D(n6177) );
  SDFFARX1 P2_addr_reg_0_ ( .QN(n19003), .CLK(clock_G1B2I26_1), .RSTB(n7544), 
        .SE(n7452), .SI(n6688), .D(n6197) );
  SDFFARX1 P2_IR_reg_23_ ( .QN(n19001), .CLK(clock_G1B2I30_1), .RSTB(n7590), 
        .SE(Scan_Enable), .SI(n6608), .D(n6293) );
  SDFFARX1 P2_reg2_reg_0_ ( .QN(n18999), .CLK(clock_G1B2I12_1), .RSTB(n7547), 
        .SE(n7552), .SI(n18882), .D(n6229) );
  SDFFARX1 P2_reg2_reg_1_ ( .QN(n18997), .CLK(clock_G1B2I12_1), .RSTB(n7547), 
        .SE(n7552), .SI(n18998), .D(n6228) );
  SDFFARX1 P2_reg2_reg_2_ ( .QN(n18995), .CLK(clock_G1B2I12_1), .RSTB(n7547), 
        .SE(n7551), .SI(n6720), .D(n6227) );
  AND2X1 P1_C20200 ( .IN1(n6716), .IN2(P1_N106), .Q(P1_N5897) );
  AND2X1 P1_C20201 ( .IN1(n6715), .IN2(n6628), .Q(P1_N5898) );
  OR2X1 P1_C20203 ( .IN2(P1_N5900), .IN1(P1_N5899), .Q(P1_N423) );
  AND2X1 P1_C20204 ( .IN1(n6704), .IN2(P1_N105), .Q(P1_N5899) );
  AND2X1 P1_C20205 ( .IN1(n6703), .IN2(n6627), .Q(P1_N5900) );
  OR2X1 P1_C20207 ( .IN2(P1_N5902), .IN1(P1_N5901), .Q(P1_N424) );
  AND2X1 P1_C20208 ( .IN1(n6704), .IN2(P1_N104), .Q(P1_N5901) );
  AND2X1 P1_C20209 ( .IN1(n6703), .IN2(n6626), .Q(P1_N5902) );
  OR2X1 P1_C20211 ( .IN2(P1_N5904), .IN1(P1_N5903), .Q(P1_N425) );
  AND2X1 P1_C20212 ( .IN1(n6704), .IN2(P1_N103), .Q(P1_N5903) );
  AND2X1 P1_C20213 ( .IN1(n6703), .IN2(n6625), .Q(P1_N5904) );
  OR2X1 P1_C20215 ( .IN2(P1_N5906), .IN1(P1_N5905), .Q(P1_N426) );
  AND2X1 P1_C20216 ( .IN1(n6704), .IN2(n6624), .Q(P1_N5905) );
  AND2X1 P1_C20217 ( .IN1(n6703), .IN2(n6624), .Q(P1_N5906) );
  AND2X1 P1_C20453 ( .IN1(P1_N536), .IN2(P1_N531), .Q(P1_N5977) );
  AND2X1 P1_C20454 ( .IN1(n7271), .IN2(n6619), .Q(P1_N5978) );
  AND2X1 P1_C20457 ( .IN1(P1_N536), .IN2(P1_N530), .Q(P1_N5979) );
  AND2X1 P1_C20458 ( .IN1(n7271), .IN2(n6620), .Q(P1_N5980) );
  AND2X1 P1_C20634 ( .IN1(P1_N536), .IN2(P1_N531), .Q(P1_N6041) );
  AND2X1 P1_C20635 ( .IN1(n7271), .IN2(n6619), .Q(P1_N6042) );
  AND2X1 P1_C20638 ( .IN1(P1_N536), .IN2(P1_N530), .Q(P1_N6043) );
  AND2X1 P1_C20639 ( .IN1(n7271), .IN2(n6620), .Q(P1_N6044) );
  AND2X1 P1_C20809 ( .IN1(P1_N536), .IN2(P1_N531), .Q(P1_N6105) );
  AND2X1 P1_C20810 ( .IN1(n7271), .IN2(n6619), .Q(P1_N6106) );
  AND2X1 P1_C20813 ( .IN1(P1_N536), .IN2(P1_N530), .Q(P1_N6107) );
  AND2X1 P1_C20814 ( .IN1(n7271), .IN2(n6620), .Q(P1_N6108) );
  AND2X1 P1_C20981 ( .IN1(P1_N536), .IN2(P1_N531), .Q(P1_N6169) );
  AND2X1 P1_C20982 ( .IN1(n7271), .IN2(n6619), .Q(P1_N6170) );
  AND2X1 P1_C20985 ( .IN1(P1_N536), .IN2(P1_N530), .Q(P1_N6171) );
  AND2X1 P1_C20986 ( .IN1(n7271), .IN2(n6620), .Q(P1_N6172) );
  AND2X1 P1_C21158 ( .IN1(P1_N536), .IN2(P1_N531), .Q(P1_N6233) );
  AND2X1 P1_C21159 ( .IN1(n7271), .IN2(n6619), .Q(P1_N6234) );
  AND2X1 P1_C21162 ( .IN1(P1_N536), .IN2(P1_N530), .Q(P1_N6235) );
  AND2X1 P1_C21163 ( .IN1(n7271), .IN2(n6620), .Q(P1_N6236) );
  AND2X1 P1_C21338 ( .IN1(P1_N536), .IN2(P1_N531), .Q(P1_N6297) );
  AND2X1 P1_C21339 ( .IN1(n7271), .IN2(n6619), .Q(P1_N6298) );
  AND2X1 P1_C21342 ( .IN1(P1_N536), .IN2(P1_N530), .Q(P1_N6299) );
  AND2X1 P1_C21343 ( .IN1(n7271), .IN2(n6620), .Q(P1_N6300) );
  AND2X1 P1_C21515 ( .IN1(P1_N536), .IN2(P1_N531), .Q(P1_N6361) );
  AND2X1 P1_C21516 ( .IN1(n7271), .IN2(n6619), .Q(P1_N6362) );
  AND2X1 P1_C20073 ( .IN1(n7480), .IN2(n6628), .Q(P1_N5834) );
  OR2X1 P1_C20075 ( .IN2(P1_N5836), .IN1(P1_N5835), .Q(P1_N360) );
  AND2X1 P1_C20076 ( .IN1(n6712), .IN2(P1_N105), .Q(P1_N5835) );
  AND2X1 P1_C20077 ( .IN1(n7480), .IN2(n6627), .Q(P1_N5836) );
  OR2X1 P1_C20079 ( .IN2(P1_N5838), .IN1(P1_N5837), .Q(P1_N361) );
  AND2X1 P1_C20080 ( .IN1(n6704), .IN2(P1_N104), .Q(P1_N5837) );
  AND2X1 P1_C20081 ( .IN1(n6703), .IN2(n6626), .Q(P1_N5838) );
  OR2X1 P1_C20083 ( .IN2(P1_N5840), .IN1(P1_N5839), .Q(P1_N362) );
  AND2X1 P1_C20084 ( .IN1(n6718), .IN2(P1_N103), .Q(P1_N5839) );
  AND2X1 P1_C20085 ( .IN1(n6705), .IN2(n6625), .Q(P1_N5840) );
  OR2X1 P1_C20087 ( .IN2(P1_N5842), .IN1(P1_N5841), .Q(P1_N363) );
  AND2X1 P1_C20088 ( .IN1(n6718), .IN2(n6624), .Q(P1_N5841) );
  AND2X1 P1_C20089 ( .IN1(n6705), .IN2(n6624), .Q(P1_N5842) );
  AND2X1 P1_C20092 ( .IN1(n6706), .IN2(P1_N133), .Q(P1_N395) );
  OR2X1 P1_C20095 ( .IN2(P1_N5846), .IN1(P1_N5845), .Q(P1_N396) );
  AND2X1 P1_C20096 ( .IN1(n6708), .IN2(P1_N132), .Q(P1_N5845) );
  AND2X1 P1_C20097 ( .IN1(n19009), .IN2(n10129), .Q(P1_N5846) );
  OR2X1 P1_C20099 ( .IN2(P1_N5848), .IN1(P1_N5847), .Q(P1_N397) );
  AND2X1 P1_C20100 ( .IN1(n6708), .IN2(P1_N131), .Q(P1_N5847) );
  AND2X1 P1_C20101 ( .IN1(n19009), .IN2(n10125), .Q(P1_N5848) );
  OR2X1 P1_C20103 ( .IN2(P1_N5850), .IN1(P1_N5849), .Q(P1_N398) );
  AND2X1 P1_C20104 ( .IN1(n6708), .IN2(P1_N130), .Q(P1_N5849) );
  AND2X1 P1_C20105 ( .IN1(n19009), .IN2(n10145), .Q(P1_N5850) );
  OR2X1 P1_C20107 ( .IN2(P1_N5852), .IN1(P1_N5851), .Q(P1_N399) );
  AND2X1 P1_C20108 ( .IN1(n6708), .IN2(P1_N129), .Q(P1_N5851) );
  AND2X1 P1_C20109 ( .IN1(n19009), .IN2(n10373), .Q(P1_N5852) );
  OR2X1 P1_C20111 ( .IN2(P1_N5854), .IN1(P1_N5853), .Q(P1_N400) );
  AND2X1 P1_C20112 ( .IN1(n6708), .IN2(P1_N128), .Q(P1_N5853) );
  AND2X1 P1_C20113 ( .IN1(n19009), .IN2(n10187), .Q(P1_N5854) );
  OR2X1 P1_C20115 ( .IN2(P1_N5856), .IN1(P1_N5855), .Q(P1_N401) );
  AND2X1 P1_C20116 ( .IN1(n6706), .IN2(P1_N127), .Q(P1_N5855) );
  AND2X1 P1_C20117 ( .IN1(n6705), .IN2(n10381), .Q(P1_N5856) );
  OR2X1 P1_C20119 ( .IN2(P1_N5858), .IN1(P1_N5857), .Q(P1_N402) );
  AND2X1 P1_C20120 ( .IN1(n6706), .IN2(P1_N126), .Q(P1_N5857) );
  AND2X1 P1_C20121 ( .IN1(n6705), .IN2(n10195), .Q(P1_N5858) );
  OR2X1 P1_C20123 ( .IN2(P1_N5860), .IN1(P1_N5859), .Q(P1_N403) );
  AND2X1 P1_C20124 ( .IN1(n6706), .IN2(P1_N125), .Q(P1_N5859) );
  AND2X1 P1_C20125 ( .IN1(n6705), .IN2(n6637), .Q(P1_N5860) );
  OR2X1 P1_C20127 ( .IN2(P1_N5862), .IN1(P1_N5861), .Q(P1_N404) );
  AND2X1 P1_C20128 ( .IN1(n6706), .IN2(P1_N124), .Q(P1_N5861) );
  AND2X1 P1_C20129 ( .IN1(n6705), .IN2(n6638), .Q(P1_N5862) );
  OR2X1 P1_C20131 ( .IN2(P1_N5864), .IN1(P1_N5863), .Q(P1_N405) );
  AND2X1 P1_C20132 ( .IN1(n6714), .IN2(P1_N123), .Q(P1_N5863) );
  AND2X1 P1_C20133 ( .IN1(n6713), .IN2(n6639), .Q(P1_N5864) );
  OR2X1 P1_C20135 ( .IN2(P1_N5866), .IN1(P1_N5865), .Q(P1_N406) );
  AND2X1 P1_C20136 ( .IN1(n6714), .IN2(P1_N122), .Q(P1_N5865) );
  AND2X1 P1_C20137 ( .IN1(n6713), .IN2(n6640), .Q(P1_N5866) );
  OR2X1 P1_C20139 ( .IN2(P1_N5868), .IN1(P1_N5867), .Q(P1_N407) );
  AND2X1 P1_C20140 ( .IN1(n6714), .IN2(P1_N121), .Q(P1_N5867) );
  AND2X1 P1_C20141 ( .IN1(n6713), .IN2(n6641), .Q(P1_N5868) );
  OR2X1 P1_C20143 ( .IN2(P1_N5870), .IN1(P1_N5869), .Q(P1_N408) );
  AND2X1 P1_C20144 ( .IN1(n6714), .IN2(P1_N120), .Q(P1_N5869) );
  AND2X1 P1_C20145 ( .IN1(n6713), .IN2(n6642), .Q(P1_N5870) );
  OR2X1 P1_C20147 ( .IN2(P1_N5872), .IN1(P1_N5871), .Q(P1_N409) );
  AND2X1 P1_C20148 ( .IN1(n6718), .IN2(P1_N119), .Q(P1_N5871) );
  AND2X1 P1_C20149 ( .IN1(n6705), .IN2(n6643), .Q(P1_N5872) );
  OR2X1 P1_C20151 ( .IN2(P1_N5874), .IN1(P1_N5873), .Q(P1_N410) );
  AND2X1 P1_C20152 ( .IN1(n6718), .IN2(P1_N118), .Q(P1_N5873) );
  AND2X1 P1_C20153 ( .IN1(n6705), .IN2(n6644), .Q(P1_N5874) );
  OR2X1 P1_C20155 ( .IN2(P1_N5876), .IN1(P1_N5875), .Q(P1_N411) );
  AND2X1 P1_C20156 ( .IN1(n6704), .IN2(P1_N117), .Q(P1_N5875) );
  AND2X1 P1_C20157 ( .IN1(n6703), .IN2(n6645), .Q(P1_N5876) );
  OR2X1 P1_C20159 ( .IN2(P1_N5878), .IN1(P1_N5877), .Q(P1_N412) );
  AND2X1 P1_C20160 ( .IN1(n6704), .IN2(P1_N116), .Q(P1_N5877) );
  AND2X1 P1_C20161 ( .IN1(n6703), .IN2(n6646), .Q(P1_N5878) );
  OR2X1 P1_C20163 ( .IN2(P1_N5880), .IN1(P1_N5879), .Q(P1_N413) );
  AND2X1 P1_C20164 ( .IN1(n6716), .IN2(P1_N115), .Q(P1_N5879) );
  AND2X1 P1_C20165 ( .IN1(n6715), .IN2(n6647), .Q(P1_N5880) );
  OR2X1 P1_C20167 ( .IN2(P1_N5882), .IN1(P1_N5881), .Q(P1_N414) );
  AND2X1 P1_C20168 ( .IN1(n6712), .IN2(P1_N114), .Q(P1_N5881) );
  AND2X1 P1_C20169 ( .IN1(n7480), .IN2(n6636), .Q(P1_N5882) );
  OR2X1 P1_C20171 ( .IN2(P1_N5884), .IN1(P1_N5883), .Q(P1_N415) );
  AND2X1 P1_C20172 ( .IN1(n6712), .IN2(P1_N113), .Q(P1_N5883) );
  AND2X1 P1_C20173 ( .IN1(n7480), .IN2(n6635), .Q(P1_N5884) );
  OR2X1 P1_C20175 ( .IN2(P1_N5886), .IN1(P1_N5885), .Q(P1_N416) );
  AND2X1 P1_C20176 ( .IN1(n6710), .IN2(P1_N112), .Q(P1_N5885) );
  AND2X1 P1_C20177 ( .IN1(n19009), .IN2(n6634), .Q(P1_N5886) );
  OR2X1 P1_C20179 ( .IN2(P1_N5888), .IN1(P1_N5887), .Q(P1_N417) );
  AND2X1 P1_C20180 ( .IN1(n6710), .IN2(P1_N111), .Q(P1_N5887) );
  AND2X1 P1_C20181 ( .IN1(n19009), .IN2(n6633), .Q(P1_N5888) );
  OR2X1 P1_C20183 ( .IN2(P1_N5890), .IN1(P1_N5889), .Q(P1_N418) );
  AND2X1 P1_C20184 ( .IN1(n6716), .IN2(P1_N110), .Q(P1_N5889) );
  AND2X1 P1_C20185 ( .IN1(n6715), .IN2(n6632), .Q(P1_N5890) );
  OR2X1 P1_C20187 ( .IN2(P1_N5892), .IN1(P1_N5891), .Q(P1_N419) );
  AND2X1 P1_C20188 ( .IN1(n6716), .IN2(P1_N109), .Q(P1_N5891) );
  AND2X1 P1_C20189 ( .IN1(n6715), .IN2(n6631), .Q(P1_N5892) );
  OR2X1 P1_C20191 ( .IN2(P1_N5894), .IN1(P1_N5893), .Q(P1_N420) );
  AND2X1 P1_C20192 ( .IN1(n6716), .IN2(P1_N108), .Q(P1_N5893) );
  AND2X1 P1_C20193 ( .IN1(n6715), .IN2(n6630), .Q(P1_N5894) );
  OR2X1 P1_C20195 ( .IN2(P1_N5896), .IN1(P1_N5895), .Q(P1_N421) );
  AND2X1 P1_C20196 ( .IN1(n6716), .IN2(P1_N107), .Q(P1_N5895) );
  AND2X1 P1_C20197 ( .IN1(n6715), .IN2(n6629), .Q(P1_N5896) );
  OR2X1 P1_C20199 ( .IN2(P1_N5898), .IN1(P1_N5897), .Q(P1_N422) );
  AND2X1 P1_C19926 ( .IN1(n6705), .IN2(n6645), .Q(P1_N5772) );
  OR2X1 P1_C19928 ( .IN2(P1_N5774), .IN1(P1_N5773), .Q(P1_N305) );
  AND2X1 P1_C19929 ( .IN1(n6704), .IN2(P1_N116), .Q(P1_N5773) );
  AND2X1 P1_C19930 ( .IN1(n6703), .IN2(n6646), .Q(P1_N5774) );
  OR2X1 P1_C19932 ( .IN2(P1_N5776), .IN1(P1_N5775), .Q(P1_N306) );
  AND2X1 P1_C19933 ( .IN1(n6712), .IN2(P1_N115), .Q(P1_N5775) );
  AND2X1 P1_C19934 ( .IN1(n7480), .IN2(n6647), .Q(P1_N5776) );
  OR2X1 P1_C19936 ( .IN2(P1_N5778), .IN1(P1_N5777), .Q(P1_N307) );
  AND2X1 P1_C19937 ( .IN1(n6712), .IN2(P1_N114), .Q(P1_N5777) );
  AND2X1 P1_C19938 ( .IN1(n7480), .IN2(n6636), .Q(P1_N5778) );
  OR2X1 P1_C19940 ( .IN2(P1_N5780), .IN1(P1_N5779), .Q(P1_N308) );
  AND2X1 P1_C19941 ( .IN1(n6712), .IN2(P1_N113), .Q(P1_N5779) );
  AND2X1 P1_C19942 ( .IN1(n7480), .IN2(n6635), .Q(P1_N5780) );
  OR2X1 P1_C19944 ( .IN2(P1_N5782), .IN1(P1_N5781), .Q(P1_N309) );
  AND2X1 P1_C19945 ( .IN1(n6710), .IN2(P1_N112), .Q(P1_N5781) );
  AND2X1 P1_C19946 ( .IN1(n7480), .IN2(n6634), .Q(P1_N5782) );
  OR2X1 P1_C19948 ( .IN2(P1_N5784), .IN1(P1_N5783), .Q(P1_N310) );
  AND2X1 P1_C19949 ( .IN1(n6710), .IN2(P1_N111), .Q(P1_N5783) );
  AND2X1 P1_C19950 ( .IN1(n19009), .IN2(n6633), .Q(P1_N5784) );
  OR2X1 P1_C19952 ( .IN2(P1_N5786), .IN1(P1_N5785), .Q(P1_N311) );
  AND2X1 P1_C19953 ( .IN1(n6710), .IN2(P1_N110), .Q(P1_N5785) );
  AND2X1 P1_C19954 ( .IN1(n19009), .IN2(n6632), .Q(P1_N5786) );
  OR2X1 P1_C19956 ( .IN2(P1_N5788), .IN1(P1_N5787), .Q(P1_N312) );
  AND2X1 P1_C19957 ( .IN1(n6710), .IN2(P1_N109), .Q(P1_N5787) );
  AND2X1 P1_C19958 ( .IN1(n19009), .IN2(n6631), .Q(P1_N5788) );
  OR2X1 P1_C19960 ( .IN2(P1_N5790), .IN1(P1_N5789), .Q(P1_N313) );
  AND2X1 P1_C19961 ( .IN1(n6710), .IN2(P1_N108), .Q(P1_N5789) );
  AND2X1 P1_C19962 ( .IN1(n19009), .IN2(n6630), .Q(P1_N5790) );
  OR2X1 P1_C19964 ( .IN2(P1_N5792), .IN1(P1_N5791), .Q(P1_N314) );
  AND2X1 P1_C19965 ( .IN1(n6716), .IN2(P1_N107), .Q(P1_N5791) );
  AND2X1 P1_C19966 ( .IN1(n6715), .IN2(n6629), .Q(P1_N5792) );
  OR2X1 P1_C19968 ( .IN2(P1_N5794), .IN1(P1_N5793), .Q(P1_N315) );
  AND2X1 P1_C19969 ( .IN1(n6716), .IN2(P1_N106), .Q(P1_N5793) );
  AND2X1 P1_C19970 ( .IN1(n6715), .IN2(n6628), .Q(P1_N5794) );
  OR2X1 P1_C19972 ( .IN2(P1_N5796), .IN1(P1_N5795), .Q(P1_N316) );
  AND2X1 P1_C19973 ( .IN1(n6716), .IN2(P1_N105), .Q(P1_N5795) );
  AND2X1 P1_C19974 ( .IN1(n6715), .IN2(n6627), .Q(P1_N5796) );
  OR2X1 P1_C19976 ( .IN2(P1_N5798), .IN1(P1_N5797), .Q(P1_N317) );
  AND2X1 P1_C19977 ( .IN1(n6704), .IN2(P1_N104), .Q(P1_N5797) );
  AND2X1 P1_C19978 ( .IN1(n6703), .IN2(n6626), .Q(P1_N5798) );
  OR2X1 P1_C19980 ( .IN2(P1_N5800), .IN1(P1_N5799), .Q(P1_N318) );
  AND2X1 P1_C19981 ( .IN1(n6704), .IN2(P1_N103), .Q(P1_N5799) );
  AND2X1 P1_C19982 ( .IN1(n6703), .IN2(n6625), .Q(P1_N5800) );
  OR2X1 P1_C19984 ( .IN2(P1_N5802), .IN1(P1_N5801), .Q(P1_N319) );
  AND2X1 P1_C19985 ( .IN1(n6704), .IN2(n6624), .Q(P1_N5801) );
  AND2X1 P1_C19986 ( .IN1(n6703), .IN2(n6624), .Q(P1_N5802) );
  OR2X1 P1_C20011 ( .IN2(P1_N5804), .IN1(P1_N5803), .Q(P1_N344) );
  AND2X1 P1_C20012 ( .IN1(n6714), .IN2(P1_N121), .Q(P1_N5803) );
  AND2X1 P1_C20013 ( .IN1(n6713), .IN2(n6641), .Q(P1_N5804) );
  OR2X1 P1_C20015 ( .IN2(P1_N5806), .IN1(P1_N5805), .Q(P1_N345) );
  AND2X1 P1_C20016 ( .IN1(n6718), .IN2(P1_N120), .Q(P1_N5805) );
  AND2X1 P1_C20017 ( .IN1(n6713), .IN2(n6642), .Q(P1_N5806) );
  OR2X1 P1_C20019 ( .IN2(P1_N5808), .IN1(P1_N5807), .Q(P1_N346) );
  AND2X1 P1_C20020 ( .IN1(n6718), .IN2(P1_N119), .Q(P1_N5807) );
  AND2X1 P1_C20021 ( .IN1(n6705), .IN2(n6643), .Q(P1_N5808) );
  OR2X1 P1_C20023 ( .IN2(P1_N5810), .IN1(P1_N5809), .Q(P1_N347) );
  AND2X1 P1_C20024 ( .IN1(n6718), .IN2(P1_N118), .Q(P1_N5809) );
  AND2X1 P1_C20025 ( .IN1(n6705), .IN2(n6644), .Q(P1_N5810) );
  OR2X1 P1_C20027 ( .IN2(P1_N5812), .IN1(P1_N5811), .Q(P1_N348) );
  AND2X1 P1_C20028 ( .IN1(n6718), .IN2(P1_N117), .Q(P1_N5811) );
  AND2X1 P1_C20029 ( .IN1(n6705), .IN2(n6645), .Q(P1_N5812) );
  OR2X1 P1_C20031 ( .IN2(P1_N5814), .IN1(P1_N5813), .Q(P1_N349) );
  AND2X1 P1_C20032 ( .IN1(n6712), .IN2(P1_N116), .Q(P1_N5813) );
  AND2X1 P1_C20033 ( .IN1(n7480), .IN2(n6646), .Q(P1_N5814) );
  OR2X1 P1_C20035 ( .IN2(P1_N5816), .IN1(P1_N5815), .Q(P1_N350) );
  AND2X1 P1_C20036 ( .IN1(n6712), .IN2(P1_N115), .Q(P1_N5815) );
  AND2X1 P1_C20037 ( .IN1(n7480), .IN2(n6647), .Q(P1_N5816) );
  OR2X1 P1_C20039 ( .IN2(P1_N5818), .IN1(P1_N5817), .Q(P1_N351) );
  AND2X1 P1_C20040 ( .IN1(n6712), .IN2(P1_N114), .Q(P1_N5817) );
  AND2X1 P1_C20041 ( .IN1(n7480), .IN2(n6636), .Q(P1_N5818) );
  OR2X1 P1_C20043 ( .IN2(P1_N5820), .IN1(P1_N5819), .Q(P1_N352) );
  AND2X1 P1_C20044 ( .IN1(n6712), .IN2(P1_N113), .Q(P1_N5819) );
  AND2X1 P1_C20045 ( .IN1(n7480), .IN2(n6635), .Q(P1_N5820) );
  OR2X1 P1_C20047 ( .IN2(P1_N5822), .IN1(P1_N5821), .Q(P1_N353) );
  AND2X1 P1_C20048 ( .IN1(n6710), .IN2(P1_N112), .Q(P1_N5821) );
  AND2X1 P1_C20049 ( .IN1(n7480), .IN2(n6634), .Q(P1_N5822) );
  OR2X1 P1_C20051 ( .IN2(P1_N5824), .IN1(P1_N5823), .Q(P1_N354) );
  AND2X1 P1_C20052 ( .IN1(n6710), .IN2(P1_N111), .Q(P1_N5823) );
  AND2X1 P1_C20053 ( .IN1(n19009), .IN2(n6633), .Q(P1_N5824) );
  OR2X1 P1_C20055 ( .IN2(P1_N5826), .IN1(P1_N5825), .Q(P1_N355) );
  AND2X1 P1_C20056 ( .IN1(n6710), .IN2(P1_N110), .Q(P1_N5825) );
  AND2X1 P1_C20057 ( .IN1(n19009), .IN2(n6632), .Q(P1_N5826) );
  OR2X1 P1_C20059 ( .IN2(P1_N5828), .IN1(P1_N5827), .Q(P1_N356) );
  AND2X1 P1_C20060 ( .IN1(n6710), .IN2(P1_N109), .Q(P1_N5827) );
  AND2X1 P1_C20061 ( .IN1(n19009), .IN2(n6631), .Q(P1_N5828) );
  OR2X1 P1_C20063 ( .IN2(P1_N5830), .IN1(P1_N5829), .Q(P1_N357) );
  AND2X1 P1_C20064 ( .IN1(n6710), .IN2(P1_N108), .Q(P1_N5829) );
  AND2X1 P1_C20065 ( .IN1(n19009), .IN2(n6630), .Q(P1_N5830) );
  OR2X1 P1_C20067 ( .IN2(P1_N5832), .IN1(P1_N5831), .Q(P1_N358) );
  AND2X1 P1_C20068 ( .IN1(n6710), .IN2(P1_N107), .Q(P1_N5831) );
  AND2X1 P1_C20069 ( .IN1(n19009), .IN2(n6629), .Q(P1_N5832) );
  OR2X1 P1_C20071 ( .IN2(P1_N5834), .IN1(P1_N5833), .Q(P1_N359) );
  AND2X1 P1_C20072 ( .IN1(n6712), .IN2(P1_N106), .Q(P1_N5833) );
  AND2X1 P1_C19782 ( .IN1(n6706), .IN2(P1_N123), .Q(P1_N5709) );
  AND2X1 P1_C19783 ( .IN1(n6705), .IN2(n6639), .Q(P1_N5710) );
  OR2X1 P1_C19785 ( .IN2(P1_N5712), .IN1(P1_N5711), .Q(P1_N251) );
  AND2X1 P1_C19786 ( .IN1(n6714), .IN2(P1_N122), .Q(P1_N5711) );
  AND2X1 P1_C19787 ( .IN1(n6713), .IN2(n6640), .Q(P1_N5712) );
  OR2X1 P1_C19789 ( .IN2(P1_N5714), .IN1(P1_N5713), .Q(P1_N252) );
  AND2X1 P1_C19790 ( .IN1(n6714), .IN2(P1_N121), .Q(P1_N5713) );
  AND2X1 P1_C19791 ( .IN1(n6713), .IN2(n6641), .Q(P1_N5714) );
  OR2X1 P1_C19793 ( .IN2(P1_N5716), .IN1(P1_N5715), .Q(P1_N253) );
  AND2X1 P1_C19794 ( .IN1(n6718), .IN2(P1_N120), .Q(P1_N5715) );
  AND2X1 P1_C19795 ( .IN1(n6705), .IN2(n6642), .Q(P1_N5716) );
  OR2X1 P1_C19797 ( .IN2(P1_N5718), .IN1(P1_N5717), .Q(P1_N254) );
  AND2X1 P1_C19798 ( .IN1(n6718), .IN2(P1_N119), .Q(P1_N5717) );
  AND2X1 P1_C19799 ( .IN1(n6705), .IN2(n6643), .Q(P1_N5718) );
  OR2X1 P1_C19801 ( .IN2(P1_N5720), .IN1(P1_N5719), .Q(P1_N255) );
  AND2X1 P1_C19802 ( .IN1(n6718), .IN2(P1_N118), .Q(P1_N5719) );
  AND2X1 P1_C19803 ( .IN1(n6713), .IN2(n6644), .Q(P1_N5720) );
  OR2X1 P1_C19805 ( .IN2(P1_N5722), .IN1(P1_N5721), .Q(P1_N256) );
  AND2X1 P1_C19806 ( .IN1(n6718), .IN2(P1_N117), .Q(P1_N5721) );
  AND2X1 P1_C19807 ( .IN1(n6705), .IN2(n6645), .Q(P1_N5722) );
  OR2X1 P1_C19809 ( .IN2(P1_N5724), .IN1(P1_N5723), .Q(P1_N257) );
  AND2X1 P1_C19810 ( .IN1(n6712), .IN2(P1_N116), .Q(P1_N5723) );
  AND2X1 P1_C19811 ( .IN1(n7480), .IN2(n6646), .Q(P1_N5724) );
  OR2X1 P1_C19813 ( .IN2(P1_N5726), .IN1(P1_N5725), .Q(P1_N258) );
  AND2X1 P1_C19814 ( .IN1(n6712), .IN2(P1_N115), .Q(P1_N5725) );
  AND2X1 P1_C19815 ( .IN1(n7480), .IN2(n6647), .Q(P1_N5726) );
  OR2X1 P1_C19817 ( .IN2(P1_N5728), .IN1(P1_N5727), .Q(P1_N259) );
  AND2X1 P1_C19818 ( .IN1(n6712), .IN2(P1_N114), .Q(P1_N5727) );
  AND2X1 P1_C19819 ( .IN1(n7480), .IN2(n6636), .Q(P1_N5728) );
  OR2X1 P1_C19821 ( .IN2(P1_N5730), .IN1(P1_N5729), .Q(P1_N260) );
  AND2X1 P1_C19822 ( .IN1(n6712), .IN2(P1_N113), .Q(P1_N5729) );
  AND2X1 P1_C19823 ( .IN1(n7480), .IN2(n6635), .Q(P1_N5730) );
  OR2X1 P1_C19825 ( .IN2(P1_N5732), .IN1(P1_N5731), .Q(P1_N261) );
  AND2X1 P1_C19826 ( .IN1(n6712), .IN2(P1_N112), .Q(P1_N5731) );
  AND2X1 P1_C19827 ( .IN1(n7480), .IN2(n6634), .Q(P1_N5732) );
  OR2X1 P1_C19829 ( .IN2(P1_N5734), .IN1(P1_N5733), .Q(P1_N262) );
  AND2X1 P1_C19830 ( .IN1(n6710), .IN2(P1_N111), .Q(P1_N5733) );
  AND2X1 P1_C19831 ( .IN1(n19009), .IN2(n6633), .Q(P1_N5734) );
  OR2X1 P1_C19833 ( .IN2(P1_N5736), .IN1(P1_N5735), .Q(P1_N263) );
  AND2X1 P1_C19834 ( .IN1(n6710), .IN2(P1_N110), .Q(P1_N5735) );
  AND2X1 P1_C19835 ( .IN1(n19009), .IN2(n6632), .Q(P1_N5736) );
  OR2X1 P1_C19837 ( .IN2(P1_N5738), .IN1(P1_N5737), .Q(P1_N264) );
  AND2X1 P1_C19838 ( .IN1(n6710), .IN2(P1_N109), .Q(P1_N5737) );
  AND2X1 P1_C19839 ( .IN1(n19009), .IN2(n6631), .Q(P1_N5738) );
  OR2X1 P1_C19841 ( .IN2(P1_N5740), .IN1(P1_N5739), .Q(P1_N265) );
  AND2X1 P1_C19842 ( .IN1(n6710), .IN2(P1_N108), .Q(P1_N5739) );
  AND2X1 P1_C19843 ( .IN1(n19009), .IN2(n6630), .Q(P1_N5740) );
  OR2X1 P1_C19845 ( .IN2(P1_N5742), .IN1(P1_N5741), .Q(P1_N266) );
  AND2X1 P1_C19846 ( .IN1(n6710), .IN2(P1_N107), .Q(P1_N5741) );
  AND2X1 P1_C19847 ( .IN1(n19009), .IN2(n6629), .Q(P1_N5742) );
  OR2X1 P1_C19849 ( .IN2(P1_N5744), .IN1(P1_N5743), .Q(P1_N267) );
  AND2X1 P1_C19850 ( .IN1(n6716), .IN2(P1_N106), .Q(P1_N5743) );
  AND2X1 P1_C19851 ( .IN1(n6703), .IN2(n6628), .Q(P1_N5744) );
  OR2X1 P1_C19853 ( .IN2(P1_N5746), .IN1(P1_N5745), .Q(P1_N268) );
  AND2X1 P1_C19854 ( .IN1(n6704), .IN2(P1_N105), .Q(P1_N5745) );
  AND2X1 P1_C19855 ( .IN1(n6703), .IN2(n6627), .Q(P1_N5746) );
  OR2X1 P1_C19857 ( .IN2(P1_N5748), .IN1(P1_N5747), .Q(P1_N269) );
  AND2X1 P1_C19858 ( .IN1(n6704), .IN2(P1_N104), .Q(P1_N5747) );
  AND2X1 P1_C19859 ( .IN1(n6703), .IN2(n6626), .Q(P1_N5748) );
  OR2X1 P1_C19861 ( .IN2(P1_N5750), .IN1(P1_N5749), .Q(P1_N270) );
  AND2X1 P1_C19862 ( .IN1(n6704), .IN2(P1_N103), .Q(P1_N5749) );
  AND2X1 P1_C19863 ( .IN1(n6703), .IN2(n6625), .Q(P1_N5750) );
  OR2X1 P1_C19865 ( .IN2(P1_N5752), .IN1(P1_N5751), .Q(P1_N271) );
  AND2X1 P1_C19866 ( .IN1(n6704), .IN2(n6624), .Q(P1_N5751) );
  AND2X1 P1_C19867 ( .IN1(n6703), .IN2(n6624), .Q(P1_N5752) );
  AND2X1 P1_C19889 ( .IN1(n6706), .IN2(P1_N133), .Q(P1_N295) );
  AND2X1 P1_C19893 ( .IN1(n6706), .IN2(P1_N125), .Q(P1_N5755) );
  AND2X1 P1_C19894 ( .IN1(n6705), .IN2(n6637), .Q(P1_N5756) );
  OR2X1 P1_C19896 ( .IN2(P1_N5758), .IN1(P1_N5757), .Q(P1_N297) );
  AND2X1 P1_C19897 ( .IN1(n6706), .IN2(P1_N124), .Q(P1_N5757) );
  AND2X1 P1_C19898 ( .IN1(n6705), .IN2(n6638), .Q(P1_N5758) );
  OR2X1 P1_C19900 ( .IN2(P1_N5760), .IN1(P1_N5759), .Q(P1_N298) );
  AND2X1 P1_C19901 ( .IN1(n6706), .IN2(P1_N123), .Q(P1_N5759) );
  AND2X1 P1_C19902 ( .IN1(n6705), .IN2(n6639), .Q(P1_N5760) );
  OR2X1 P1_C19904 ( .IN2(P1_N5762), .IN1(P1_N5761), .Q(P1_N299) );
  AND2X1 P1_C19905 ( .IN1(n6714), .IN2(P1_N122), .Q(P1_N5761) );
  AND2X1 P1_C19906 ( .IN1(n6713), .IN2(n6640), .Q(P1_N5762) );
  OR2X1 P1_C19908 ( .IN2(P1_N5764), .IN1(P1_N5763), .Q(P1_N300) );
  AND2X1 P1_C19909 ( .IN1(n6714), .IN2(P1_N121), .Q(P1_N5763) );
  AND2X1 P1_C19910 ( .IN1(n6713), .IN2(n6641), .Q(P1_N5764) );
  OR2X1 P1_C19912 ( .IN2(P1_N5766), .IN1(P1_N5765), .Q(P1_N301) );
  AND2X1 P1_C19913 ( .IN1(n6714), .IN2(P1_N120), .Q(P1_N5765) );
  AND2X1 P1_C19914 ( .IN1(n6705), .IN2(n6642), .Q(P1_N5766) );
  OR2X1 P1_C19916 ( .IN2(P1_N5768), .IN1(P1_N5767), .Q(P1_N302) );
  AND2X1 P1_C19917 ( .IN1(n6718), .IN2(P1_N119), .Q(P1_N5767) );
  AND2X1 P1_C19918 ( .IN1(n6705), .IN2(n6643), .Q(P1_N5768) );
  OR2X1 P1_C19920 ( .IN2(P1_N5770), .IN1(P1_N5769), .Q(P1_N303) );
  AND2X1 P1_C19921 ( .IN1(n6718), .IN2(P1_N118), .Q(P1_N5769) );
  AND2X1 P1_C19922 ( .IN1(n6713), .IN2(n6644), .Q(P1_N5770) );
  OR2X1 P1_C19924 ( .IN2(P1_N5772), .IN1(P1_N5771), .Q(P1_N304) );
  AND2X1 P1_C19925 ( .IN1(n6718), .IN2(P1_N117), .Q(P1_N5771) );
  AND2X1 P1_C19600 ( .IN1(n6703), .IN2(n6626), .Q(P1_N5644) );
  OR2X1 P1_C19602 ( .IN2(P1_N5646), .IN1(P1_N5645), .Q(P1_N162) );
  AND2X1 P1_C19603 ( .IN1(n6704), .IN2(P1_N103), .Q(P1_N5645) );
  AND2X1 P1_C19604 ( .IN1(n6703), .IN2(n6625), .Q(P1_N5646) );
  OR2X1 P1_C19606 ( .IN2(P1_N5648), .IN1(P1_N5647), .Q(P1_N163) );
  AND2X1 P1_C19607 ( .IN1(n6704), .IN2(n6624), .Q(P1_N5647) );
  AND2X1 P1_C19608 ( .IN1(n6703), .IN2(n6624), .Q(P1_N5648) );
  AND2X1 P1_C19638 ( .IN1(n6706), .IN2(P1_N133), .Q(P1_N193) );
  OR2X1 P1_C19641 ( .IN2(P1_N5652), .IN1(P1_N5651), .Q(P1_N194) );
  AND2X1 P1_C19642 ( .IN1(n6708), .IN2(P1_N128), .Q(P1_N5651) );
  AND2X1 P1_C19643 ( .IN1(n19009), .IN2(n10187), .Q(P1_N5652) );
  AND2X1 P1_C19646 ( .IN1(n6708), .IN2(P1_N127), .Q(P1_N5653) );
  AND2X1 P1_C19647 ( .IN1(n19009), .IN2(n10381), .Q(P1_N5654) );
  OR2X1 P1_C19649 ( .IN2(P1_N5656), .IN1(P1_N5655), .Q(P1_N196) );
  AND2X1 P1_C19650 ( .IN1(n6708), .IN2(P1_N126), .Q(P1_N5655) );
  AND2X1 P1_C19651 ( .IN1(n19009), .IN2(n10195), .Q(P1_N5656) );
  OR2X1 P1_C19653 ( .IN2(P1_N5658), .IN1(P1_N5657), .Q(P1_N197) );
  AND2X1 P1_C19654 ( .IN1(n6706), .IN2(P1_N125), .Q(P1_N5657) );
  AND2X1 P1_C19655 ( .IN1(n6705), .IN2(n6637), .Q(P1_N5658) );
  OR2X1 P1_C19657 ( .IN2(P1_N5660), .IN1(P1_N5659), .Q(P1_N198) );
  AND2X1 P1_C19658 ( .IN1(n6706), .IN2(P1_N124), .Q(P1_N5659) );
  AND2X1 P1_C19659 ( .IN1(n6705), .IN2(n6638), .Q(P1_N5660) );
  OR2X1 P1_C19661 ( .IN2(P1_N5662), .IN1(P1_N5661), .Q(P1_N199) );
  AND2X1 P1_C19662 ( .IN1(n6706), .IN2(P1_N123), .Q(P1_N5661) );
  AND2X1 P1_C19663 ( .IN1(n6705), .IN2(n6639), .Q(P1_N5662) );
  OR2X1 P1_C19665 ( .IN2(P1_N5664), .IN1(P1_N5663), .Q(P1_N200) );
  AND2X1 P1_C19666 ( .IN1(n6714), .IN2(P1_N122), .Q(P1_N5663) );
  AND2X1 P1_C19667 ( .IN1(n6713), .IN2(n6640), .Q(P1_N5664) );
  OR2X1 P1_C19669 ( .IN2(P1_N5666), .IN1(P1_N5665), .Q(P1_N201) );
  AND2X1 P1_C19670 ( .IN1(n6714), .IN2(P1_N121), .Q(P1_N5665) );
  AND2X1 P1_C19671 ( .IN1(n6713), .IN2(n6641), .Q(P1_N5666) );
  OR2X1 P1_C19673 ( .IN2(P1_N5668), .IN1(P1_N5667), .Q(P1_N202) );
  AND2X1 P1_C19674 ( .IN1(n6714), .IN2(P1_N120), .Q(P1_N5667) );
  AND2X1 P1_C19675 ( .IN1(n6713), .IN2(n6642), .Q(P1_N5668) );
  OR2X1 P1_C19677 ( .IN2(P1_N5670), .IN1(P1_N5669), .Q(P1_N203) );
  AND2X1 P1_C19678 ( .IN1(n6718), .IN2(P1_N119), .Q(P1_N5669) );
  AND2X1 P1_C19679 ( .IN1(n6705), .IN2(n6643), .Q(P1_N5670) );
  OR2X1 P1_C19681 ( .IN2(P1_N5672), .IN1(P1_N5671), .Q(P1_N204) );
  AND2X1 P1_C19682 ( .IN1(n6718), .IN2(P1_N118), .Q(P1_N5671) );
  AND2X1 P1_C19683 ( .IN1(n6705), .IN2(n6644), .Q(P1_N5672) );
  OR2X1 P1_C19685 ( .IN2(P1_N5674), .IN1(P1_N5673), .Q(P1_N205) );
  AND2X1 P1_C19686 ( .IN1(n6704), .IN2(P1_N117), .Q(P1_N5673) );
  AND2X1 P1_C19687 ( .IN1(n6703), .IN2(n6645), .Q(P1_N5674) );
  OR2X1 P1_C19689 ( .IN2(P1_N5676), .IN1(P1_N5675), .Q(P1_N206) );
  AND2X1 P1_C19690 ( .IN1(n6704), .IN2(P1_N116), .Q(P1_N5675) );
  AND2X1 P1_C19691 ( .IN1(n6703), .IN2(n6646), .Q(P1_N5676) );
  OR2X1 P1_C19693 ( .IN2(P1_N5678), .IN1(P1_N5677), .Q(P1_N207) );
  AND2X1 P1_C19694 ( .IN1(n6716), .IN2(P1_N115), .Q(P1_N5677) );
  AND2X1 P1_C19695 ( .IN1(n6715), .IN2(n6647), .Q(P1_N5678) );
  OR2X1 P1_C19697 ( .IN2(P1_N5680), .IN1(P1_N5679), .Q(P1_N208) );
  AND2X1 P1_C19698 ( .IN1(n6716), .IN2(P1_N114), .Q(P1_N5679) );
  AND2X1 P1_C19699 ( .IN1(n6715), .IN2(n6636), .Q(P1_N5680) );
  OR2X1 P1_C19701 ( .IN2(P1_N5682), .IN1(P1_N5681), .Q(P1_N209) );
  AND2X1 P1_C19702 ( .IN1(n6712), .IN2(P1_N113), .Q(P1_N5681) );
  AND2X1 P1_C19703 ( .IN1(n6715), .IN2(n6635), .Q(P1_N5682) );
  OR2X1 P1_C19705 ( .IN2(P1_N5684), .IN1(P1_N5683), .Q(P1_N210) );
  AND2X1 P1_C19706 ( .IN1(n6716), .IN2(P1_N112), .Q(P1_N5683) );
  AND2X1 P1_C19707 ( .IN1(n6715), .IN2(n6634), .Q(P1_N5684) );
  OR2X1 P1_C19709 ( .IN2(P1_N5686), .IN1(P1_N5685), .Q(P1_N211) );
  AND2X1 P1_C19710 ( .IN1(n6710), .IN2(P1_N111), .Q(P1_N5685) );
  AND2X1 P1_C19711 ( .IN1(n19009), .IN2(n6633), .Q(P1_N5686) );
  OR2X1 P1_C19713 ( .IN2(P1_N5688), .IN1(P1_N5687), .Q(P1_N212) );
  AND2X1 P1_C19714 ( .IN1(n6716), .IN2(P1_N110), .Q(P1_N5687) );
  AND2X1 P1_C19715 ( .IN1(n6715), .IN2(n6632), .Q(P1_N5688) );
  OR2X1 P1_C19717 ( .IN2(P1_N5690), .IN1(P1_N5689), .Q(P1_N213) );
  AND2X1 P1_C19718 ( .IN1(n6716), .IN2(P1_N109), .Q(P1_N5689) );
  AND2X1 P1_C19719 ( .IN1(n6715), .IN2(n6631), .Q(P1_N5690) );
  OR2X1 P1_C19721 ( .IN2(P1_N5692), .IN1(P1_N5691), .Q(P1_N214) );
  AND2X1 P1_C19722 ( .IN1(n6716), .IN2(P1_N108), .Q(P1_N5691) );
  AND2X1 P1_C19723 ( .IN1(n6715), .IN2(n6630), .Q(P1_N5692) );
  OR2X1 P1_C19725 ( .IN2(P1_N5694), .IN1(P1_N5693), .Q(P1_N215) );
  AND2X1 P1_C19726 ( .IN1(n6716), .IN2(P1_N107), .Q(P1_N5693) );
  AND2X1 P1_C19727 ( .IN1(n6715), .IN2(n6629), .Q(P1_N5694) );
  OR2X1 P1_C19729 ( .IN2(P1_N5696), .IN1(P1_N5695), .Q(P1_N216) );
  AND2X1 P1_C19730 ( .IN1(n6716), .IN2(P1_N106), .Q(P1_N5695) );
  AND2X1 P1_C19731 ( .IN1(n6715), .IN2(n6628), .Q(P1_N5696) );
  OR2X1 P1_C19733 ( .IN2(P1_N5698), .IN1(P1_N5697), .Q(P1_N217) );
  AND2X1 P1_C19734 ( .IN1(n6704), .IN2(P1_N105), .Q(P1_N5697) );
  AND2X1 P1_C19735 ( .IN1(n6715), .IN2(n6627), .Q(P1_N5698) );
  OR2X1 P1_C19737 ( .IN2(P1_N5700), .IN1(P1_N5699), .Q(P1_N218) );
  AND2X1 P1_C19738 ( .IN1(n6704), .IN2(P1_N104), .Q(P1_N5699) );
  AND2X1 P1_C19739 ( .IN1(n6703), .IN2(n6626), .Q(P1_N5700) );
  OR2X1 P1_C19741 ( .IN2(P1_N5702), .IN1(P1_N5701), .Q(P1_N219) );
  AND2X1 P1_C19742 ( .IN1(n6704), .IN2(P1_N103), .Q(P1_N5701) );
  AND2X1 P1_C19743 ( .IN1(n6703), .IN2(n6625), .Q(P1_N5702) );
  OR2X1 P1_C19745 ( .IN2(P1_N5704), .IN1(P1_N5703), .Q(P1_N220) );
  AND2X1 P1_C19746 ( .IN1(n6704), .IN2(n6624), .Q(P1_N5703) );
  AND2X1 P1_C19747 ( .IN1(n6703), .IN2(n6624), .Q(P1_N5704) );
  AND2X1 P1_C19774 ( .IN1(n6706), .IN2(P1_N133), .Q(P1_N248) );
  OR2X1 P1_C19777 ( .IN2(P1_N5708), .IN1(P1_N5707), .Q(P1_N249) );
  AND2X1 P1_C19778 ( .IN1(n6706), .IN2(P1_N124), .Q(P1_N5707) );
  AND2X1 P1_C19779 ( .IN1(n6705), .IN2(n6638), .Q(P1_N5708) );
  OR2X1 P2_C22593 ( .IN2(n6591), .IN1(P2_N6610), .Q(P2_N5354) );
  AND2X1 P1_C1092 ( .IN1(n6980), .IN2(n6958), .Q(P1_N541) );
  AND2X1 P1_C1093 ( .IN1(n6882), .IN2(n6856), .Q(P1_N542) );
  OR2X1 P1_C16110 ( .IN2(n6996), .IN1(P1_N583), .Q(P1_N5570) );
  OR2X1 P1_C16112 ( .IN2(n7340), .IN1(n7337), .Q(P1_N5571) );
  AND2X1 P1_C19491 ( .IN1(n6706), .IN2(P1_N133), .Q(P1_N134) );
  OR2X1 P1_C19494 ( .IN2(P1_N5592), .IN1(P1_N5591), .Q(P1_N135) );
  AND2X1 P1_C19495 ( .IN1(n6708), .IN2(P1_N130), .Q(P1_N5591) );
  AND2X1 P1_C19496 ( .IN1(n19009), .IN2(n10145), .Q(P1_N5592) );
  OR2X1 P1_C19498 ( .IN2(P1_N5594), .IN1(P1_N5593), .Q(P1_N136) );
  AND2X1 P1_C19499 ( .IN1(n6708), .IN2(P1_N129), .Q(P1_N5593) );
  AND2X1 P1_C19500 ( .IN1(n19009), .IN2(n10373), .Q(P1_N5594) );
  OR2X1 P1_C19502 ( .IN2(P1_N5596), .IN1(P1_N5595), .Q(P1_N137) );
  AND2X1 P1_C19503 ( .IN1(n6708), .IN2(P1_N128), .Q(P1_N5595) );
  AND2X1 P1_C19504 ( .IN1(n19009), .IN2(n10187), .Q(P1_N5596) );
  OR2X1 P1_C19506 ( .IN2(P1_N5598), .IN1(P1_N5597), .Q(P1_N138) );
  AND2X1 P1_C19507 ( .IN1(n6706), .IN2(P1_N127), .Q(P1_N5597) );
  AND2X1 P1_C19508 ( .IN1(n6705), .IN2(n10381), .Q(P1_N5598) );
  OR2X1 P1_C19510 ( .IN2(P1_N5600), .IN1(P1_N5599), .Q(P1_N139) );
  AND2X1 P1_C19511 ( .IN1(n6706), .IN2(P1_N126), .Q(P1_N5599) );
  AND2X1 P1_C19512 ( .IN1(n19009), .IN2(n10195), .Q(P1_N5600) );
  OR2X1 P1_C19514 ( .IN2(P1_N5602), .IN1(P1_N5601), .Q(P1_N140) );
  AND2X1 P1_C19515 ( .IN1(n6706), .IN2(P1_N125), .Q(P1_N5601) );
  AND2X1 P1_C19516 ( .IN1(n6705), .IN2(n6637), .Q(P1_N5602) );
  OR2X1 P1_C19518 ( .IN2(P1_N5604), .IN1(P1_N5603), .Q(P1_N141) );
  AND2X1 P1_C19519 ( .IN1(n6706), .IN2(P1_N124), .Q(P1_N5603) );
  AND2X1 P1_C19520 ( .IN1(n6705), .IN2(n6638), .Q(P1_N5604) );
  OR2X1 P1_C19522 ( .IN2(P1_N5606), .IN1(P1_N5605), .Q(P1_N142) );
  AND2X1 P1_C19523 ( .IN1(n6706), .IN2(P1_N123), .Q(P1_N5605) );
  AND2X1 P1_C19524 ( .IN1(n6705), .IN2(n6639), .Q(P1_N5606) );
  OR2X1 P1_C19526 ( .IN2(P1_N5608), .IN1(P1_N5607), .Q(P1_N143) );
  AND2X1 P1_C19527 ( .IN1(n6714), .IN2(P1_N122), .Q(P1_N5607) );
  AND2X1 P1_C19528 ( .IN1(n6713), .IN2(n6640), .Q(P1_N5608) );
  OR2X1 P1_C19530 ( .IN2(P1_N5610), .IN1(P1_N5609), .Q(P1_N144) );
  AND2X1 P1_C19531 ( .IN1(n6714), .IN2(P1_N121), .Q(P1_N5609) );
  AND2X1 P1_C19532 ( .IN1(n6713), .IN2(n6641), .Q(P1_N5610) );
  OR2X1 P1_C19534 ( .IN2(P1_N5612), .IN1(P1_N5611), .Q(P1_N145) );
  AND2X1 P1_C19535 ( .IN1(n6714), .IN2(P1_N120), .Q(P1_N5611) );
  AND2X1 P1_C19536 ( .IN1(n6713), .IN2(n6642), .Q(P1_N5612) );
  OR2X1 P1_C19538 ( .IN2(P1_N5614), .IN1(P1_N5613), .Q(P1_N146) );
  AND2X1 P1_C19539 ( .IN1(n6718), .IN2(P1_N119), .Q(P1_N5613) );
  AND2X1 P1_C19540 ( .IN1(n6705), .IN2(n6643), .Q(P1_N5614) );
  OR2X1 P1_C19542 ( .IN2(P1_N5616), .IN1(P1_N5615), .Q(P1_N147) );
  AND2X1 P1_C19543 ( .IN1(n6718), .IN2(P1_N118), .Q(P1_N5615) );
  AND2X1 P1_C19544 ( .IN1(n6705), .IN2(n6644), .Q(P1_N5616) );
  OR2X1 P1_C19546 ( .IN2(P1_N5618), .IN1(P1_N5617), .Q(P1_N148) );
  AND2X1 P1_C19547 ( .IN1(n6704), .IN2(P1_N117), .Q(P1_N5617) );
  AND2X1 P1_C19548 ( .IN1(n6703), .IN2(n6645), .Q(P1_N5618) );
  OR2X1 P1_C19550 ( .IN2(P1_N5620), .IN1(P1_N5619), .Q(P1_N149) );
  AND2X1 P1_C19551 ( .IN1(n6704), .IN2(P1_N116), .Q(P1_N5619) );
  AND2X1 P1_C19552 ( .IN1(n6703), .IN2(n6646), .Q(P1_N5620) );
  OR2X1 P1_C19554 ( .IN2(P1_N5622), .IN1(P1_N5621), .Q(P1_N150) );
  AND2X1 P1_C19555 ( .IN1(n6716), .IN2(P1_N115), .Q(P1_N5621) );
  AND2X1 P1_C19556 ( .IN1(n6715), .IN2(n6647), .Q(P1_N5622) );
  OR2X1 P1_C19558 ( .IN2(P1_N5624), .IN1(P1_N5623), .Q(P1_N151) );
  AND2X1 P1_C19559 ( .IN1(n6716), .IN2(P1_N114), .Q(P1_N5623) );
  AND2X1 P1_C19560 ( .IN1(n6715), .IN2(n6636), .Q(P1_N5624) );
  OR2X1 P1_C19562 ( .IN2(P1_N5626), .IN1(P1_N5625), .Q(P1_N152) );
  AND2X1 P1_C19563 ( .IN1(n6712), .IN2(P1_N113), .Q(P1_N5625) );
  AND2X1 P1_C19564 ( .IN1(n6715), .IN2(n6635), .Q(P1_N5626) );
  OR2X1 P1_C19566 ( .IN2(P1_N5628), .IN1(P1_N5627), .Q(P1_N153) );
  AND2X1 P1_C19567 ( .IN1(n6716), .IN2(P1_N112), .Q(P1_N5627) );
  AND2X1 P1_C19568 ( .IN1(n6715), .IN2(n6634), .Q(P1_N5628) );
  OR2X1 P1_C19570 ( .IN2(P1_N5630), .IN1(P1_N5629), .Q(P1_N154) );
  AND2X1 P1_C19571 ( .IN1(n6716), .IN2(P1_N111), .Q(P1_N5629) );
  AND2X1 P1_C19572 ( .IN1(n6715), .IN2(n6633), .Q(P1_N5630) );
  OR2X1 P1_C19574 ( .IN2(P1_N5632), .IN1(P1_N5631), .Q(P1_N155) );
  AND2X1 P1_C19575 ( .IN1(n6716), .IN2(P1_N110), .Q(P1_N5631) );
  AND2X1 P1_C19576 ( .IN1(n6715), .IN2(n6632), .Q(P1_N5632) );
  OR2X1 P1_C19578 ( .IN2(P1_N5634), .IN1(P1_N5633), .Q(P1_N156) );
  AND2X1 P1_C19579 ( .IN1(n6716), .IN2(P1_N109), .Q(P1_N5633) );
  AND2X1 P1_C19580 ( .IN1(n6715), .IN2(n6631), .Q(P1_N5634) );
  OR2X1 P1_C19582 ( .IN2(P1_N5636), .IN1(P1_N5635), .Q(P1_N157) );
  AND2X1 P1_C19583 ( .IN1(n6716), .IN2(P1_N108), .Q(P1_N5635) );
  AND2X1 P1_C19584 ( .IN1(n6715), .IN2(n6630), .Q(P1_N5636) );
  OR2X1 P1_C19586 ( .IN2(P1_N5638), .IN1(P1_N5637), .Q(P1_N158) );
  AND2X1 P1_C19587 ( .IN1(n6716), .IN2(P1_N107), .Q(P1_N5637) );
  AND2X1 P1_C19588 ( .IN1(n6715), .IN2(n6629), .Q(P1_N5638) );
  OR2X1 P1_C19590 ( .IN2(P1_N5640), .IN1(P1_N5639), .Q(P1_N159) );
  AND2X1 P1_C19591 ( .IN1(n6716), .IN2(P1_N106), .Q(P1_N5639) );
  AND2X1 P1_C19592 ( .IN1(n6715), .IN2(n6628), .Q(P1_N5640) );
  OR2X1 P1_C19594 ( .IN2(P1_N5642), .IN1(P1_N5641), .Q(P1_N160) );
  AND2X1 P1_C19595 ( .IN1(n6704), .IN2(P1_N105), .Q(P1_N5641) );
  AND2X1 P1_C19596 ( .IN1(n6703), .IN2(n6627), .Q(P1_N5642) );
  OR2X1 P1_C19598 ( .IN2(P1_N5644), .IN1(P1_N5643), .Q(P1_N161) );
  AND2X1 P1_C19599 ( .IN1(n6704), .IN2(P1_N104), .Q(P1_N5643) );
  AND2X1 P2_C21207 ( .IN1(P2_N536), .IN2(P2_N531), .Q(P2_N6155) );
  AND2X1 P2_C21208 ( .IN1(n7272), .IN2(n6592), .Q(P2_N6156) );
  AND2X1 P2_C21211 ( .IN1(P2_N536), .IN2(P2_N530), .Q(P2_N6157) );
  AND2X1 P2_C21212 ( .IN1(n7272), .IN2(n6593), .Q(P2_N6158) );
  AND2X1 P2_C21387 ( .IN1(P2_N536), .IN2(P2_N531), .Q(P2_N6219) );
  AND2X1 P2_C21388 ( .IN1(n7272), .IN2(n6592), .Q(P2_N6220) );
  AND2X1 P2_C21391 ( .IN1(P2_N536), .IN2(P2_N530), .Q(P2_N6221) );
  AND2X1 P2_C21392 ( .IN1(n7272), .IN2(n6593), .Q(P2_N6222) );
  AND2X1 P2_C21564 ( .IN1(P2_N536), .IN2(P2_N531), .Q(P2_N6283) );
  AND2X1 P2_C21565 ( .IN1(n7272), .IN2(n6592), .Q(P2_N6284) );
  AND2X1 P2_C21568 ( .IN1(P2_N536), .IN2(P2_N530), .Q(P2_N6285) );
  AND2X1 P2_C21569 ( .IN1(n7272), .IN2(n6593), .Q(P2_N6286) );
  AND2X1 P2_C21741 ( .IN1(P2_N536), .IN2(P2_N531), .Q(P2_N6347) );
  AND2X1 P2_C21742 ( .IN1(n7272), .IN2(n6592), .Q(P2_N6348) );
  AND2X1 P2_C21745 ( .IN1(P2_N536), .IN2(P2_N530), .Q(P2_N6349) );
  AND2X1 P2_C21746 ( .IN1(n7272), .IN2(n6593), .Q(P2_N6350) );
  AND2X1 P2_C21921 ( .IN1(P2_N536), .IN2(P2_N531), .Q(P2_N6411) );
  AND2X1 P2_C21922 ( .IN1(n7272), .IN2(n6592), .Q(P2_N6412) );
  AND2X1 P2_C21925 ( .IN1(P2_N536), .IN2(P2_N530), .Q(P2_N6413) );
  AND2X1 P2_C21926 ( .IN1(n7272), .IN2(n6593), .Q(P2_N6414) );
  AND2X1 P2_C22098 ( .IN1(P2_N536), .IN2(P2_N531), .Q(P2_N6475) );
  AND2X1 P2_C22099 ( .IN1(n7272), .IN2(n6592), .Q(P2_N6476) );
  AND2X1 P2_C22102 ( .IN1(P2_N536), .IN2(P2_N530), .Q(P2_N6477) );
  AND2X1 P2_C22103 ( .IN1(n7272), .IN2(n6593), .Q(P2_N6478) );
  OR2X1 P2_C22274 ( .IN2(P2_N6540), .IN1(P2_N6539), .Q(P2_N4178) );
  AND2X1 P2_C22275 ( .IN1(P2_N536), .IN2(P2_N531), .Q(P2_N6539) );
  AND2X1 P2_C22276 ( .IN1(n7272), .IN2(n6592), .Q(P2_N6540) );
  AND2X1 P2_C22279 ( .IN1(P2_N536), .IN2(P2_N530), .Q(P2_N6541) );
  AND2X1 P2_C22280 ( .IN1(n7272), .IN2(n6593), .Q(P2_N6542) );
  OR2X1 P2_C22458 ( .IN2(P2_N6604), .IN1(P2_N6603), .Q(P2_N4561) );
  AND2X1 P2_C22459 ( .IN1(P2_N536), .IN2(P2_N531), .Q(P2_N6603) );
  AND2X1 P2_C22460 ( .IN1(n7272), .IN2(n6592), .Q(P2_N6604) );
  AND2X1 P2_C22463 ( .IN1(P2_N536), .IN2(P2_N530), .Q(P2_N6605) );
  AND2X1 P2_C22464 ( .IN1(n7272), .IN2(n6593), .Q(P2_N6606) );
  OR2X1 P2_C22563 ( .IN2(n6591), .IN1(P2_N5059), .Q(P2_N5206) );
  OR2X1 P2_C22566 ( .IN2(n6591), .IN1(P2_N6607), .Q(P2_N5208) );
  OR2X1 P2_C22570 ( .IN2(n6591), .IN1(P2_N5062), .Q(P2_N5210) );
  OR2X1 P2_C22573 ( .IN2(n6591), .IN1(P2_N6608), .Q(P2_N5212) );
  OR2X1 P2_C22577 ( .IN2(n6591), .IN1(n17734), .Q(P2_N5214) );
  OR2X1 P2_C22581 ( .IN2(n6591), .IN1(P2_N5065), .Q(P2_N5216) );
  OR2X1 P2_C22587 ( .IN2(n6591), .IN1(P2_N5284), .Q(P2_N5285) );
  AND2X1 P2_C20222 ( .IN1(n6694), .IN2(P2_N114), .Q(P2_N5803) );
  AND2X1 P2_C20223 ( .IN1(n6693), .IN2(n6607), .Q(P2_N5804) );
  OR2X1 P2_C20225 ( .IN2(P2_N5806), .IN1(P2_N5805), .Q(P2_N415) );
  AND2X1 P2_C20226 ( .IN1(n6694), .IN2(P2_N113), .Q(P2_N5805) );
  AND2X1 P2_C20227 ( .IN1(n7479), .IN2(n6606), .Q(P2_N5806) );
  OR2X1 P2_C20229 ( .IN2(P2_N5808), .IN1(P2_N5807), .Q(P2_N416) );
  AND2X1 P2_C20230 ( .IN1(n6698), .IN2(P2_N112), .Q(P2_N5807) );
  AND2X1 P2_C20231 ( .IN1(n7479), .IN2(n6605), .Q(P2_N5808) );
  OR2X1 P2_C20233 ( .IN2(P2_N5810), .IN1(P2_N5809), .Q(P2_N417) );
  AND2X1 P2_C20234 ( .IN1(n6698), .IN2(P2_N111), .Q(P2_N5809) );
  AND2X1 P2_C20235 ( .IN1(n6685), .IN2(n6604), .Q(P2_N5810) );
  OR2X1 P2_C20237 ( .IN2(P2_N5812), .IN1(P2_N5811), .Q(P2_N418) );
  AND2X1 P2_C20238 ( .IN1(n6686), .IN2(P2_N110), .Q(P2_N5811) );
  AND2X1 P2_C20239 ( .IN1(n6685), .IN2(n6603), .Q(P2_N5812) );
  OR2X1 P2_C20241 ( .IN2(P2_N5814), .IN1(P2_N5813), .Q(P2_N419) );
  AND2X1 P2_C20242 ( .IN1(n6686), .IN2(P2_N109), .Q(P2_N5813) );
  AND2X1 P2_C20243 ( .IN1(n6685), .IN2(n6602), .Q(P2_N5814) );
  OR2X1 P2_C20245 ( .IN2(P2_N5816), .IN1(P2_N5815), .Q(P2_N420) );
  AND2X1 P2_C20246 ( .IN1(n6686), .IN2(P2_N108), .Q(P2_N5815) );
  AND2X1 P2_C20247 ( .IN1(n6699), .IN2(n6601), .Q(P2_N5816) );
  OR2X1 P2_C20249 ( .IN2(P2_N5818), .IN1(P2_N5817), .Q(P2_N421) );
  AND2X1 P2_C20250 ( .IN1(n6700), .IN2(P2_N107), .Q(P2_N5817) );
  AND2X1 P2_C20251 ( .IN1(n6699), .IN2(n6600), .Q(P2_N5818) );
  OR2X1 P2_C20253 ( .IN2(P2_N5820), .IN1(P2_N5819), .Q(P2_N422) );
  AND2X1 P2_C20254 ( .IN1(n6700), .IN2(P2_N106), .Q(P2_N5819) );
  AND2X1 P2_C20255 ( .IN1(n6699), .IN2(n6599), .Q(P2_N5820) );
  OR2X1 P2_C20257 ( .IN2(P2_N5822), .IN1(P2_N5821), .Q(P2_N423) );
  AND2X1 P2_C20258 ( .IN1(n6700), .IN2(P2_N105), .Q(P2_N5821) );
  AND2X1 P2_C20259 ( .IN1(n6699), .IN2(n6598), .Q(P2_N5822) );
  OR2X1 P2_C20261 ( .IN2(P2_N5824), .IN1(P2_N5823), .Q(P2_N424) );
  AND2X1 P2_C20262 ( .IN1(n6702), .IN2(P2_N104), .Q(P2_N5823) );
  AND2X1 P2_C20263 ( .IN1(n19025), .IN2(n6597), .Q(P2_N5824) );
  OR2X1 P2_C20265 ( .IN2(P2_N5826), .IN1(P2_N5825), .Q(P2_N425) );
  AND2X1 P2_C20266 ( .IN1(n6702), .IN2(P2_N103), .Q(P2_N5825) );
  AND2X1 P2_C20267 ( .IN1(n19025), .IN2(n6596), .Q(P2_N5826) );
  OR2X1 P2_C20269 ( .IN2(P2_N5828), .IN1(P2_N5827), .Q(P2_N426) );
  AND2X1 P2_C20270 ( .IN1(n6692), .IN2(n6595), .Q(P2_N5827) );
  AND2X1 P2_C20271 ( .IN1(n7479), .IN2(n6595), .Q(P2_N5828) );
  AND2X1 P2_C20507 ( .IN1(P2_N536), .IN2(P2_N531), .Q(P2_N5899) );
  AND2X1 P2_C20508 ( .IN1(n7272), .IN2(n6592), .Q(P2_N5900) );
  AND2X1 P2_C20511 ( .IN1(P2_N536), .IN2(P2_N530), .Q(P2_N5901) );
  AND2X1 P2_C20512 ( .IN1(n7272), .IN2(n6593), .Q(P2_N5902) );
  AND2X1 P2_C20683 ( .IN1(P2_N536), .IN2(P2_N531), .Q(P2_N5963) );
  AND2X1 P2_C20684 ( .IN1(n7272), .IN2(n6592), .Q(P2_N5964) );
  AND2X1 P2_C20687 ( .IN1(P2_N536), .IN2(P2_N530), .Q(P2_N5965) );
  AND2X1 P2_C20688 ( .IN1(n7272), .IN2(n6593), .Q(P2_N5966) );
  AND2X1 P2_C20858 ( .IN1(P2_N536), .IN2(P2_N531), .Q(P2_N6027) );
  AND2X1 P2_C20859 ( .IN1(n7272), .IN2(n6592), .Q(P2_N6028) );
  AND2X1 P2_C20862 ( .IN1(P2_N536), .IN2(P2_N530), .Q(P2_N6029) );
  AND2X1 P2_C20863 ( .IN1(n7272), .IN2(n6593), .Q(P2_N6030) );
  AND2X1 P2_C21030 ( .IN1(P2_N536), .IN2(P2_N531), .Q(P2_N6091) );
  AND2X1 P2_C21031 ( .IN1(n7272), .IN2(n6592), .Q(P2_N6092) );
  AND2X1 P2_C21034 ( .IN1(P2_N536), .IN2(P2_N530), .Q(P2_N6093) );
  AND2X1 P2_C21035 ( .IN1(n7272), .IN2(n6593), .Q(P2_N6094) );
  AND2X1 P2_C20095 ( .IN1(n6693), .IN2(n6607), .Q(P2_N5740) );
  OR2X1 P2_C20097 ( .IN2(P2_N5742), .IN1(P2_N5741), .Q(P2_N352) );
  AND2X1 P2_C20098 ( .IN1(n6694), .IN2(P2_N113), .Q(P2_N5741) );
  AND2X1 P2_C20099 ( .IN1(n6693), .IN2(n6606), .Q(P2_N5742) );
  OR2X1 P2_C20101 ( .IN2(P2_N5744), .IN1(P2_N5743), .Q(P2_N353) );
  AND2X1 P2_C20102 ( .IN1(n6698), .IN2(P2_N112), .Q(P2_N5743) );
  AND2X1 P2_C20103 ( .IN1(n7479), .IN2(n6605), .Q(P2_N5744) );
  OR2X1 P2_C20105 ( .IN2(P2_N5746), .IN1(P2_N5745), .Q(P2_N354) );
  AND2X1 P2_C20106 ( .IN1(n6698), .IN2(P2_N111), .Q(P2_N5745) );
  AND2X1 P2_C20107 ( .IN1(n7479), .IN2(n6604), .Q(P2_N5746) );
  OR2X1 P2_C20109 ( .IN2(P2_N5748), .IN1(P2_N5747), .Q(P2_N355) );
  AND2X1 P2_C20110 ( .IN1(n6686), .IN2(P2_N110), .Q(P2_N5747) );
  AND2X1 P2_C20111 ( .IN1(n6685), .IN2(n6603), .Q(P2_N5748) );
  OR2X1 P2_C20113 ( .IN2(P2_N5750), .IN1(P2_N5749), .Q(P2_N356) );
  AND2X1 P2_C20114 ( .IN1(n6686), .IN2(P2_N109), .Q(P2_N5749) );
  AND2X1 P2_C20115 ( .IN1(n6685), .IN2(n6602), .Q(P2_N5750) );
  OR2X1 P2_C20117 ( .IN2(P2_N5752), .IN1(P2_N5751), .Q(P2_N357) );
  AND2X1 P2_C20118 ( .IN1(n6700), .IN2(P2_N108), .Q(P2_N5751) );
  AND2X1 P2_C20119 ( .IN1(n6699), .IN2(n6601), .Q(P2_N5752) );
  OR2X1 P2_C20121 ( .IN2(P2_N5754), .IN1(P2_N5753), .Q(P2_N358) );
  AND2X1 P2_C20122 ( .IN1(n6700), .IN2(P2_N107), .Q(P2_N5753) );
  AND2X1 P2_C20123 ( .IN1(n7479), .IN2(n6600), .Q(P2_N5754) );
  OR2X1 P2_C20125 ( .IN2(P2_N5756), .IN1(P2_N5755), .Q(P2_N359) );
  AND2X1 P2_C20126 ( .IN1(n6700), .IN2(P2_N106), .Q(P2_N5755) );
  AND2X1 P2_C20127 ( .IN1(n6699), .IN2(n6599), .Q(P2_N5756) );
  OR2X1 P2_C20129 ( .IN2(P2_N5758), .IN1(P2_N5757), .Q(P2_N360) );
  AND2X1 P2_C20130 ( .IN1(n6702), .IN2(P2_N105), .Q(P2_N5757) );
  AND2X1 P2_C20131 ( .IN1(n7479), .IN2(n6598), .Q(P2_N5758) );
  OR2X1 P2_C20133 ( .IN2(P2_N5760), .IN1(P2_N5759), .Q(P2_N361) );
  AND2X1 P2_C20134 ( .IN1(n6690), .IN2(P2_N104), .Q(P2_N5759) );
  AND2X1 P2_C20135 ( .IN1(n19025), .IN2(n6597), .Q(P2_N5760) );
  OR2X1 P2_C20137 ( .IN2(P2_N5762), .IN1(P2_N5761), .Q(P2_N362) );
  AND2X1 P2_C20138 ( .IN1(n6690), .IN2(P2_N103), .Q(P2_N5761) );
  AND2X1 P2_C20139 ( .IN1(n19025), .IN2(n6596), .Q(P2_N5762) );
  OR2X1 P2_C20141 ( .IN2(P2_N5764), .IN1(P2_N5763), .Q(P2_N363) );
  AND2X1 P2_C20142 ( .IN1(n6690), .IN2(n6595), .Q(P2_N5763) );
  AND2X1 P2_C20143 ( .IN1(n19025), .IN2(n6595), .Q(P2_N5764) );
  AND2X1 P2_C20146 ( .IN1(n6688), .IN2(P2_N133), .Q(P2_N395) );
  OR2X1 P2_C20149 ( .IN2(P2_N5768), .IN1(P2_N5767), .Q(P2_N396) );
  AND2X1 P2_C20150 ( .IN1(n6688), .IN2(P2_N132), .Q(P2_N5767) );
  AND2X1 P2_C20151 ( .IN1(n6687), .IN2(n10137), .Q(P2_N5768) );
  OR2X1 P2_C20153 ( .IN2(P2_N5770), .IN1(P2_N5769), .Q(P2_N397) );
  AND2X1 P2_C20154 ( .IN1(n6688), .IN2(P2_N131), .Q(P2_N5769) );
  AND2X1 P2_C20155 ( .IN1(n6687), .IN2(n10133), .Q(P2_N5770) );
  OR2X1 P2_C20157 ( .IN2(P2_N5772), .IN1(P2_N5771), .Q(P2_N398) );
  AND2X1 P2_C20158 ( .IN1(n6688), .IN2(P2_N130), .Q(P2_N5771) );
  AND2X1 P2_C20159 ( .IN1(n6687), .IN2(n10141), .Q(P2_N5772) );
  OR2X1 P2_C20161 ( .IN2(P2_N5774), .IN1(P2_N5773), .Q(P2_N399) );
  AND2X1 P2_C20162 ( .IN1(n6688), .IN2(P2_N129), .Q(P2_N5773) );
  AND2X1 P2_C20163 ( .IN1(n6687), .IN2(n10369), .Q(P2_N5774) );
  OR2X1 P2_C20165 ( .IN2(P2_N5776), .IN1(P2_N5775), .Q(P2_N400) );
  AND2X1 P2_C20166 ( .IN1(n6688), .IN2(P2_N128), .Q(P2_N5775) );
  AND2X1 P2_C20167 ( .IN1(n6687), .IN2(n10183), .Q(P2_N5776) );
  OR2X1 P2_C20169 ( .IN2(P2_N5778), .IN1(P2_N5777), .Q(P2_N401) );
  AND2X1 P2_C20170 ( .IN1(n6688), .IN2(P2_N127), .Q(P2_N5777) );
  AND2X1 P2_C20171 ( .IN1(n6687), .IN2(n10377), .Q(P2_N5778) );
  OR2X1 P2_C20173 ( .IN2(P2_N5780), .IN1(P2_N5779), .Q(P2_N402) );
  AND2X1 P2_C20174 ( .IN1(n6688), .IN2(P2_N126), .Q(P2_N5779) );
  AND2X1 P2_C20175 ( .IN1(n6687), .IN2(n10191), .Q(P2_N5780) );
  OR2X1 P2_C20177 ( .IN2(P2_N5782), .IN1(P2_N5781), .Q(P2_N403) );
  AND2X1 P2_C20178 ( .IN1(n6688), .IN2(P2_N125), .Q(P2_N5781) );
  AND2X1 P2_C20179 ( .IN1(n6687), .IN2(n6719), .Q(P2_N5782) );
  OR2X1 P2_C20181 ( .IN2(P2_N5784), .IN1(P2_N5783), .Q(P2_N404) );
  AND2X1 P2_C20182 ( .IN1(n6690), .IN2(P2_N124), .Q(P2_N5783) );
  AND2X1 P2_C20183 ( .IN1(n19025), .IN2(n6608), .Q(P2_N5784) );
  OR2X1 P2_C20185 ( .IN2(P2_N5786), .IN1(P2_N5785), .Q(P2_N405) );
  AND2X1 P2_C20186 ( .IN1(n6690), .IN2(P2_N123), .Q(P2_N5785) );
  AND2X1 P2_C20187 ( .IN1(n19025), .IN2(n6609), .Q(P2_N5786) );
  OR2X1 P2_C20189 ( .IN2(P2_N5788), .IN1(P2_N5787), .Q(P2_N406) );
  AND2X1 P2_C20190 ( .IN1(n6696), .IN2(P2_N122), .Q(P2_N5787) );
  AND2X1 P2_C20191 ( .IN1(n19025), .IN2(n6610), .Q(P2_N5788) );
  OR2X1 P2_C20193 ( .IN2(P2_N5790), .IN1(P2_N5789), .Q(P2_N407) );
  AND2X1 P2_C20194 ( .IN1(n6696), .IN2(P2_N121), .Q(P2_N5789) );
  AND2X1 P2_C20195 ( .IN1(n19025), .IN2(n6611), .Q(P2_N5790) );
  OR2X1 P2_C20197 ( .IN2(P2_N5792), .IN1(P2_N5791), .Q(P2_N408) );
  AND2X1 P2_C20198 ( .IN1(n6696), .IN2(P2_N120), .Q(P2_N5791) );
  AND2X1 P2_C20199 ( .IN1(n6687), .IN2(n6612), .Q(P2_N5792) );
  OR2X1 P2_C20201 ( .IN2(P2_N5794), .IN1(P2_N5793), .Q(P2_N409) );
  AND2X1 P2_C20202 ( .IN1(n6692), .IN2(P2_N119), .Q(P2_N5793) );
  AND2X1 P2_C20203 ( .IN1(n7479), .IN2(n6613), .Q(P2_N5794) );
  OR2X1 P2_C20205 ( .IN2(P2_N5796), .IN1(P2_N5795), .Q(P2_N410) );
  AND2X1 P2_C20206 ( .IN1(n6692), .IN2(P2_N118), .Q(P2_N5795) );
  AND2X1 P2_C20207 ( .IN1(n7479), .IN2(n6614), .Q(P2_N5796) );
  OR2X1 P2_C20209 ( .IN2(P2_N5798), .IN1(P2_N5797), .Q(P2_N411) );
  AND2X1 P2_C20210 ( .IN1(n6692), .IN2(P2_N117), .Q(P2_N5797) );
  AND2X1 P2_C20211 ( .IN1(n7479), .IN2(n6615), .Q(P2_N5798) );
  OR2X1 P2_C20213 ( .IN2(P2_N5800), .IN1(P2_N5799), .Q(P2_N412) );
  AND2X1 P2_C20214 ( .IN1(n6694), .IN2(P2_N116), .Q(P2_N5799) );
  AND2X1 P2_C20215 ( .IN1(n6693), .IN2(n6616), .Q(P2_N5800) );
  OR2X1 P2_C20217 ( .IN2(P2_N5802), .IN1(P2_N5801), .Q(P2_N413) );
  AND2X1 P2_C20218 ( .IN1(n6694), .IN2(P2_N115), .Q(P2_N5801) );
  AND2X1 P2_C20219 ( .IN1(n6693), .IN2(n6617), .Q(P2_N5802) );
  OR2X1 P2_C20221 ( .IN2(P2_N5804), .IN1(P2_N5803), .Q(P2_N414) );
  AND2X1 P2_C19948 ( .IN1(n6687), .IN2(n6719), .Q(P2_N5678) );
  OR2X1 P2_C19950 ( .IN2(P2_N5680), .IN1(P2_N5679), .Q(P2_N297) );
  AND2X1 P2_C19951 ( .IN1(n6690), .IN2(P2_N124), .Q(P2_N5679) );
  AND2X1 P2_C19952 ( .IN1(n19025), .IN2(n6608), .Q(P2_N5680) );
  OR2X1 P2_C19954 ( .IN2(P2_N5682), .IN1(P2_N5681), .Q(P2_N298) );
  AND2X1 P2_C19955 ( .IN1(n6690), .IN2(P2_N123), .Q(P2_N5681) );
  AND2X1 P2_C19956 ( .IN1(n19025), .IN2(n6609), .Q(P2_N5682) );
  OR2X1 P2_C19958 ( .IN2(P2_N5684), .IN1(P2_N5683), .Q(P2_N299) );
  AND2X1 P2_C19959 ( .IN1(n6696), .IN2(P2_N122), .Q(P2_N5683) );
  AND2X1 P2_C19960 ( .IN1(n6687), .IN2(n6610), .Q(P2_N5684) );
  OR2X1 P2_C19962 ( .IN2(P2_N5686), .IN1(P2_N5685), .Q(P2_N300) );
  AND2X1 P2_C19963 ( .IN1(n6696), .IN2(P2_N121), .Q(P2_N5685) );
  AND2X1 P2_C19964 ( .IN1(n6687), .IN2(n6611), .Q(P2_N5686) );
  OR2X1 P2_C19966 ( .IN2(P2_N5688), .IN1(P2_N5687), .Q(P2_N301) );
  AND2X1 P2_C19967 ( .IN1(n6696), .IN2(P2_N120), .Q(P2_N5687) );
  AND2X1 P2_C19968 ( .IN1(n6687), .IN2(n6612), .Q(P2_N5688) );
  OR2X1 P2_C19970 ( .IN2(P2_N5690), .IN1(P2_N5689), .Q(P2_N302) );
  AND2X1 P2_C19971 ( .IN1(n6692), .IN2(P2_N119), .Q(P2_N5689) );
  AND2X1 P2_C19972 ( .IN1(n7479), .IN2(n6613), .Q(P2_N5690) );
  OR2X1 P2_C19974 ( .IN2(P2_N5692), .IN1(P2_N5691), .Q(P2_N303) );
  AND2X1 P2_C19975 ( .IN1(n6692), .IN2(P2_N118), .Q(P2_N5691) );
  AND2X1 P2_C19976 ( .IN1(n7479), .IN2(n6614), .Q(P2_N5692) );
  OR2X1 P2_C19978 ( .IN2(P2_N5694), .IN1(P2_N5693), .Q(P2_N304) );
  AND2X1 P2_C19979 ( .IN1(n6692), .IN2(P2_N117), .Q(P2_N5693) );
  AND2X1 P2_C19980 ( .IN1(n7479), .IN2(n6615), .Q(P2_N5694) );
  OR2X1 P2_C19982 ( .IN2(P2_N5696), .IN1(P2_N5695), .Q(P2_N305) );
  AND2X1 P2_C19983 ( .IN1(n6694), .IN2(P2_N116), .Q(P2_N5695) );
  AND2X1 P2_C19984 ( .IN1(n6693), .IN2(n6616), .Q(P2_N5696) );
  OR2X1 P2_C19986 ( .IN2(P2_N5698), .IN1(P2_N5697), .Q(P2_N306) );
  AND2X1 P2_C19987 ( .IN1(n6694), .IN2(P2_N115), .Q(P2_N5697) );
  AND2X1 P2_C19988 ( .IN1(n6693), .IN2(n6617), .Q(P2_N5698) );
  OR2X1 P2_C19990 ( .IN2(P2_N5700), .IN1(P2_N5699), .Q(P2_N307) );
  AND2X1 P2_C19991 ( .IN1(n6694), .IN2(P2_N114), .Q(P2_N5699) );
  AND2X1 P2_C19992 ( .IN1(n6693), .IN2(n6607), .Q(P2_N5700) );
  OR2X1 P2_C19994 ( .IN2(P2_N5702), .IN1(P2_N5701), .Q(P2_N308) );
  AND2X1 P2_C19995 ( .IN1(n6698), .IN2(P2_N113), .Q(P2_N5701) );
  AND2X1 P2_C19996 ( .IN1(n7479), .IN2(n6606), .Q(P2_N5702) );
  OR2X1 P2_C19998 ( .IN2(P2_N5704), .IN1(P2_N5703), .Q(P2_N309) );
  AND2X1 P2_C19999 ( .IN1(n6698), .IN2(P2_N112), .Q(P2_N5703) );
  AND2X1 P2_C20000 ( .IN1(n7479), .IN2(n6605), .Q(P2_N5704) );
  OR2X1 P2_C20002 ( .IN2(P2_N5706), .IN1(P2_N5705), .Q(P2_N310) );
  AND2X1 P2_C20003 ( .IN1(n6698), .IN2(P2_N111), .Q(P2_N5705) );
  AND2X1 P2_C20004 ( .IN1(n7479), .IN2(n6604), .Q(P2_N5706) );
  OR2X1 P2_C20006 ( .IN2(P2_N5708), .IN1(P2_N5707), .Q(P2_N311) );
  AND2X1 P2_C20007 ( .IN1(n6686), .IN2(P2_N110), .Q(P2_N5707) );
  AND2X1 P2_C20008 ( .IN1(n6685), .IN2(n6603), .Q(P2_N5708) );
  OR2X1 P2_C20010 ( .IN2(P2_N5710), .IN1(P2_N5709), .Q(P2_N312) );
  AND2X1 P2_C20011 ( .IN1(n6686), .IN2(P2_N109), .Q(P2_N5709) );
  AND2X1 P2_C20012 ( .IN1(n6685), .IN2(n6602), .Q(P2_N5710) );
  OR2X1 P2_C20014 ( .IN2(P2_N5712), .IN1(P2_N5711), .Q(P2_N313) );
  AND2X1 P2_C20015 ( .IN1(n6686), .IN2(P2_N108), .Q(P2_N5711) );
  AND2X1 P2_C20016 ( .IN1(n6685), .IN2(n6601), .Q(P2_N5712) );
  OR2X1 P2_C20018 ( .IN2(P2_N5714), .IN1(P2_N5713), .Q(P2_N314) );
  AND2X1 P2_C20019 ( .IN1(n6700), .IN2(P2_N107), .Q(P2_N5713) );
  AND2X1 P2_C20020 ( .IN1(n6699), .IN2(n6600), .Q(P2_N5714) );
  OR2X1 P2_C20022 ( .IN2(P2_N5716), .IN1(P2_N5715), .Q(P2_N315) );
  AND2X1 P2_C20023 ( .IN1(n6700), .IN2(P2_N106), .Q(P2_N5715) );
  AND2X1 P2_C20024 ( .IN1(n6699), .IN2(n6599), .Q(P2_N5716) );
  OR2X1 P2_C20026 ( .IN2(P2_N5718), .IN1(P2_N5717), .Q(P2_N316) );
  AND2X1 P2_C20027 ( .IN1(n6700), .IN2(P2_N105), .Q(P2_N5717) );
  AND2X1 P2_C20028 ( .IN1(n6699), .IN2(n6598), .Q(P2_N5718) );
  OR2X1 P2_C20030 ( .IN2(P2_N5720), .IN1(P2_N5719), .Q(P2_N317) );
  AND2X1 P2_C20031 ( .IN1(n6702), .IN2(P2_N104), .Q(P2_N5719) );
  AND2X1 P2_C20032 ( .IN1(n19025), .IN2(n6597), .Q(P2_N5720) );
  OR2X1 P2_C20034 ( .IN2(P2_N5722), .IN1(P2_N5721), .Q(P2_N318) );
  AND2X1 P2_C20035 ( .IN1(n6702), .IN2(P2_N103), .Q(P2_N5721) );
  AND2X1 P2_C20036 ( .IN1(n19025), .IN2(n6596), .Q(P2_N5722) );
  OR2X1 P2_C20038 ( .IN2(P2_N5724), .IN1(P2_N5723), .Q(P2_N319) );
  AND2X1 P2_C20039 ( .IN1(n6696), .IN2(n6595), .Q(P2_N5723) );
  AND2X1 P2_C20040 ( .IN1(n19025), .IN2(n6595), .Q(P2_N5724) );
  OR2X1 P2_C20065 ( .IN2(P2_N5726), .IN1(P2_N5725), .Q(P2_N344) );
  AND2X1 P2_C20066 ( .IN1(n6690), .IN2(P2_N121), .Q(P2_N5725) );
  AND2X1 P2_C20067 ( .IN1(n19025), .IN2(n6611), .Q(P2_N5726) );
  OR2X1 P2_C20069 ( .IN2(P2_N5728), .IN1(P2_N5727), .Q(P2_N345) );
  AND2X1 P2_C20070 ( .IN1(n6696), .IN2(P2_N120), .Q(P2_N5727) );
  AND2X1 P2_C20071 ( .IN1(n6687), .IN2(n6612), .Q(P2_N5728) );
  OR2X1 P2_C20073 ( .IN2(P2_N5730), .IN1(P2_N5729), .Q(P2_N346) );
  AND2X1 P2_C20074 ( .IN1(n6696), .IN2(P2_N119), .Q(P2_N5729) );
  AND2X1 P2_C20075 ( .IN1(n6687), .IN2(n6613), .Q(P2_N5730) );
  OR2X1 P2_C20077 ( .IN2(P2_N5732), .IN1(P2_N5731), .Q(P2_N347) );
  AND2X1 P2_C20078 ( .IN1(n6692), .IN2(P2_N118), .Q(P2_N5731) );
  AND2X1 P2_C20079 ( .IN1(n7479), .IN2(n6614), .Q(P2_N5732) );
  OR2X1 P2_C20081 ( .IN2(P2_N5734), .IN1(P2_N5733), .Q(P2_N348) );
  AND2X1 P2_C20082 ( .IN1(n6692), .IN2(P2_N117), .Q(P2_N5733) );
  AND2X1 P2_C20083 ( .IN1(n7479), .IN2(n6615), .Q(P2_N5734) );
  OR2X1 P2_C20085 ( .IN2(P2_N5736), .IN1(P2_N5735), .Q(P2_N349) );
  AND2X1 P2_C20086 ( .IN1(n6694), .IN2(P2_N116), .Q(P2_N5735) );
  AND2X1 P2_C20087 ( .IN1(n6693), .IN2(n6616), .Q(P2_N5736) );
  OR2X1 P2_C20089 ( .IN2(P2_N5738), .IN1(P2_N5737), .Q(P2_N350) );
  AND2X1 P2_C20090 ( .IN1(n6694), .IN2(P2_N115), .Q(P2_N5737) );
  AND2X1 P2_C20091 ( .IN1(n6693), .IN2(n6617), .Q(P2_N5738) );
  OR2X1 P2_C20093 ( .IN2(P2_N5740), .IN1(P2_N5739), .Q(P2_N351) );
  AND2X1 P2_C20094 ( .IN1(n6694), .IN2(P2_N114), .Q(P2_N5739) );
  AND2X1 P2_C19776 ( .IN1(n6686), .IN2(P2_N108), .Q(P2_N5613) );
  AND2X1 P2_C19777 ( .IN1(n6685), .IN2(n6601), .Q(P2_N5614) );
  OR2X1 P2_C19779 ( .IN2(P2_N5616), .IN1(P2_N5615), .Q(P2_N215) );
  AND2X1 P2_C19780 ( .IN1(n6700), .IN2(P2_N107), .Q(P2_N5615) );
  AND2X1 P2_C19781 ( .IN1(n6699), .IN2(n6600), .Q(P2_N5616) );
  OR2X1 P2_C19783 ( .IN2(P2_N5618), .IN1(P2_N5617), .Q(P2_N216) );
  AND2X1 P2_C19784 ( .IN1(n6700), .IN2(P2_N106), .Q(P2_N5617) );
  AND2X1 P2_C19785 ( .IN1(n6699), .IN2(n6599), .Q(P2_N5618) );
  OR2X1 P2_C19787 ( .IN2(P2_N5620), .IN1(P2_N5619), .Q(P2_N217) );
  AND2X1 P2_C19788 ( .IN1(n6700), .IN2(P2_N105), .Q(P2_N5619) );
  AND2X1 P2_C19789 ( .IN1(n6699), .IN2(n6598), .Q(P2_N5620) );
  OR2X1 P2_C19791 ( .IN2(P2_N5622), .IN1(P2_N5621), .Q(P2_N218) );
  AND2X1 P2_C19792 ( .IN1(n6702), .IN2(P2_N104), .Q(P2_N5621) );
  AND2X1 P2_C19793 ( .IN1(n19025), .IN2(n6597), .Q(P2_N5622) );
  OR2X1 P2_C19795 ( .IN2(P2_N5624), .IN1(P2_N5623), .Q(P2_N219) );
  AND2X1 P2_C19796 ( .IN1(n6702), .IN2(P2_N103), .Q(P2_N5623) );
  AND2X1 P2_C19797 ( .IN1(n19025), .IN2(n6596), .Q(P2_N5624) );
  OR2X1 P2_C19799 ( .IN2(P2_N5626), .IN1(P2_N5625), .Q(P2_N220) );
  AND2X1 P2_C19800 ( .IN1(n6702), .IN2(n6595), .Q(P2_N5625) );
  AND2X1 P2_C19801 ( .IN1(n19025), .IN2(n6595), .Q(P2_N5626) );
  AND2X1 P2_C19828 ( .IN1(n6690), .IN2(P2_N133), .Q(P2_N248) );
  OR2X1 P2_C19831 ( .IN2(P2_N5630), .IN1(P2_N5629), .Q(P2_N249) );
  AND2X1 P2_C19832 ( .IN1(n6690), .IN2(P2_N124), .Q(P2_N5629) );
  AND2X1 P2_C19833 ( .IN1(n19025), .IN2(n6608), .Q(P2_N5630) );
  AND2X1 P2_C19836 ( .IN1(n6690), .IN2(P2_N123), .Q(P2_N5631) );
  AND2X1 P2_C19837 ( .IN1(n19025), .IN2(n6609), .Q(P2_N5632) );
  OR2X1 P2_C19839 ( .IN2(P2_N5634), .IN1(P2_N5633), .Q(P2_N251) );
  AND2X1 P2_C19840 ( .IN1(n6690), .IN2(P2_N122), .Q(P2_N5633) );
  AND2X1 P2_C19841 ( .IN1(n19025), .IN2(n6610), .Q(P2_N5634) );
  OR2X1 P2_C19843 ( .IN2(P2_N5636), .IN1(P2_N5635), .Q(P2_N252) );
  AND2X1 P2_C19844 ( .IN1(n6690), .IN2(P2_N121), .Q(P2_N5635) );
  AND2X1 P2_C19845 ( .IN1(n19025), .IN2(n6611), .Q(P2_N5636) );
  OR2X1 P2_C19847 ( .IN2(P2_N5638), .IN1(P2_N5637), .Q(P2_N253) );
  AND2X1 P2_C19848 ( .IN1(n6696), .IN2(P2_N120), .Q(P2_N5637) );
  AND2X1 P2_C19849 ( .IN1(n6687), .IN2(n6612), .Q(P2_N5638) );
  OR2X1 P2_C19851 ( .IN2(P2_N5640), .IN1(P2_N5639), .Q(P2_N254) );
  AND2X1 P2_C19852 ( .IN1(n6692), .IN2(P2_N119), .Q(P2_N5639) );
  AND2X1 P2_C19853 ( .IN1(n7479), .IN2(n6613), .Q(P2_N5640) );
  OR2X1 P2_C19855 ( .IN2(P2_N5642), .IN1(P2_N5641), .Q(P2_N255) );
  AND2X1 P2_C19856 ( .IN1(n6692), .IN2(P2_N118), .Q(P2_N5641) );
  AND2X1 P2_C19857 ( .IN1(n7479), .IN2(n6614), .Q(P2_N5642) );
  OR2X1 P2_C19859 ( .IN2(P2_N5644), .IN1(P2_N5643), .Q(P2_N256) );
  AND2X1 P2_C19860 ( .IN1(n6694), .IN2(P2_N117), .Q(P2_N5643) );
  AND2X1 P2_C19861 ( .IN1(n7479), .IN2(n6615), .Q(P2_N5644) );
  OR2X1 P2_C19863 ( .IN2(P2_N5646), .IN1(P2_N5645), .Q(P2_N257) );
  AND2X1 P2_C19864 ( .IN1(n6694), .IN2(P2_N116), .Q(P2_N5645) );
  AND2X1 P2_C19865 ( .IN1(n6693), .IN2(n6616), .Q(P2_N5646) );
  OR2X1 P2_C19867 ( .IN2(P2_N5648), .IN1(P2_N5647), .Q(P2_N258) );
  AND2X1 P2_C19868 ( .IN1(n6694), .IN2(P2_N115), .Q(P2_N5647) );
  AND2X1 P2_C19869 ( .IN1(n6693), .IN2(n6617), .Q(P2_N5648) );
  OR2X1 P2_C19871 ( .IN2(P2_N5650), .IN1(P2_N5649), .Q(P2_N259) );
  AND2X1 P2_C19872 ( .IN1(n6694), .IN2(P2_N114), .Q(P2_N5649) );
  AND2X1 P2_C19873 ( .IN1(n6693), .IN2(n6607), .Q(P2_N5650) );
  OR2X1 P2_C19875 ( .IN2(P2_N5652), .IN1(P2_N5651), .Q(P2_N260) );
  AND2X1 P2_C19876 ( .IN1(n6698), .IN2(P2_N113), .Q(P2_N5651) );
  AND2X1 P2_C19877 ( .IN1(n7479), .IN2(n6606), .Q(P2_N5652) );
  OR2X1 P2_C19879 ( .IN2(P2_N5654), .IN1(P2_N5653), .Q(P2_N261) );
  AND2X1 P2_C19880 ( .IN1(n6698), .IN2(P2_N112), .Q(P2_N5653) );
  AND2X1 P2_C19881 ( .IN1(n7479), .IN2(n6605), .Q(P2_N5654) );
  OR2X1 P2_C19883 ( .IN2(P2_N5656), .IN1(P2_N5655), .Q(P2_N262) );
  AND2X1 P2_C19884 ( .IN1(n6698), .IN2(P2_N111), .Q(P2_N5655) );
  AND2X1 P2_C19885 ( .IN1(n7479), .IN2(n6604), .Q(P2_N5656) );
  OR2X1 P2_C19887 ( .IN2(P2_N5658), .IN1(P2_N5657), .Q(P2_N263) );
  AND2X1 P2_C19888 ( .IN1(n6686), .IN2(P2_N110), .Q(P2_N5657) );
  AND2X1 P2_C19889 ( .IN1(n6685), .IN2(n6603), .Q(P2_N5658) );
  OR2X1 P2_C19891 ( .IN2(P2_N5660), .IN1(P2_N5659), .Q(P2_N264) );
  AND2X1 P2_C19892 ( .IN1(n6686), .IN2(P2_N109), .Q(P2_N5659) );
  AND2X1 P2_C19893 ( .IN1(n6685), .IN2(n6602), .Q(P2_N5660) );
  OR2X1 P2_C19895 ( .IN2(P2_N5662), .IN1(P2_N5661), .Q(P2_N265) );
  AND2X1 P2_C19896 ( .IN1(n6686), .IN2(P2_N108), .Q(P2_N5661) );
  AND2X1 P2_C19897 ( .IN1(n6685), .IN2(n6601), .Q(P2_N5662) );
  OR2X1 P2_C19899 ( .IN2(P2_N5664), .IN1(P2_N5663), .Q(P2_N266) );
  AND2X1 P2_C19900 ( .IN1(n6686), .IN2(P2_N107), .Q(P2_N5663) );
  AND2X1 P2_C19901 ( .IN1(n6685), .IN2(n6600), .Q(P2_N5664) );
  OR2X1 P2_C19903 ( .IN2(P2_N5666), .IN1(P2_N5665), .Q(P2_N267) );
  AND2X1 P2_C19904 ( .IN1(n6700), .IN2(P2_N106), .Q(P2_N5665) );
  AND2X1 P2_C19905 ( .IN1(n6699), .IN2(n6599), .Q(P2_N5666) );
  OR2X1 P2_C19907 ( .IN2(P2_N5668), .IN1(P2_N5667), .Q(P2_N268) );
  AND2X1 P2_C19908 ( .IN1(n6700), .IN2(P2_N105), .Q(P2_N5667) );
  AND2X1 P2_C19909 ( .IN1(n6699), .IN2(n6598), .Q(P2_N5668) );
  OR2X1 P2_C19911 ( .IN2(P2_N5670), .IN1(P2_N5669), .Q(P2_N269) );
  AND2X1 P2_C19912 ( .IN1(n6702), .IN2(P2_N104), .Q(P2_N5669) );
  AND2X1 P2_C19913 ( .IN1(n19025), .IN2(n6597), .Q(P2_N5670) );
  OR2X1 P2_C19915 ( .IN2(P2_N5672), .IN1(P2_N5671), .Q(P2_N270) );
  AND2X1 P2_C19916 ( .IN1(n6696), .IN2(P2_N103), .Q(P2_N5671) );
  AND2X1 P2_C19917 ( .IN1(n19025), .IN2(n6596), .Q(P2_N5672) );
  OR2X1 P2_C19919 ( .IN2(P2_N5674), .IN1(P2_N5673), .Q(P2_N271) );
  AND2X1 P2_C19920 ( .IN1(n6696), .IN2(n6595), .Q(P2_N5673) );
  AND2X1 P2_C19921 ( .IN1(n6687), .IN2(n6595), .Q(P2_N5674) );
  AND2X1 P2_C19943 ( .IN1(n6690), .IN2(P2_N133), .Q(P2_N295) );
  AND2X1 P2_C19947 ( .IN1(n6688), .IN2(P2_N125), .Q(P2_N5677) );
  AND2X1 P2_C19622 ( .IN1(n7479), .IN2(n6605), .Q(P2_N5550) );
  OR2X1 P2_C19624 ( .IN2(P2_N5552), .IN1(P2_N5551), .Q(P2_N154) );
  AND2X1 P2_C19625 ( .IN1(n6686), .IN2(P2_N111), .Q(P2_N5551) );
  AND2X1 P2_C19626 ( .IN1(n6685), .IN2(n6604), .Q(P2_N5552) );
  OR2X1 P2_C19628 ( .IN2(P2_N5554), .IN1(P2_N5553), .Q(P2_N155) );
  AND2X1 P2_C19629 ( .IN1(n6686), .IN2(P2_N110), .Q(P2_N5553) );
  AND2X1 P2_C19630 ( .IN1(n6685), .IN2(n6603), .Q(P2_N5554) );
  OR2X1 P2_C19632 ( .IN2(P2_N5556), .IN1(P2_N5555), .Q(P2_N156) );
  AND2X1 P2_C19633 ( .IN1(n6686), .IN2(P2_N109), .Q(P2_N5555) );
  AND2X1 P2_C19634 ( .IN1(n6685), .IN2(n6602), .Q(P2_N5556) );
  OR2X1 P2_C19636 ( .IN2(P2_N5558), .IN1(P2_N5557), .Q(P2_N157) );
  AND2X1 P2_C19637 ( .IN1(n6700), .IN2(P2_N108), .Q(P2_N5557) );
  AND2X1 P2_C19638 ( .IN1(n6699), .IN2(n6601), .Q(P2_N5558) );
  OR2X1 P2_C19640 ( .IN2(P2_N5560), .IN1(P2_N5559), .Q(P2_N158) );
  AND2X1 P2_C19641 ( .IN1(n6700), .IN2(P2_N107), .Q(P2_N5559) );
  AND2X1 P2_C19642 ( .IN1(n6699), .IN2(n6600), .Q(P2_N5560) );
  OR2X1 P2_C19644 ( .IN2(P2_N5562), .IN1(P2_N5561), .Q(P2_N159) );
  AND2X1 P2_C19645 ( .IN1(n6700), .IN2(P2_N106), .Q(P2_N5561) );
  AND2X1 P2_C19646 ( .IN1(n6699), .IN2(n6599), .Q(P2_N5562) );
  OR2X1 P2_C19648 ( .IN2(P2_N5564), .IN1(P2_N5563), .Q(P2_N160) );
  AND2X1 P2_C19649 ( .IN1(n6702), .IN2(P2_N105), .Q(P2_N5563) );
  AND2X1 P2_C19650 ( .IN1(n19025), .IN2(n6598), .Q(P2_N5564) );
  OR2X1 P2_C19652 ( .IN2(P2_N5566), .IN1(P2_N5565), .Q(P2_N161) );
  AND2X1 P2_C19653 ( .IN1(n6702), .IN2(P2_N104), .Q(P2_N5565) );
  AND2X1 P2_C19654 ( .IN1(n19025), .IN2(n6597), .Q(P2_N5566) );
  OR2X1 P2_C19656 ( .IN2(P2_N5568), .IN1(P2_N5567), .Q(P2_N162) );
  AND2X1 P2_C19657 ( .IN1(n6702), .IN2(P2_N103), .Q(P2_N5567) );
  AND2X1 P2_C19658 ( .IN1(n19025), .IN2(n6596), .Q(P2_N5568) );
  OR2X1 P2_C19660 ( .IN2(P2_N5570), .IN1(P2_N5569), .Q(P2_N163) );
  AND2X1 P2_C19661 ( .IN1(n6692), .IN2(n6595), .Q(P2_N5569) );
  AND2X1 P2_C19662 ( .IN1(n19025), .IN2(n6595), .Q(P2_N5570) );
  AND2X1 P2_C19692 ( .IN1(n6688), .IN2(P2_N133), .Q(P2_N193) );
  OR2X1 P2_C19695 ( .IN2(P2_N5574), .IN1(P2_N5573), .Q(P2_N194) );
  AND2X1 P2_C19696 ( .IN1(n6688), .IN2(P2_N128), .Q(P2_N5573) );
  AND2X1 P2_C19697 ( .IN1(n6687), .IN2(n10183), .Q(P2_N5574) );
  AND2X1 P2_C19700 ( .IN1(n6688), .IN2(P2_N127), .Q(P2_N5575) );
  AND2X1 P2_C19701 ( .IN1(n6687), .IN2(n10377), .Q(P2_N5576) );
  OR2X1 P2_C19703 ( .IN2(P2_N5578), .IN1(P2_N5577), .Q(P2_N196) );
  AND2X1 P2_C19704 ( .IN1(n6688), .IN2(P2_N126), .Q(P2_N5577) );
  AND2X1 P2_C19705 ( .IN1(n6687), .IN2(n10191), .Q(P2_N5578) );
  OR2X1 P2_C19707 ( .IN2(P2_N5580), .IN1(P2_N5579), .Q(P2_N197) );
  AND2X1 P2_C19708 ( .IN1(n6688), .IN2(P2_N125), .Q(P2_N5579) );
  AND2X1 P2_C19709 ( .IN1(n6687), .IN2(n6719), .Q(P2_N5580) );
  OR2X1 P2_C19711 ( .IN2(P2_N5582), .IN1(P2_N5581), .Q(P2_N198) );
  AND2X1 P2_C19712 ( .IN1(n6690), .IN2(P2_N124), .Q(P2_N5581) );
  AND2X1 P2_C19713 ( .IN1(n19025), .IN2(n6608), .Q(P2_N5582) );
  OR2X1 P2_C19715 ( .IN2(P2_N5584), .IN1(P2_N5583), .Q(P2_N199) );
  AND2X1 P2_C19716 ( .IN1(n6690), .IN2(P2_N123), .Q(P2_N5583) );
  AND2X1 P2_C19717 ( .IN1(n19025), .IN2(n6609), .Q(P2_N5584) );
  OR2X1 P2_C19719 ( .IN2(P2_N5586), .IN1(P2_N5585), .Q(P2_N200) );
  AND2X1 P2_C19720 ( .IN1(n6696), .IN2(P2_N122), .Q(P2_N5585) );
  AND2X1 P2_C19721 ( .IN1(n6687), .IN2(n6610), .Q(P2_N5586) );
  OR2X1 P2_C19723 ( .IN2(P2_N5588), .IN1(P2_N5587), .Q(P2_N201) );
  AND2X1 P2_C19724 ( .IN1(n6696), .IN2(P2_N121), .Q(P2_N5587) );
  AND2X1 P2_C19725 ( .IN1(n6687), .IN2(n6611), .Q(P2_N5588) );
  OR2X1 P2_C19727 ( .IN2(P2_N5590), .IN1(P2_N5589), .Q(P2_N202) );
  AND2X1 P2_C19728 ( .IN1(n6696), .IN2(P2_N120), .Q(P2_N5589) );
  AND2X1 P2_C19729 ( .IN1(n6687), .IN2(n6612), .Q(P2_N5590) );
  OR2X1 P2_C19731 ( .IN2(P2_N5592), .IN1(P2_N5591), .Q(P2_N203) );
  AND2X1 P2_C19732 ( .IN1(n6692), .IN2(P2_N119), .Q(P2_N5591) );
  AND2X1 P2_C19733 ( .IN1(n7479), .IN2(n6613), .Q(P2_N5592) );
  OR2X1 P2_C19735 ( .IN2(P2_N5594), .IN1(P2_N5593), .Q(P2_N204) );
  AND2X1 P2_C19736 ( .IN1(n6692), .IN2(P2_N118), .Q(P2_N5593) );
  AND2X1 P2_C19737 ( .IN1(n7479), .IN2(n6614), .Q(P2_N5594) );
  OR2X1 P2_C19739 ( .IN2(P2_N5596), .IN1(P2_N5595), .Q(P2_N205) );
  AND2X1 P2_C19740 ( .IN1(n6692), .IN2(P2_N117), .Q(P2_N5595) );
  AND2X1 P2_C19741 ( .IN1(n7479), .IN2(n6615), .Q(P2_N5596) );
  OR2X1 P2_C19743 ( .IN2(P2_N5598), .IN1(P2_N5597), .Q(P2_N206) );
  AND2X1 P2_C19744 ( .IN1(n6694), .IN2(P2_N116), .Q(P2_N5597) );
  AND2X1 P2_C19745 ( .IN1(n6693), .IN2(n6616), .Q(P2_N5598) );
  OR2X1 P2_C19747 ( .IN2(P2_N5600), .IN1(P2_N5599), .Q(P2_N207) );
  AND2X1 P2_C19748 ( .IN1(n6694), .IN2(P2_N115), .Q(P2_N5599) );
  AND2X1 P2_C19749 ( .IN1(n6693), .IN2(n6617), .Q(P2_N5600) );
  OR2X1 P2_C19751 ( .IN2(P2_N5602), .IN1(P2_N5601), .Q(P2_N208) );
  AND2X1 P2_C19752 ( .IN1(n6694), .IN2(P2_N114), .Q(P2_N5601) );
  AND2X1 P2_C19753 ( .IN1(n6693), .IN2(n6607), .Q(P2_N5602) );
  OR2X1 P2_C19755 ( .IN2(P2_N5604), .IN1(P2_N5603), .Q(P2_N209) );
  AND2X1 P2_C19756 ( .IN1(n6698), .IN2(P2_N113), .Q(P2_N5603) );
  AND2X1 P2_C19757 ( .IN1(n7479), .IN2(n6606), .Q(P2_N5604) );
  OR2X1 P2_C19759 ( .IN2(P2_N5606), .IN1(P2_N5605), .Q(P2_N210) );
  AND2X1 P2_C19760 ( .IN1(n6698), .IN2(P2_N112), .Q(P2_N5605) );
  AND2X1 P2_C19761 ( .IN1(n7479), .IN2(n6605), .Q(P2_N5606) );
  OR2X1 P2_C19763 ( .IN2(P2_N5608), .IN1(P2_N5607), .Q(P2_N211) );
  AND2X1 P2_C19764 ( .IN1(n6698), .IN2(P2_N111), .Q(P2_N5607) );
  AND2X1 P2_C19765 ( .IN1(n7479), .IN2(n6604), .Q(P2_N5608) );
  OR2X1 P2_C19767 ( .IN2(P2_N5610), .IN1(P2_N5609), .Q(P2_N212) );
  AND2X1 P2_C19768 ( .IN1(n6686), .IN2(P2_N110), .Q(P2_N5609) );
  AND2X1 P2_C19769 ( .IN1(n6685), .IN2(n6603), .Q(P2_N5610) );
  OR2X1 P2_C19771 ( .IN2(P2_N5612), .IN1(P2_N5611), .Q(P2_N213) );
  AND2X1 P2_C19772 ( .IN1(n6686), .IN2(P2_N109), .Q(P2_N5611) );
  AND2X1 P2_C19773 ( .IN1(n6685), .IN2(n6602), .Q(P2_N5612) );
  OR2X1 P2_C19775 ( .IN2(P2_N5614), .IN1(P2_N5613), .Q(P2_N214) );
  AND2X1 P2_C1092 ( .IN1(n6972), .IN2(n6940), .Q(P2_N541) );
  AND2X1 P2_C1093 ( .IN1(n6838), .IN2(n6784), .Q(P2_N542) );
  OR2X1 P2_C16127 ( .IN2(n7341), .IN1(n7334), .Q(P2_N5492) );
  OR2X1 P2_C16167 ( .IN2(n7334), .IN1(n6999), .Q(P2_N5493) );
  AND2X1 P2_C19545 ( .IN1(n6688), .IN2(P2_N133), .Q(P2_N134) );
  OR2X1 P2_C19548 ( .IN2(P2_N5514), .IN1(P2_N5513), .Q(P2_N135) );
  AND2X1 P2_C19549 ( .IN1(n6688), .IN2(P2_N130), .Q(P2_N5513) );
  AND2X1 P2_C19550 ( .IN1(n6687), .IN2(n10141), .Q(P2_N5514) );
  OR2X1 P2_C19552 ( .IN2(P2_N5516), .IN1(P2_N5515), .Q(P2_N136) );
  AND2X1 P2_C19553 ( .IN1(n6688), .IN2(P2_N129), .Q(P2_N5515) );
  AND2X1 P2_C19554 ( .IN1(n6687), .IN2(n10369), .Q(P2_N5516) );
  OR2X1 P2_C19556 ( .IN2(P2_N5518), .IN1(P2_N5517), .Q(P2_N137) );
  AND2X1 P2_C19557 ( .IN1(n6688), .IN2(P2_N128), .Q(P2_N5517) );
  AND2X1 P2_C19558 ( .IN1(n6687), .IN2(n10183), .Q(P2_N5518) );
  OR2X1 P2_C19560 ( .IN2(P2_N5520), .IN1(P2_N5519), .Q(P2_N138) );
  AND2X1 P2_C19561 ( .IN1(n6688), .IN2(P2_N127), .Q(P2_N5519) );
  AND2X1 P2_C19562 ( .IN1(n6687), .IN2(n10377), .Q(P2_N5520) );
  OR2X1 P2_C19564 ( .IN2(P2_N5522), .IN1(P2_N5521), .Q(P2_N139) );
  AND2X1 P2_C19565 ( .IN1(n6688), .IN2(P2_N126), .Q(P2_N5521) );
  AND2X1 P2_C19566 ( .IN1(n6687), .IN2(n10191), .Q(P2_N5522) );
  OR2X1 P2_C19568 ( .IN2(P2_N5524), .IN1(P2_N5523), .Q(P2_N140) );
  AND2X1 P2_C19569 ( .IN1(n6688), .IN2(P2_N125), .Q(P2_N5523) );
  AND2X1 P2_C19570 ( .IN1(n6687), .IN2(n6719), .Q(P2_N5524) );
  OR2X1 P2_C19572 ( .IN2(P2_N5526), .IN1(P2_N5525), .Q(P2_N141) );
  AND2X1 P2_C19573 ( .IN1(n6690), .IN2(P2_N124), .Q(P2_N5525) );
  AND2X1 P2_C19574 ( .IN1(n19025), .IN2(n6608), .Q(P2_N5526) );
  OR2X1 P2_C19576 ( .IN2(P2_N5528), .IN1(P2_N5527), .Q(P2_N142) );
  AND2X1 P2_C19577 ( .IN1(n6690), .IN2(P2_N123), .Q(P2_N5527) );
  AND2X1 P2_C19578 ( .IN1(n19025), .IN2(n6609), .Q(P2_N5528) );
  OR2X1 P2_C19580 ( .IN2(P2_N5530), .IN1(P2_N5529), .Q(P2_N143) );
  AND2X1 P2_C19581 ( .IN1(n6696), .IN2(P2_N122), .Q(P2_N5529) );
  AND2X1 P2_C19582 ( .IN1(n6687), .IN2(n6610), .Q(P2_N5530) );
  OR2X1 P2_C19584 ( .IN2(P2_N5532), .IN1(P2_N5531), .Q(P2_N144) );
  AND2X1 P2_C19585 ( .IN1(n6696), .IN2(P2_N121), .Q(P2_N5531) );
  AND2X1 P2_C19586 ( .IN1(n6687), .IN2(n6611), .Q(P2_N5532) );
  OR2X1 P2_C19588 ( .IN2(P2_N5534), .IN1(P2_N5533), .Q(P2_N145) );
  AND2X1 P2_C19589 ( .IN1(n6696), .IN2(P2_N120), .Q(P2_N5533) );
  AND2X1 P2_C19590 ( .IN1(n6687), .IN2(n6612), .Q(P2_N5534) );
  OR2X1 P2_C19592 ( .IN2(P2_N5536), .IN1(P2_N5535), .Q(P2_N146) );
  AND2X1 P2_C19593 ( .IN1(n6692), .IN2(P2_N119), .Q(P2_N5535) );
  AND2X1 P2_C19594 ( .IN1(n7479), .IN2(n6613), .Q(P2_N5536) );
  OR2X1 P2_C19596 ( .IN2(P2_N5538), .IN1(P2_N5537), .Q(P2_N147) );
  AND2X1 P2_C19597 ( .IN1(n6692), .IN2(P2_N118), .Q(P2_N5537) );
  AND2X1 P2_C19598 ( .IN1(n7479), .IN2(n6614), .Q(P2_N5538) );
  OR2X1 P2_C19600 ( .IN2(P2_N5540), .IN1(P2_N5539), .Q(P2_N148) );
  AND2X1 P2_C19601 ( .IN1(n6692), .IN2(P2_N117), .Q(P2_N5539) );
  AND2X1 P2_C19602 ( .IN1(n7479), .IN2(n6615), .Q(P2_N5540) );
  OR2X1 P2_C19604 ( .IN2(P2_N5542), .IN1(P2_N5541), .Q(P2_N149) );
  AND2X1 P2_C19605 ( .IN1(n6694), .IN2(P2_N116), .Q(P2_N5541) );
  AND2X1 P2_C19606 ( .IN1(n6693), .IN2(n6616), .Q(P2_N5542) );
  OR2X1 P2_C19608 ( .IN2(P2_N5544), .IN1(P2_N5543), .Q(P2_N150) );
  AND2X1 P2_C19609 ( .IN1(n6694), .IN2(P2_N115), .Q(P2_N5543) );
  AND2X1 P2_C19610 ( .IN1(n6693), .IN2(n6617), .Q(P2_N5544) );
  OR2X1 P2_C19612 ( .IN2(P2_N5546), .IN1(P2_N5545), .Q(P2_N151) );
  AND2X1 P2_C19613 ( .IN1(n6694), .IN2(P2_N114), .Q(P2_N5545) );
  AND2X1 P2_C19614 ( .IN1(n6693), .IN2(n6607), .Q(P2_N5546) );
  OR2X1 P2_C19616 ( .IN2(P2_N5548), .IN1(P2_N5547), .Q(P2_N152) );
  AND2X1 P2_C19617 ( .IN1(n6698), .IN2(P2_N113), .Q(P2_N5547) );
  AND2X1 P2_C19618 ( .IN1(n7479), .IN2(n6606), .Q(P2_N5548) );
  OR2X1 P2_C19620 ( .IN2(P2_N5550), .IN1(P2_N5549), .Q(P2_N153) );
  AND2X1 P2_C19621 ( .IN1(n6698), .IN2(P2_N112), .Q(P2_N5549) );
  NAND2X0 P2_lt_696_U21 ( .IN1(P2_N5032), .IN2(P2_lt_696_n28), 
        .QN(P2_lt_696_n27) );
  NAND2X0 P2_lt_696_U20 ( .IN1(P2_lt_696_n26), .IN2(P2_lt_696_n27), 
        .QN(P2_lt_696_n25) );
  NOR2X0 P2_lt_696_U19 ( .QN(P2_lt_696_n21), .IN1(P2_lt_696_n24), 
        .IN2(P2_lt_696_n25) );
  NOR2X0 P2_lt_696_U18 ( .QN(P2_lt_696_n22), .IN1(P2_N5033), 
        .IN2(P2_lt_696_n23) );
  NOR2X0 P2_lt_696_U17 ( .QN(P2_lt_696_n19), .IN1(P2_lt_696_n21), 
        .IN2(P2_lt_696_n22) );
  INVX0 P2_lt_696_U16 ( .ZN(P2_lt_696_n18), .INP(P2_N5349) );
  OR2X1 P2_lt_696_U15 ( .IN2(P2_N5034), .IN1(P2_lt_696_n18), .Q(P2_lt_696_n20)
         );
  NAND2X0 P2_lt_696_U14 ( .IN1(P2_lt_696_n19), .IN2(P2_lt_696_n20), 
        .QN(P2_lt_696_n16) );
  NAND2X0 P2_lt_696_U13 ( .IN1(P2_N5034), .IN2(P2_lt_696_n18), 
        .QN(P2_lt_696_n17) );
  NAND2X0 P2_lt_696_U12 ( .IN1(P2_lt_696_n16), .IN2(P2_lt_696_n17), 
        .QN(P2_lt_696_n15) );
  NOR2X0 P2_lt_696_U11 ( .QN(P2_lt_696_n11), .IN1(P2_lt_696_n14), 
        .IN2(P2_lt_696_n15) );
  NOR2X0 P2_lt_696_U10 ( .QN(P2_lt_696_n12), .IN1(P2_N5035), 
        .IN2(P2_lt_696_n13) );
  NOR2X0 P2_lt_696_U9 ( .QN(P2_lt_696_n9), .IN1(P2_lt_696_n11), 
        .IN2(P2_lt_696_n12) );
  INVX0 P2_lt_696_U8 ( .ZN(P2_lt_696_n8), .INP(P2_N5351) );
  OR2X1 P2_lt_696_U7 ( .IN2(P2_N5036), .IN1(P2_lt_696_n8), .Q(P2_lt_696_n10)
         );
  NAND2X0 P2_lt_696_U6 ( .IN1(P2_lt_696_n9), .IN2(P2_lt_696_n10), 
        .QN(P2_lt_696_n6) );
  NAND2X0 P2_lt_696_U5 ( .IN1(P2_N5036), .IN2(P2_lt_696_n8), .QN(P2_lt_696_n7)
         );
  NAND2X0 P2_lt_696_U4 ( .IN1(P2_lt_696_n6), .IN2(P2_lt_696_n7), 
        .QN(P2_lt_696_n3) );
  NAND2X0 P2_lt_696_U3 ( .IN1(P2_N5037), .IN2(P2_lt_696_n5), .QN(P2_lt_696_n4)
         );
  NAND2X0 P2_lt_696_U2 ( .IN1(P2_lt_696_n3), .IN2(P2_lt_696_n4), 
        .QN(P2_lt_696_n2) );
  NAND2X0 P2_lt_696_U1 ( .IN1(P2_lt_696_n1), .IN2(P2_lt_696_n2), .QN(P2_N5203)
         );
  NOR2X0 P2_lt_696_U114 ( .QN(P2_lt_696_n142), .IN1(P2_N5009), 
        .IN2(P2_lt_696_n143) );
  NOR2X0 P2_lt_696_U113 ( .QN(P2_lt_696_n139), .IN1(P2_lt_696_n141), 
        .IN2(P2_lt_696_n142) );
  INVX0 P2_lt_696_U112 ( .ZN(P2_lt_696_n138), .INP(P2_N5325) );
  OR2X1 P2_lt_696_U111 ( .IN2(P2_N5010), .IN1(P2_lt_696_n138), 
        .Q(P2_lt_696_n140) );
  NAND2X0 P2_lt_696_U110 ( .IN1(P2_lt_696_n139), .IN2(P2_lt_696_n140), 
        .QN(P2_lt_696_n136) );
  NAND2X0 P2_lt_696_U109 ( .IN1(P2_N5010), .IN2(P2_lt_696_n138), 
        .QN(P2_lt_696_n137) );
  NAND2X0 P2_lt_696_U108 ( .IN1(P2_lt_696_n136), .IN2(P2_lt_696_n137), 
        .QN(P2_lt_696_n135) );
  NOR2X0 P2_lt_696_U107 ( .QN(P2_lt_696_n131), .IN1(P2_lt_696_n134), 
        .IN2(P2_lt_696_n135) );
  NOR2X0 P2_lt_696_U106 ( .QN(P2_lt_696_n132), .IN1(P2_N5011), 
        .IN2(P2_lt_696_n133) );
  NOR2X0 P2_lt_696_U105 ( .QN(P2_lt_696_n129), .IN1(P2_lt_696_n131), 
        .IN2(P2_lt_696_n132) );
  INVX0 P2_lt_696_U104 ( .ZN(P2_lt_696_n128), .INP(P2_N5327) );
  OR2X1 P2_lt_696_U103 ( .IN2(P2_N5012), .IN1(P2_lt_696_n128), 
        .Q(P2_lt_696_n130) );
  NAND2X0 P2_lt_696_U102 ( .IN1(P2_lt_696_n129), .IN2(P2_lt_696_n130), 
        .QN(P2_lt_696_n126) );
  NAND2X0 P2_lt_696_U101 ( .IN1(P2_N5012), .IN2(P2_lt_696_n128), 
        .QN(P2_lt_696_n127) );
  NAND2X0 P2_lt_696_U100 ( .IN1(P2_lt_696_n126), .IN2(P2_lt_696_n127), 
        .QN(P2_lt_696_n125) );
  NOR2X0 P2_lt_696_U99 ( .QN(P2_lt_696_n121), .IN1(P2_lt_696_n124), 
        .IN2(P2_lt_696_n125) );
  NOR2X0 P2_lt_696_U98 ( .QN(P2_lt_696_n122), .IN1(P2_N5013), 
        .IN2(P2_lt_696_n123) );
  NOR2X0 P2_lt_696_U97 ( .QN(P2_lt_696_n119), .IN1(P2_lt_696_n121), 
        .IN2(P2_lt_696_n122) );
  INVX0 P2_lt_696_U96 ( .ZN(P2_lt_696_n118), .INP(P2_N5329) );
  OR2X1 P2_lt_696_U95 ( .IN2(P2_N5014), .IN1(P2_lt_696_n118), 
        .Q(P2_lt_696_n120) );
  NAND2X0 P2_lt_696_U94 ( .IN1(P2_lt_696_n119), .IN2(P2_lt_696_n120), 
        .QN(P2_lt_696_n116) );
  NAND2X0 P2_lt_696_U93 ( .IN1(P2_N5014), .IN2(P2_lt_696_n118), 
        .QN(P2_lt_696_n117) );
  NAND2X0 P2_lt_696_U92 ( .IN1(P2_lt_696_n116), .IN2(P2_lt_696_n117), 
        .QN(P2_lt_696_n115) );
  NOR2X0 P2_lt_696_U91 ( .QN(P2_lt_696_n112), .IN1(P2_lt_696_n114), 
        .IN2(P2_lt_696_n115) );
  INVX0 P2_lt_696_U90 ( .ZN(P2_lt_696_n108), .INP(P2_N5331) );
  NOR2X0 P2_lt_696_U89 ( .QN(P2_lt_696_n113), .IN1(P2_N5016), 
        .IN2(P2_lt_696_n108) );
  NOR2X0 P2_lt_696_U88 ( .QN(P2_lt_696_n109), .IN1(P2_lt_696_n112), 
        .IN2(P2_lt_696_n113) );
  NAND2X0 P2_lt_696_U87 ( .IN1(P2_N5330), .IN2(n7275), .QN(P2_lt_696_n110) );
  NAND2X0 P2_lt_696_U86 ( .IN1(P2_lt_696_n109), .IN2(P2_lt_696_n110), 
        .QN(P2_lt_696_n106) );
  NAND2X0 P2_lt_696_U85 ( .IN1(P2_N5016), .IN2(P2_lt_696_n108), 
        .QN(P2_lt_696_n107) );
  NAND2X0 P2_lt_696_U84 ( .IN1(P2_lt_696_n106), .IN2(P2_lt_696_n107), 
        .QN(P2_lt_696_n105) );
  NOR2X0 P2_lt_696_U83 ( .QN(P2_lt_696_n101), .IN1(P2_lt_696_n104), 
        .IN2(P2_lt_696_n105) );
  NOR2X0 P2_lt_696_U82 ( .QN(P2_lt_696_n102), .IN1(P2_N5017), 
        .IN2(P2_lt_696_n103) );
  NOR2X0 P2_lt_696_U81 ( .QN(P2_lt_696_n99), .IN1(P2_lt_696_n101), 
        .IN2(P2_lt_696_n102) );
  INVX0 P2_lt_696_U80 ( .ZN(P2_lt_696_n98), .INP(P2_N5333) );
  OR2X1 P2_lt_696_U79 ( .IN2(P2_N5018), .IN1(P2_lt_696_n98), 
        .Q(P2_lt_696_n100) );
  NAND2X0 P2_lt_696_U78 ( .IN1(P2_lt_696_n99), .IN2(P2_lt_696_n100), 
        .QN(P2_lt_696_n96) );
  NAND2X0 P2_lt_696_U77 ( .IN1(P2_N5018), .IN2(P2_lt_696_n98), 
        .QN(P2_lt_696_n97) );
  NAND2X0 P2_lt_696_U76 ( .IN1(P2_lt_696_n96), .IN2(P2_lt_696_n97), 
        .QN(P2_lt_696_n95) );
  NOR2X0 P2_lt_696_U75 ( .QN(P2_lt_696_n91), .IN1(P2_lt_696_n94), 
        .IN2(P2_lt_696_n95) );
  NOR2X0 P2_lt_696_U74 ( .QN(P2_lt_696_n92), .IN1(P2_N5019), 
        .IN2(P2_lt_696_n93) );
  NOR2X0 P2_lt_696_U73 ( .QN(P2_lt_696_n89), .IN1(P2_lt_696_n91), 
        .IN2(P2_lt_696_n92) );
  INVX0 P2_lt_696_U72 ( .ZN(P2_lt_696_n88), .INP(P2_N5335) );
  OR2X1 P2_lt_696_U71 ( .IN2(P2_N5020), .IN1(P2_lt_696_n88), .Q(P2_lt_696_n90)
         );
  NAND2X0 P2_lt_696_U70 ( .IN1(P2_lt_696_n89), .IN2(P2_lt_696_n90), 
        .QN(P2_lt_696_n86) );
  NAND2X0 P2_lt_696_U69 ( .IN1(P2_N5020), .IN2(P2_lt_696_n88), 
        .QN(P2_lt_696_n87) );
  NAND2X0 P2_lt_696_U68 ( .IN1(P2_lt_696_n86), .IN2(P2_lt_696_n87), 
        .QN(P2_lt_696_n85) );
  NOR2X0 P2_lt_696_U67 ( .QN(P2_lt_696_n81), .IN1(P2_lt_696_n84), 
        .IN2(P2_lt_696_n85) );
  NOR2X0 P2_lt_696_U66 ( .QN(P2_lt_696_n82), .IN1(P2_N5021), 
        .IN2(P2_lt_696_n83) );
  NOR2X0 P2_lt_696_U65 ( .QN(P2_lt_696_n79), .IN1(P2_lt_696_n81), 
        .IN2(P2_lt_696_n82) );
  INVX0 P2_lt_696_U64 ( .ZN(P2_lt_696_n78), .INP(P2_N5337) );
  OR2X1 P2_lt_696_U63 ( .IN2(P2_N5022), .IN1(P2_lt_696_n78), .Q(P2_lt_696_n80)
         );
  NAND2X0 P2_lt_696_U62 ( .IN1(P2_lt_696_n79), .IN2(P2_lt_696_n80), 
        .QN(P2_lt_696_n76) );
  NAND2X0 P2_lt_696_U61 ( .IN1(P2_N5022), .IN2(P2_lt_696_n78), 
        .QN(P2_lt_696_n77) );
  NAND2X0 P2_lt_696_U60 ( .IN1(P2_lt_696_n76), .IN2(P2_lt_696_n77), 
        .QN(P2_lt_696_n75) );
  NOR2X0 P2_lt_696_U59 ( .QN(P2_lt_696_n71), .IN1(P2_lt_696_n74), 
        .IN2(P2_lt_696_n75) );
  NOR2X0 P2_lt_696_U58 ( .QN(P2_lt_696_n72), .IN1(P2_N5023), 
        .IN2(P2_lt_696_n73) );
  NOR2X0 P2_lt_696_U57 ( .QN(P2_lt_696_n69), .IN1(P2_lt_696_n71), 
        .IN2(P2_lt_696_n72) );
  INVX0 P2_lt_696_U56 ( .ZN(P2_lt_696_n68), .INP(P2_N5339) );
  OR2X1 P2_lt_696_U55 ( .IN2(P2_N5024), .IN1(P2_lt_696_n68), .Q(P2_lt_696_n70)
         );
  NAND2X0 P2_lt_696_U54 ( .IN1(P2_lt_696_n69), .IN2(P2_lt_696_n70), 
        .QN(P2_lt_696_n66) );
  NAND2X0 P2_lt_696_U53 ( .IN1(P2_N5024), .IN2(P2_lt_696_n68), 
        .QN(P2_lt_696_n67) );
  NAND2X0 P2_lt_696_U52 ( .IN1(P2_lt_696_n66), .IN2(P2_lt_696_n67), 
        .QN(P2_lt_696_n65) );
  NOR2X0 P2_lt_696_U51 ( .QN(P2_lt_696_n61), .IN1(P2_lt_696_n64), 
        .IN2(P2_lt_696_n65) );
  NOR2X0 P2_lt_696_U50 ( .QN(P2_lt_696_n62), .IN1(P2_N5025), 
        .IN2(P2_lt_696_n63) );
  NOR2X0 P2_lt_696_U49 ( .QN(P2_lt_696_n59), .IN1(P2_lt_696_n61), 
        .IN2(P2_lt_696_n62) );
  INVX0 P2_lt_696_U48 ( .ZN(P2_lt_696_n58), .INP(P2_N5341) );
  OR2X1 P2_lt_696_U47 ( .IN2(P2_N5026), .IN1(P2_lt_696_n58), .Q(P2_lt_696_n60)
         );
  NAND2X0 P2_lt_696_U46 ( .IN1(P2_lt_696_n59), .IN2(P2_lt_696_n60), 
        .QN(P2_lt_696_n56) );
  NAND2X0 P2_lt_696_U45 ( .IN1(P2_N5026), .IN2(P2_lt_696_n58), 
        .QN(P2_lt_696_n57) );
  NAND2X0 P2_lt_696_U44 ( .IN1(P2_lt_696_n56), .IN2(P2_lt_696_n57), 
        .QN(P2_lt_696_n55) );
  NOR2X0 P2_lt_696_U43 ( .QN(P2_lt_696_n51), .IN1(P2_lt_696_n54), 
        .IN2(P2_lt_696_n55) );
  NOR2X0 P2_lt_696_U42 ( .QN(P2_lt_696_n52), .IN1(P2_N5027), 
        .IN2(P2_lt_696_n53) );
  NOR2X0 P2_lt_696_U41 ( .QN(P2_lt_696_n49), .IN1(P2_lt_696_n51), 
        .IN2(P2_lt_696_n52) );
  INVX0 P2_lt_696_U40 ( .ZN(P2_lt_696_n48), .INP(P2_N5343) );
  OR2X1 P2_lt_696_U39 ( .IN2(P2_N5028), .IN1(P2_lt_696_n48), .Q(P2_lt_696_n50)
         );
  NAND2X0 P2_lt_696_U38 ( .IN1(P2_lt_696_n49), .IN2(P2_lt_696_n50), 
        .QN(P2_lt_696_n46) );
  NAND2X0 P2_lt_696_U37 ( .IN1(P2_N5028), .IN2(P2_lt_696_n48), 
        .QN(P2_lt_696_n47) );
  NAND2X0 P2_lt_696_U36 ( .IN1(P2_lt_696_n46), .IN2(P2_lt_696_n47), 
        .QN(P2_lt_696_n45) );
  NOR2X0 P2_lt_696_U35 ( .QN(P2_lt_696_n41), .IN1(P2_lt_696_n44), 
        .IN2(P2_lt_696_n45) );
  NOR2X0 P2_lt_696_U34 ( .QN(P2_lt_696_n42), .IN1(P2_N5029), 
        .IN2(P2_lt_696_n43) );
  NOR2X0 P2_lt_696_U33 ( .QN(P2_lt_696_n39), .IN1(P2_lt_696_n41), 
        .IN2(P2_lt_696_n42) );
  INVX0 P2_lt_696_U32 ( .ZN(P2_lt_696_n38), .INP(P2_N5345) );
  OR2X1 P2_lt_696_U31 ( .IN2(P2_N5030), .IN1(P2_lt_696_n38), .Q(P2_lt_696_n40)
         );
  NAND2X0 P2_lt_696_U30 ( .IN1(P2_lt_696_n39), .IN2(P2_lt_696_n40), 
        .QN(P2_lt_696_n36) );
  NAND2X0 P2_lt_696_U29 ( .IN1(P2_N5030), .IN2(P2_lt_696_n38), 
        .QN(P2_lt_696_n37) );
  NAND2X0 P2_lt_696_U28 ( .IN1(P2_lt_696_n36), .IN2(P2_lt_696_n37), 
        .QN(P2_lt_696_n35) );
  NOR2X0 P2_lt_696_U27 ( .QN(P2_lt_696_n31), .IN1(P2_lt_696_n34), 
        .IN2(P2_lt_696_n35) );
  NOR2X0 P2_lt_696_U26 ( .QN(P2_lt_696_n32), .IN1(P2_N5031), 
        .IN2(P2_lt_696_n33) );
  NOR2X0 P2_lt_696_U25 ( .QN(P2_lt_696_n29), .IN1(P2_lt_696_n31), 
        .IN2(P2_lt_696_n32) );
  INVX0 P2_lt_696_U24 ( .ZN(P2_lt_696_n28), .INP(P2_N5347) );
  OR2X1 P2_lt_696_U23 ( .IN2(P2_N5032), .IN1(P2_lt_696_n28), .Q(P2_lt_696_n30)
         );
  NAND2X0 P2_lt_696_U22 ( .IN1(P2_lt_696_n29), .IN2(P2_lt_696_n30), 
        .QN(P2_lt_696_n26) );
  INVX0 P2_lt_696_U157 ( .ZN(P2_lt_696_n5), .INP(P2_N5352) );
  OR2X1 P2_lt_696_U156 ( .IN2(P2_N5037), .IN1(P2_lt_696_n5), .Q(P2_lt_696_n1)
         );
  INVX0 P2_lt_696_U155 ( .ZN(P2_lt_696_n13), .INP(P2_N5350) );
  AND2X1 P2_lt_696_U154 ( .IN1(P2_lt_696_n13), .IN2(P2_N5035), 
        .Q(P2_lt_696_n14) );
  INVX0 P2_lt_696_U153 ( .ZN(P2_lt_696_n23), .INP(P2_N5348) );
  AND2X1 P2_lt_696_U152 ( .IN1(P2_lt_696_n23), .IN2(P2_N5033), 
        .Q(P2_lt_696_n24) );
  INVX0 P2_lt_696_U151 ( .ZN(P2_lt_696_n33), .INP(P2_N5346) );
  AND2X1 P2_lt_696_U150 ( .IN1(P2_lt_696_n33), .IN2(P2_N5031), 
        .Q(P2_lt_696_n34) );
  INVX0 P2_lt_696_U149 ( .ZN(P2_lt_696_n43), .INP(P2_N5344) );
  AND2X1 P2_lt_696_U148 ( .IN1(P2_lt_696_n43), .IN2(P2_N5029), 
        .Q(P2_lt_696_n44) );
  INVX0 P2_lt_696_U147 ( .ZN(P2_lt_696_n53), .INP(P2_N5342) );
  AND2X1 P2_lt_696_U146 ( .IN1(P2_lt_696_n53), .IN2(P2_N5027), 
        .Q(P2_lt_696_n54) );
  INVX0 P2_lt_696_U145 ( .ZN(P2_lt_696_n63), .INP(P2_N5340) );
  AND2X1 P2_lt_696_U144 ( .IN1(P2_lt_696_n63), .IN2(P2_N5025), 
        .Q(P2_lt_696_n64) );
  INVX0 P2_lt_696_U143 ( .ZN(P2_lt_696_n73), .INP(P2_N5338) );
  AND2X1 P2_lt_696_U142 ( .IN1(P2_lt_696_n73), .IN2(P2_N5023), 
        .Q(P2_lt_696_n74) );
  INVX0 P2_lt_696_U141 ( .ZN(P2_lt_696_n83), .INP(P2_N5336) );
  AND2X1 P2_lt_696_U140 ( .IN1(P2_lt_696_n83), .IN2(P2_N5021), 
        .Q(P2_lt_696_n84) );
  INVX0 P2_lt_696_U139 ( .ZN(P2_lt_696_n93), .INP(P2_N5334) );
  AND2X1 P2_lt_696_U138 ( .IN1(P2_lt_696_n93), .IN2(P2_N5019), 
        .Q(P2_lt_696_n94) );
  INVX0 P2_lt_696_U137 ( .ZN(P2_lt_696_n103), .INP(P2_N5332) );
  AND2X1 P2_lt_696_U136 ( .IN1(P2_lt_696_n103), .IN2(P2_N5017), 
        .Q(P2_lt_696_n104) );
  NOR2X0 P2_lt_696_U134 ( .QN(P2_lt_696_n114), .IN1(P2_N5330), .IN2(n7275) );
  INVX0 P2_lt_696_U133 ( .ZN(P2_lt_696_n123), .INP(P2_N5328) );
  AND2X1 P2_lt_696_U132 ( .IN1(P2_lt_696_n123), .IN2(P2_N5013), 
        .Q(P2_lt_696_n124) );
  INVX0 P2_lt_696_U131 ( .ZN(P2_lt_696_n133), .INP(P2_N5326) );
  AND2X1 P2_lt_696_U130 ( .IN1(P2_lt_696_n133), .IN2(P2_N5011), 
        .Q(P2_lt_696_n134) );
  INVX0 P2_lt_696_U129 ( .ZN(P2_lt_696_n143), .INP(P2_N5324) );
  AND2X1 P2_lt_696_U128 ( .IN1(P2_lt_696_n143), .IN2(P2_N5009), 
        .Q(P2_lt_696_n144) );
  INVX0 P2_lt_696_U127 ( .ZN(P2_lt_696_n154), .INP(P2_N5322) );
  INVX0 P2_lt_696_U126 ( .ZN(P2_lt_696_n156), .INP(P2_N5006) );
  NOR2X0 P2_lt_696_U125 ( .QN(P2_lt_696_n153), .IN1(P2_lt_696_n156), 
        .IN2(P2_N5321) );
  AND2X1 P2_lt_696_U124 ( .IN1(P2_lt_696_n154), .IN2(P2_lt_696_n153), 
        .Q(P2_lt_696_n155) );
  NOR2X0 P2_lt_696_U123 ( .QN(P2_lt_696_n151), .IN1(P2_N5007), 
        .IN2(P2_lt_696_n155) );
  NOR2X0 P2_lt_696_U122 ( .QN(P2_lt_696_n152), .IN1(P2_lt_696_n153), 
        .IN2(P2_lt_696_n154) );
  NOR2X0 P2_lt_696_U121 ( .QN(P2_lt_696_n149), .IN1(P2_lt_696_n151), 
        .IN2(P2_lt_696_n152) );
  INVX0 P2_lt_696_U120 ( .ZN(P2_lt_696_n148), .INP(P2_N5323) );
  OR2X1 P2_lt_696_U119 ( .IN2(P2_N5008), .IN1(P2_lt_696_n148), 
        .Q(P2_lt_696_n150) );
  NAND2X0 P2_lt_696_U118 ( .IN1(P2_lt_696_n149), .IN2(P2_lt_696_n150), 
        .QN(P2_lt_696_n146) );
  NAND2X0 P2_lt_696_U117 ( .IN1(P2_N5008), .IN2(P2_lt_696_n148), 
        .QN(P2_lt_696_n147) );
  NAND2X0 P2_lt_696_U116 ( .IN1(P2_lt_696_n146), .IN2(P2_lt_696_n147), 
        .QN(P2_lt_696_n145) );
  NOR2X0 P2_lt_696_U115 ( .QN(P2_lt_696_n141), .IN1(P2_lt_696_n144), 
        .IN2(P2_lt_696_n145) );
  NAND2X0 P2_lt_734_U85 ( .IN1(P2_N5016), .IN2(P2_lt_734_n108), 
        .QN(P2_lt_734_n107) );
  NAND2X0 P2_lt_734_U84 ( .IN1(P2_lt_734_n106), .IN2(P2_lt_734_n107), 
        .QN(P2_lt_734_n105) );
  NOR2X0 P2_lt_734_U83 ( .QN(P2_lt_734_n101), .IN1(P2_lt_734_n104), 
        .IN2(P2_lt_734_n105) );
  NOR2X0 P2_lt_734_U82 ( .QN(P2_lt_734_n102), .IN1(P2_N5017), 
        .IN2(P2_lt_734_n103) );
  NOR2X0 P2_lt_734_U81 ( .QN(P2_lt_734_n99), .IN1(P2_lt_734_n101), 
        .IN2(P2_lt_734_n102) );
  INVX0 P2_lt_734_U80 ( .ZN(P2_lt_734_n98), .INP(P2_N5333) );
  OR2X1 P2_lt_734_U79 ( .IN2(P2_N5018), .IN1(P2_lt_734_n98), 
        .Q(P2_lt_734_n100) );
  NAND2X0 P2_lt_734_U78 ( .IN1(P2_lt_734_n99), .IN2(P2_lt_734_n100), 
        .QN(P2_lt_734_n96) );
  NAND2X0 P2_lt_734_U77 ( .IN1(P2_N5018), .IN2(P2_lt_734_n98), 
        .QN(P2_lt_734_n97) );
  NAND2X0 P2_lt_734_U76 ( .IN1(P2_lt_734_n96), .IN2(P2_lt_734_n97), 
        .QN(P2_lt_734_n95) );
  NOR2X0 P2_lt_734_U75 ( .QN(P2_lt_734_n91), .IN1(P2_lt_734_n94), 
        .IN2(P2_lt_734_n95) );
  NOR2X0 P2_lt_734_U74 ( .QN(P2_lt_734_n92), .IN1(P2_N5019), 
        .IN2(P2_lt_734_n93) );
  NOR2X0 P2_lt_734_U73 ( .QN(P2_lt_734_n89), .IN1(P2_lt_734_n91), 
        .IN2(P2_lt_734_n92) );
  INVX0 P2_lt_734_U72 ( .ZN(P2_lt_734_n88), .INP(P2_N5335) );
  OR2X1 P2_lt_734_U71 ( .IN2(P2_N5020), .IN1(P2_lt_734_n88), .Q(P2_lt_734_n90)
         );
  NAND2X0 P2_lt_734_U70 ( .IN1(P2_lt_734_n89), .IN2(P2_lt_734_n90), 
        .QN(P2_lt_734_n86) );
  NAND2X0 P2_lt_734_U69 ( .IN1(P2_N5020), .IN2(P2_lt_734_n88), 
        .QN(P2_lt_734_n87) );
  NAND2X0 P2_lt_734_U68 ( .IN1(P2_lt_734_n86), .IN2(P2_lt_734_n87), 
        .QN(P2_lt_734_n85) );
  NOR2X0 P2_lt_734_U67 ( .QN(P2_lt_734_n81), .IN1(P2_lt_734_n84), 
        .IN2(P2_lt_734_n85) );
  NOR2X0 P2_lt_734_U66 ( .QN(P2_lt_734_n82), .IN1(P2_N5021), 
        .IN2(P2_lt_734_n83) );
  NOR2X0 P2_lt_734_U65 ( .QN(P2_lt_734_n79), .IN1(P2_lt_734_n81), 
        .IN2(P2_lt_734_n82) );
  INVX0 P2_lt_734_U64 ( .ZN(P2_lt_734_n78), .INP(P2_N5337) );
  OR2X1 P2_lt_734_U63 ( .IN2(P2_N5022), .IN1(P2_lt_734_n78), .Q(P2_lt_734_n80)
         );
  NAND2X0 P2_lt_734_U62 ( .IN1(P2_lt_734_n79), .IN2(P2_lt_734_n80), 
        .QN(P2_lt_734_n76) );
  NAND2X0 P2_lt_734_U61 ( .IN1(P2_N5022), .IN2(P2_lt_734_n78), 
        .QN(P2_lt_734_n77) );
  NAND2X0 P2_lt_734_U60 ( .IN1(P2_lt_734_n76), .IN2(P2_lt_734_n77), 
        .QN(P2_lt_734_n75) );
  NOR2X0 P2_lt_734_U59 ( .QN(P2_lt_734_n71), .IN1(P2_lt_734_n74), 
        .IN2(P2_lt_734_n75) );
  NOR2X0 P2_lt_734_U58 ( .QN(P2_lt_734_n72), .IN1(P2_N5023), 
        .IN2(P2_lt_734_n73) );
  NOR2X0 P2_lt_734_U57 ( .QN(P2_lt_734_n69), .IN1(P2_lt_734_n71), 
        .IN2(P2_lt_734_n72) );
  INVX0 P2_lt_734_U56 ( .ZN(P2_lt_734_n68), .INP(P2_N5339) );
  OR2X1 P2_lt_734_U55 ( .IN2(P2_N5024), .IN1(P2_lt_734_n68), .Q(P2_lt_734_n70)
         );
  NAND2X0 P2_lt_734_U54 ( .IN1(P2_lt_734_n69), .IN2(P2_lt_734_n70), 
        .QN(P2_lt_734_n66) );
  NAND2X0 P2_lt_734_U53 ( .IN1(P2_N5024), .IN2(P2_lt_734_n68), 
        .QN(P2_lt_734_n67) );
  NAND2X0 P2_lt_734_U52 ( .IN1(P2_lt_734_n66), .IN2(P2_lt_734_n67), 
        .QN(P2_lt_734_n65) );
  NOR2X0 P2_lt_734_U51 ( .QN(P2_lt_734_n61), .IN1(P2_lt_734_n64), 
        .IN2(P2_lt_734_n65) );
  NOR2X0 P2_lt_734_U50 ( .QN(P2_lt_734_n62), .IN1(P2_N5025), 
        .IN2(P2_lt_734_n63) );
  NOR2X0 P2_lt_734_U49 ( .QN(P2_lt_734_n59), .IN1(P2_lt_734_n61), 
        .IN2(P2_lt_734_n62) );
  INVX0 P2_lt_734_U48 ( .ZN(P2_lt_734_n58), .INP(P2_N5341) );
  OR2X1 P2_lt_734_U47 ( .IN2(P2_N5026), .IN1(P2_lt_734_n58), .Q(P2_lt_734_n60)
         );
  NAND2X0 P2_lt_734_U46 ( .IN1(P2_lt_734_n59), .IN2(P2_lt_734_n60), 
        .QN(P2_lt_734_n56) );
  NAND2X0 P2_lt_734_U45 ( .IN1(P2_N5026), .IN2(P2_lt_734_n58), 
        .QN(P2_lt_734_n57) );
  NAND2X0 P2_lt_734_U44 ( .IN1(P2_lt_734_n56), .IN2(P2_lt_734_n57), 
        .QN(P2_lt_734_n55) );
  NOR2X0 P2_lt_734_U43 ( .QN(P2_lt_734_n51), .IN1(P2_lt_734_n54), 
        .IN2(P2_lt_734_n55) );
  NOR2X0 P2_lt_734_U42 ( .QN(P2_lt_734_n52), .IN1(P2_N5027), 
        .IN2(P2_lt_734_n53) );
  NOR2X0 P2_lt_734_U41 ( .QN(P2_lt_734_n49), .IN1(P2_lt_734_n51), 
        .IN2(P2_lt_734_n52) );
  INVX0 P2_lt_734_U40 ( .ZN(P2_lt_734_n48), .INP(P2_N5343) );
  OR2X1 P2_lt_734_U39 ( .IN2(P2_N5028), .IN1(P2_lt_734_n48), .Q(P2_lt_734_n50)
         );
  NAND2X0 P2_lt_734_U38 ( .IN1(P2_lt_734_n49), .IN2(P2_lt_734_n50), 
        .QN(P2_lt_734_n46) );
  NAND2X0 P2_lt_734_U37 ( .IN1(P2_N5028), .IN2(P2_lt_734_n48), 
        .QN(P2_lt_734_n47) );
  NAND2X0 P2_lt_734_U36 ( .IN1(P2_lt_734_n46), .IN2(P2_lt_734_n47), 
        .QN(P2_lt_734_n45) );
  NOR2X0 P2_lt_734_U35 ( .QN(P2_lt_734_n41), .IN1(P2_lt_734_n44), 
        .IN2(P2_lt_734_n45) );
  NOR2X0 P2_lt_734_U34 ( .QN(P2_lt_734_n42), .IN1(P2_N5029), 
        .IN2(P2_lt_734_n43) );
  NOR2X0 P2_lt_734_U33 ( .QN(P2_lt_734_n39), .IN1(P2_lt_734_n41), 
        .IN2(P2_lt_734_n42) );
  INVX0 P2_lt_734_U32 ( .ZN(P2_lt_734_n38), .INP(P2_N5345) );
  OR2X1 P2_lt_734_U31 ( .IN2(P2_N5030), .IN1(P2_lt_734_n38), .Q(P2_lt_734_n40)
         );
  NAND2X0 P2_lt_734_U30 ( .IN1(P2_lt_734_n39), .IN2(P2_lt_734_n40), 
        .QN(P2_lt_734_n36) );
  NAND2X0 P2_lt_734_U29 ( .IN1(P2_N5030), .IN2(P2_lt_734_n38), 
        .QN(P2_lt_734_n37) );
  NAND2X0 P2_lt_734_U28 ( .IN1(P2_lt_734_n36), .IN2(P2_lt_734_n37), 
        .QN(P2_lt_734_n35) );
  NOR2X0 P2_lt_734_U27 ( .QN(P2_lt_734_n31), .IN1(P2_lt_734_n34), 
        .IN2(P2_lt_734_n35) );
  NOR2X0 P2_lt_734_U26 ( .QN(P2_lt_734_n32), .IN1(P2_N5031), 
        .IN2(P2_lt_734_n33) );
  NOR2X0 P2_lt_734_U25 ( .QN(P2_lt_734_n29), .IN1(P2_lt_734_n31), 
        .IN2(P2_lt_734_n32) );
  INVX0 P2_lt_734_U24 ( .ZN(P2_lt_734_n28), .INP(P2_N5347) );
  OR2X1 P2_lt_734_U23 ( .IN2(P2_N5032), .IN1(P2_lt_734_n28), .Q(P2_lt_734_n30)
         );
  NAND2X0 P2_lt_734_U22 ( .IN1(P2_lt_734_n29), .IN2(P2_lt_734_n30), 
        .QN(P2_lt_734_n26) );
  NAND2X0 P2_lt_734_U21 ( .IN1(P2_N5032), .IN2(P2_lt_734_n28), 
        .QN(P2_lt_734_n27) );
  NAND2X0 P2_lt_734_U20 ( .IN1(P2_lt_734_n26), .IN2(P2_lt_734_n27), 
        .QN(P2_lt_734_n25) );
  NOR2X0 P2_lt_734_U19 ( .QN(P2_lt_734_n21), .IN1(P2_lt_734_n24), 
        .IN2(P2_lt_734_n25) );
  NOR2X0 P2_lt_734_U18 ( .QN(P2_lt_734_n22), .IN1(P2_N5033), 
        .IN2(P2_lt_734_n23) );
  NOR2X0 P2_lt_734_U17 ( .QN(P2_lt_734_n19), .IN1(P2_lt_734_n21), 
        .IN2(P2_lt_734_n22) );
  INVX0 P2_lt_734_U16 ( .ZN(P2_lt_734_n18), .INP(P2_N5349) );
  OR2X1 P2_lt_734_U15 ( .IN2(P2_N5034), .IN1(P2_lt_734_n18), .Q(P2_lt_734_n20)
         );
  NAND2X0 P2_lt_734_U14 ( .IN1(P2_lt_734_n19), .IN2(P2_lt_734_n20), 
        .QN(P2_lt_734_n16) );
  NAND2X0 P2_lt_734_U13 ( .IN1(P2_N5034), .IN2(P2_lt_734_n18), 
        .QN(P2_lt_734_n17) );
  NAND2X0 P2_lt_734_U12 ( .IN1(P2_lt_734_n16), .IN2(P2_lt_734_n17), 
        .QN(P2_lt_734_n15) );
  NOR2X0 P2_lt_734_U11 ( .QN(P2_lt_734_n11), .IN1(P2_lt_734_n14), 
        .IN2(P2_lt_734_n15) );
  NOR2X0 P2_lt_734_U10 ( .QN(P2_lt_734_n12), .IN1(P2_N5035), 
        .IN2(P2_lt_734_n13) );
  NOR2X0 P2_lt_734_U9 ( .QN(P2_lt_734_n9), .IN1(P2_lt_734_n11), 
        .IN2(P2_lt_734_n12) );
  INVX0 P2_lt_734_U8 ( .ZN(P2_lt_734_n8), .INP(P2_N5351) );
  OR2X1 P2_lt_734_U7 ( .IN2(P2_N5036), .IN1(P2_lt_734_n8), .Q(P2_lt_734_n10)
         );
  NAND2X0 P2_lt_734_U6 ( .IN1(P2_lt_734_n9), .IN2(P2_lt_734_n10), 
        .QN(P2_lt_734_n6) );
  NAND2X0 P2_lt_734_U5 ( .IN1(P2_N5036), .IN2(P2_lt_734_n8), .QN(P2_lt_734_n7)
         );
  NAND2X0 P2_lt_734_U4 ( .IN1(P2_lt_734_n6), .IN2(P2_lt_734_n7), 
        .QN(P2_lt_734_n3) );
  NAND2X0 P2_lt_734_U3 ( .IN1(P2_N5037), .IN2(P2_lt_734_n5), .QN(P2_lt_734_n4)
         );
  NAND2X0 P2_lt_734_U2 ( .IN1(P2_lt_734_n3), .IN2(P2_lt_734_n4), 
        .QN(P2_lt_734_n2) );
  NAND2X0 P2_lt_734_U1 ( .IN1(P2_lt_734_n1), .IN2(P2_lt_734_n2), .QN(P2_N5284)
         );
  INVX0 P2_lt_734_U157 ( .ZN(P2_lt_734_n5), .INP(P2_N5352) );
  OR2X1 P2_lt_734_U156 ( .IN2(P2_N5037), .IN1(P2_lt_734_n5), .Q(P2_lt_734_n1)
         );
  INVX0 P2_lt_734_U155 ( .ZN(P2_lt_734_n13), .INP(P2_N5350) );
  AND2X1 P2_lt_734_U154 ( .IN1(P2_lt_734_n13), .IN2(P2_N5035), 
        .Q(P2_lt_734_n14) );
  INVX0 P2_lt_734_U153 ( .ZN(P2_lt_734_n23), .INP(P2_N5348) );
  AND2X1 P2_lt_734_U152 ( .IN1(P2_lt_734_n23), .IN2(P2_N5033), 
        .Q(P2_lt_734_n24) );
  INVX0 P2_lt_734_U151 ( .ZN(P2_lt_734_n33), .INP(P2_N5346) );
  AND2X1 P2_lt_734_U150 ( .IN1(P2_lt_734_n33), .IN2(P2_N5031), 
        .Q(P2_lt_734_n34) );
  INVX0 P2_lt_734_U149 ( .ZN(P2_lt_734_n43), .INP(P2_N5344) );
  AND2X1 P2_lt_734_U148 ( .IN1(P2_lt_734_n43), .IN2(P2_N5029), 
        .Q(P2_lt_734_n44) );
  INVX0 P2_lt_734_U147 ( .ZN(P2_lt_734_n53), .INP(P2_N5342) );
  AND2X1 P2_lt_734_U146 ( .IN1(P2_lt_734_n53), .IN2(P2_N5027), 
        .Q(P2_lt_734_n54) );
  INVX0 P2_lt_734_U145 ( .ZN(P2_lt_734_n63), .INP(P2_N5340) );
  AND2X1 P2_lt_734_U144 ( .IN1(P2_lt_734_n63), .IN2(P2_N5025), 
        .Q(P2_lt_734_n64) );
  INVX0 P2_lt_734_U143 ( .ZN(P2_lt_734_n73), .INP(P2_N5338) );
  AND2X1 P2_lt_734_U142 ( .IN1(P2_lt_734_n73), .IN2(P2_N5023), 
        .Q(P2_lt_734_n74) );
  INVX0 P2_lt_734_U141 ( .ZN(P2_lt_734_n83), .INP(P2_N5336) );
  AND2X1 P2_lt_734_U140 ( .IN1(P2_lt_734_n83), .IN2(P2_N5021), 
        .Q(P2_lt_734_n84) );
  INVX0 P2_lt_734_U139 ( .ZN(P2_lt_734_n93), .INP(P2_N5334) );
  AND2X1 P2_lt_734_U138 ( .IN1(P2_lt_734_n93), .IN2(P2_N5019), 
        .Q(P2_lt_734_n94) );
  INVX0 P2_lt_734_U137 ( .ZN(P2_lt_734_n103), .INP(P2_N5332) );
  AND2X1 P2_lt_734_U136 ( .IN1(P2_lt_734_n103), .IN2(P2_N5017), 
        .Q(P2_lt_734_n104) );
  NOR2X0 P2_lt_734_U134 ( .QN(P2_lt_734_n114), .IN1(P2_N5330), .IN2(n7275) );
  INVX0 P2_lt_734_U133 ( .ZN(P2_lt_734_n123), .INP(P2_N5328) );
  AND2X1 P2_lt_734_U132 ( .IN1(P2_lt_734_n123), .IN2(P2_N5013), 
        .Q(P2_lt_734_n124) );
  INVX0 P2_lt_734_U131 ( .ZN(P2_lt_734_n133), .INP(P2_N5326) );
  AND2X1 P2_lt_734_U130 ( .IN1(P2_lt_734_n133), .IN2(P2_N5011), 
        .Q(P2_lt_734_n134) );
  INVX0 P2_lt_734_U129 ( .ZN(P2_lt_734_n143), .INP(P2_N5324) );
  AND2X1 P2_lt_734_U128 ( .IN1(P2_lt_734_n143), .IN2(P2_N5009), 
        .Q(P2_lt_734_n144) );
  INVX0 P2_lt_734_U127 ( .ZN(P2_lt_734_n154), .INP(P2_N5322) );
  INVX0 P2_lt_734_U126 ( .ZN(P2_lt_734_n156), .INP(P2_N5006) );
  NOR2X0 P2_lt_734_U125 ( .QN(P2_lt_734_n153), .IN1(P2_lt_734_n156), 
        .IN2(P2_N5321) );
  AND2X1 P2_lt_734_U124 ( .IN1(P2_lt_734_n154), .IN2(P2_lt_734_n153), 
        .Q(P2_lt_734_n155) );
  NOR2X0 P2_lt_734_U123 ( .QN(P2_lt_734_n151), .IN1(P2_N5007), 
        .IN2(P2_lt_734_n155) );
  NOR2X0 P2_lt_734_U122 ( .QN(P2_lt_734_n152), .IN1(P2_lt_734_n153), 
        .IN2(P2_lt_734_n154) );
  NOR2X0 P2_lt_734_U121 ( .QN(P2_lt_734_n149), .IN1(P2_lt_734_n151), 
        .IN2(P2_lt_734_n152) );
  INVX0 P2_lt_734_U120 ( .ZN(P2_lt_734_n148), .INP(P2_N5323) );
  OR2X1 P2_lt_734_U119 ( .IN2(P2_N5008), .IN1(P2_lt_734_n148), 
        .Q(P2_lt_734_n150) );
  NAND2X0 P2_lt_734_U118 ( .IN1(P2_lt_734_n149), .IN2(P2_lt_734_n150), 
        .QN(P2_lt_734_n146) );
  NAND2X0 P2_lt_734_U117 ( .IN1(P2_N5008), .IN2(P2_lt_734_n148), 
        .QN(P2_lt_734_n147) );
  NAND2X0 P2_lt_734_U116 ( .IN1(P2_lt_734_n146), .IN2(P2_lt_734_n147), 
        .QN(P2_lt_734_n145) );
  NOR2X0 P2_lt_734_U115 ( .QN(P2_lt_734_n141), .IN1(P2_lt_734_n144), 
        .IN2(P2_lt_734_n145) );
  NOR2X0 P2_lt_734_U114 ( .QN(P2_lt_734_n142), .IN1(P2_N5009), 
        .IN2(P2_lt_734_n143) );
  NOR2X0 P2_lt_734_U113 ( .QN(P2_lt_734_n139), .IN1(P2_lt_734_n141), 
        .IN2(P2_lt_734_n142) );
  INVX0 P2_lt_734_U112 ( .ZN(P2_lt_734_n138), .INP(P2_N5325) );
  OR2X1 P2_lt_734_U111 ( .IN2(P2_N5010), .IN1(P2_lt_734_n138), 
        .Q(P2_lt_734_n140) );
  NAND2X0 P2_lt_734_U110 ( .IN1(P2_lt_734_n139), .IN2(P2_lt_734_n140), 
        .QN(P2_lt_734_n136) );
  NAND2X0 P2_lt_734_U109 ( .IN1(P2_N5010), .IN2(P2_lt_734_n138), 
        .QN(P2_lt_734_n137) );
  NAND2X0 P2_lt_734_U108 ( .IN1(P2_lt_734_n136), .IN2(P2_lt_734_n137), 
        .QN(P2_lt_734_n135) );
  NOR2X0 P2_lt_734_U107 ( .QN(P2_lt_734_n131), .IN1(P2_lt_734_n134), 
        .IN2(P2_lt_734_n135) );
  NOR2X0 P2_lt_734_U106 ( .QN(P2_lt_734_n132), .IN1(P2_N5011), 
        .IN2(P2_lt_734_n133) );
  NOR2X0 P2_lt_734_U105 ( .QN(P2_lt_734_n129), .IN1(P2_lt_734_n131), 
        .IN2(P2_lt_734_n132) );
  INVX0 P2_lt_734_U104 ( .ZN(P2_lt_734_n128), .INP(P2_N5327) );
  OR2X1 P2_lt_734_U103 ( .IN2(P2_N5012), .IN1(P2_lt_734_n128), 
        .Q(P2_lt_734_n130) );
  NAND2X0 P2_lt_734_U102 ( .IN1(P2_lt_734_n129), .IN2(P2_lt_734_n130), 
        .QN(P2_lt_734_n126) );
  NAND2X0 P2_lt_734_U101 ( .IN1(P2_N5012), .IN2(P2_lt_734_n128), 
        .QN(P2_lt_734_n127) );
  NAND2X0 P2_lt_734_U100 ( .IN1(P2_lt_734_n126), .IN2(P2_lt_734_n127), 
        .QN(P2_lt_734_n125) );
  NOR2X0 P2_lt_734_U99 ( .QN(P2_lt_734_n121), .IN1(P2_lt_734_n124), 
        .IN2(P2_lt_734_n125) );
  NOR2X0 P2_lt_734_U98 ( .QN(P2_lt_734_n122), .IN1(P2_N5013), 
        .IN2(P2_lt_734_n123) );
  NOR2X0 P2_lt_734_U97 ( .QN(P2_lt_734_n119), .IN1(P2_lt_734_n121), 
        .IN2(P2_lt_734_n122) );
  INVX0 P2_lt_734_U96 ( .ZN(P2_lt_734_n118), .INP(P2_N5329) );
  OR2X1 P2_lt_734_U95 ( .IN2(P2_N5014), .IN1(P2_lt_734_n118), 
        .Q(P2_lt_734_n120) );
  NAND2X0 P2_lt_734_U94 ( .IN1(P2_lt_734_n119), .IN2(P2_lt_734_n120), 
        .QN(P2_lt_734_n116) );
  NAND2X0 P2_lt_734_U93 ( .IN1(P2_N5014), .IN2(P2_lt_734_n118), 
        .QN(P2_lt_734_n117) );
  NAND2X0 P2_lt_734_U92 ( .IN1(P2_lt_734_n116), .IN2(P2_lt_734_n117), 
        .QN(P2_lt_734_n115) );
  NOR2X0 P2_lt_734_U91 ( .QN(P2_lt_734_n112), .IN1(P2_lt_734_n114), 
        .IN2(P2_lt_734_n115) );
  INVX0 P2_lt_734_U90 ( .ZN(P2_lt_734_n108), .INP(P2_N5331) );
  NOR2X0 P2_lt_734_U89 ( .QN(P2_lt_734_n113), .IN1(P2_N5016), 
        .IN2(P2_lt_734_n108) );
  NOR2X0 P2_lt_734_U88 ( .QN(P2_lt_734_n109), .IN1(P2_lt_734_n112), 
        .IN2(P2_lt_734_n113) );
  NAND2X0 P2_lt_734_U87 ( .IN1(P2_N5330), .IN2(n7275), .QN(P2_lt_734_n110) );
  NAND2X0 P2_lt_734_U86 ( .IN1(P2_lt_734_n109), .IN2(P2_lt_734_n110), 
        .QN(P2_lt_734_n106) );
  INVX0 P2_lt_742_U56 ( .ZN(P2_lt_742_n68), .INP(P2_N5339) );
  OR2X1 P2_lt_742_U55 ( .IN2(P2_N5024), .IN1(P2_lt_742_n68), .Q(P2_lt_742_n70)
         );
  NAND2X0 P2_lt_742_U54 ( .IN1(P2_lt_742_n69), .IN2(P2_lt_742_n70), 
        .QN(P2_lt_742_n66) );
  NAND2X0 P2_lt_742_U53 ( .IN1(P2_N5024), .IN2(P2_lt_742_n68), 
        .QN(P2_lt_742_n67) );
  NAND2X0 P2_lt_742_U52 ( .IN1(P2_lt_742_n66), .IN2(P2_lt_742_n67), 
        .QN(P2_lt_742_n65) );
  NOR2X0 P2_lt_742_U51 ( .QN(P2_lt_742_n61), .IN1(P2_lt_742_n64), 
        .IN2(P2_lt_742_n65) );
  NOR2X0 P2_lt_742_U50 ( .QN(P2_lt_742_n62), .IN1(P2_N5025), 
        .IN2(P2_lt_742_n63) );
  NOR2X0 P2_lt_742_U49 ( .QN(P2_lt_742_n59), .IN1(P2_lt_742_n61), 
        .IN2(P2_lt_742_n62) );
  INVX0 P2_lt_742_U48 ( .ZN(P2_lt_742_n58), .INP(P2_N5341) );
  OR2X1 P2_lt_742_U47 ( .IN2(P2_N5026), .IN1(P2_lt_742_n58), .Q(P2_lt_742_n60)
         );
  NAND2X0 P2_lt_742_U46 ( .IN1(P2_lt_742_n59), .IN2(P2_lt_742_n60), 
        .QN(P2_lt_742_n56) );
  NAND2X0 P2_lt_742_U45 ( .IN1(P2_N5026), .IN2(P2_lt_742_n58), 
        .QN(P2_lt_742_n57) );
  NAND2X0 P2_lt_742_U44 ( .IN1(P2_lt_742_n56), .IN2(P2_lt_742_n57), 
        .QN(P2_lt_742_n55) );
  NOR2X0 P2_lt_742_U43 ( .QN(P2_lt_742_n51), .IN1(P2_lt_742_n54), 
        .IN2(P2_lt_742_n55) );
  NOR2X0 P2_lt_742_U42 ( .QN(P2_lt_742_n52), .IN1(P2_N5027), 
        .IN2(P2_lt_742_n53) );
  NOR2X0 P2_lt_742_U41 ( .QN(P2_lt_742_n49), .IN1(P2_lt_742_n51), 
        .IN2(P2_lt_742_n52) );
  INVX0 P2_lt_742_U40 ( .ZN(P2_lt_742_n48), .INP(P2_N5343) );
  OR2X1 P2_lt_742_U39 ( .IN2(P2_N5028), .IN1(P2_lt_742_n48), .Q(P2_lt_742_n50)
         );
  NAND2X0 P2_lt_742_U38 ( .IN1(P2_lt_742_n49), .IN2(P2_lt_742_n50), 
        .QN(P2_lt_742_n46) );
  NAND2X0 P2_lt_742_U37 ( .IN1(P2_N5028), .IN2(P2_lt_742_n48), 
        .QN(P2_lt_742_n47) );
  NAND2X0 P2_lt_742_U36 ( .IN1(P2_lt_742_n46), .IN2(P2_lt_742_n47), 
        .QN(P2_lt_742_n45) );
  NOR2X0 P2_lt_742_U35 ( .QN(P2_lt_742_n41), .IN1(P2_lt_742_n44), 
        .IN2(P2_lt_742_n45) );
  NOR2X0 P2_lt_742_U34 ( .QN(P2_lt_742_n42), .IN1(P2_N5029), 
        .IN2(P2_lt_742_n43) );
  NOR2X0 P2_lt_742_U33 ( .QN(P2_lt_742_n39), .IN1(P2_lt_742_n41), 
        .IN2(P2_lt_742_n42) );
  INVX0 P2_lt_742_U32 ( .ZN(P2_lt_742_n38), .INP(P2_N5345) );
  OR2X1 P2_lt_742_U31 ( .IN2(P2_N5030), .IN1(P2_lt_742_n38), .Q(P2_lt_742_n40)
         );
  NAND2X0 P2_lt_742_U30 ( .IN1(P2_lt_742_n39), .IN2(P2_lt_742_n40), 
        .QN(P2_lt_742_n36) );
  NAND2X0 P2_lt_742_U29 ( .IN1(P2_N5030), .IN2(P2_lt_742_n38), 
        .QN(P2_lt_742_n37) );
  NAND2X0 P2_lt_742_U28 ( .IN1(P2_lt_742_n36), .IN2(P2_lt_742_n37), 
        .QN(P2_lt_742_n35) );
  NOR2X0 P2_lt_742_U27 ( .QN(P2_lt_742_n31), .IN1(P2_lt_742_n34), 
        .IN2(P2_lt_742_n35) );
  NOR2X0 P2_lt_742_U26 ( .QN(P2_lt_742_n32), .IN1(P2_N5031), 
        .IN2(P2_lt_742_n33) );
  NOR2X0 P2_lt_742_U25 ( .QN(P2_lt_742_n29), .IN1(P2_lt_742_n31), 
        .IN2(P2_lt_742_n32) );
  INVX0 P2_lt_742_U24 ( .ZN(P2_lt_742_n28), .INP(P2_N5347) );
  OR2X1 P2_lt_742_U23 ( .IN2(P2_N5032), .IN1(P2_lt_742_n28), .Q(P2_lt_742_n30)
         );
  NAND2X0 P2_lt_742_U22 ( .IN1(P2_lt_742_n29), .IN2(P2_lt_742_n30), 
        .QN(P2_lt_742_n26) );
  NAND2X0 P2_lt_742_U21 ( .IN1(P2_N5032), .IN2(P2_lt_742_n28), 
        .QN(P2_lt_742_n27) );
  NAND2X0 P2_lt_742_U20 ( .IN1(P2_lt_742_n26), .IN2(P2_lt_742_n27), 
        .QN(P2_lt_742_n25) );
  NOR2X0 P2_lt_742_U19 ( .QN(P2_lt_742_n21), .IN1(P2_lt_742_n24), 
        .IN2(P2_lt_742_n25) );
  NOR2X0 P2_lt_742_U18 ( .QN(P2_lt_742_n22), .IN1(P2_N5033), 
        .IN2(P2_lt_742_n23) );
  NOR2X0 P2_lt_742_U17 ( .QN(P2_lt_742_n19), .IN1(P2_lt_742_n21), 
        .IN2(P2_lt_742_n22) );
  INVX0 P2_lt_742_U16 ( .ZN(P2_lt_742_n18), .INP(P2_N5349) );
  OR2X1 P2_lt_742_U15 ( .IN2(P2_N5034), .IN1(P2_lt_742_n18), .Q(P2_lt_742_n20)
         );
  NAND2X0 P2_lt_742_U14 ( .IN1(P2_lt_742_n19), .IN2(P2_lt_742_n20), 
        .QN(P2_lt_742_n16) );
  NAND2X0 P2_lt_742_U13 ( .IN1(P2_N5034), .IN2(P2_lt_742_n18), 
        .QN(P2_lt_742_n17) );
  NAND2X0 P2_lt_742_U12 ( .IN1(P2_lt_742_n16), .IN2(P2_lt_742_n17), 
        .QN(P2_lt_742_n15) );
  NOR2X0 P2_lt_742_U11 ( .QN(P2_lt_742_n11), .IN1(P2_lt_742_n14), 
        .IN2(P2_lt_742_n15) );
  NOR2X0 P2_lt_742_U10 ( .QN(P2_lt_742_n12), .IN1(P2_N5035), 
        .IN2(P2_lt_742_n13) );
  NOR2X0 P2_lt_742_U9 ( .QN(P2_lt_742_n9), .IN1(P2_lt_742_n11), 
        .IN2(P2_lt_742_n12) );
  INVX0 P2_lt_742_U8 ( .ZN(P2_lt_742_n8), .INP(P2_N5351) );
  OR2X1 P2_lt_742_U7 ( .IN2(P2_N5036), .IN1(P2_lt_742_n8), .Q(P2_lt_742_n10)
         );
  NAND2X0 P2_lt_742_U6 ( .IN1(P2_lt_742_n9), .IN2(P2_lt_742_n10), 
        .QN(P2_lt_742_n6) );
  NAND2X0 P2_lt_742_U5 ( .IN1(P2_N5036), .IN2(P2_lt_742_n8), .QN(P2_lt_742_n7)
         );
  NAND2X0 P2_lt_742_U4 ( .IN1(P2_lt_742_n6), .IN2(P2_lt_742_n7), 
        .QN(P2_lt_742_n3) );
  NAND2X0 P2_lt_742_U3 ( .IN1(P2_N5037), .IN2(P2_lt_742_n5), .QN(P2_lt_742_n4)
         );
  NAND2X0 P2_lt_742_U2 ( .IN1(P2_lt_742_n3), .IN2(P2_lt_742_n4), 
        .QN(P2_lt_742_n2) );
  NAND2X0 P2_lt_742_U1 ( .IN1(P2_lt_742_n1), .IN2(P2_lt_742_n2), .QN(P2_N5353)
         );
  INVX0 P2_lt_742_U149 ( .ZN(P2_lt_742_n43), .INP(P2_N5344) );
  AND2X1 P2_lt_742_U148 ( .IN1(P2_lt_742_n43), .IN2(P2_N5029), 
        .Q(P2_lt_742_n44) );
  INVX0 P2_lt_742_U147 ( .ZN(P2_lt_742_n53), .INP(P2_N5342) );
  AND2X1 P2_lt_742_U146 ( .IN1(P2_lt_742_n53), .IN2(P2_N5027), 
        .Q(P2_lt_742_n54) );
  INVX0 P2_lt_742_U145 ( .ZN(P2_lt_742_n63), .INP(P2_N5340) );
  AND2X1 P2_lt_742_U144 ( .IN1(P2_lt_742_n63), .IN2(P2_N5025), 
        .Q(P2_lt_742_n64) );
  INVX0 P2_lt_742_U143 ( .ZN(P2_lt_742_n73), .INP(P2_N5338) );
  AND2X1 P2_lt_742_U142 ( .IN1(P2_lt_742_n73), .IN2(P2_N5023), 
        .Q(P2_lt_742_n74) );
  INVX0 P2_lt_742_U141 ( .ZN(P2_lt_742_n83), .INP(P2_N5336) );
  AND2X1 P2_lt_742_U140 ( .IN1(P2_lt_742_n83), .IN2(P2_N5021), 
        .Q(P2_lt_742_n84) );
  INVX0 P2_lt_742_U139 ( .ZN(P2_lt_742_n93), .INP(P2_N5334) );
  AND2X1 P2_lt_742_U138 ( .IN1(P2_lt_742_n93), .IN2(P2_N5019), 
        .Q(P2_lt_742_n94) );
  INVX0 P2_lt_742_U137 ( .ZN(P2_lt_742_n103), .INP(P2_N5332) );
  AND2X1 P2_lt_742_U136 ( .IN1(P2_lt_742_n103), .IN2(P2_N5017), 
        .Q(P2_lt_742_n104) );
  NOR2X0 P2_lt_742_U134 ( .QN(P2_lt_742_n114), .IN1(P2_N5330), .IN2(n7275) );
  INVX0 P2_lt_742_U133 ( .ZN(P2_lt_742_n123), .INP(P2_N5328) );
  AND2X1 P2_lt_742_U132 ( .IN1(P2_lt_742_n123), .IN2(P2_N5013), 
        .Q(P2_lt_742_n124) );
  INVX0 P2_lt_742_U131 ( .ZN(P2_lt_742_n133), .INP(P2_N5326) );
  AND2X1 P2_lt_742_U130 ( .IN1(P2_lt_742_n133), .IN2(P2_N5011), 
        .Q(P2_lt_742_n134) );
  INVX0 P2_lt_742_U129 ( .ZN(P2_lt_742_n143), .INP(P2_N5324) );
  AND2X1 P2_lt_742_U128 ( .IN1(P2_lt_742_n143), .IN2(P2_N5009), 
        .Q(P2_lt_742_n144) );
  INVX0 P2_lt_742_U127 ( .ZN(P2_lt_742_n154), .INP(P2_N5322) );
  INVX0 P2_lt_742_U126 ( .ZN(P2_lt_742_n156), .INP(P2_N5006) );
  NOR2X0 P2_lt_742_U125 ( .QN(P2_lt_742_n153), .IN1(P2_lt_742_n156), 
        .IN2(P2_N5321) );
  AND2X1 P2_lt_742_U124 ( .IN1(P2_lt_742_n154), .IN2(P2_lt_742_n153), 
        .Q(P2_lt_742_n155) );
  NOR2X0 P2_lt_742_U123 ( .QN(P2_lt_742_n151), .IN1(P2_N5007), 
        .IN2(P2_lt_742_n155) );
  NOR2X0 P2_lt_742_U122 ( .QN(P2_lt_742_n152), .IN1(P2_lt_742_n153), 
        .IN2(P2_lt_742_n154) );
  NOR2X0 P2_lt_742_U121 ( .QN(P2_lt_742_n149), .IN1(P2_lt_742_n151), 
        .IN2(P2_lt_742_n152) );
  INVX0 P2_lt_742_U120 ( .ZN(P2_lt_742_n148), .INP(P2_N5323) );
  OR2X1 P2_lt_742_U119 ( .IN2(P2_N5008), .IN1(P2_lt_742_n148), 
        .Q(P2_lt_742_n150) );
  NAND2X0 P2_lt_742_U118 ( .IN1(P2_lt_742_n149), .IN2(P2_lt_742_n150), 
        .QN(P2_lt_742_n146) );
  NAND2X0 P2_lt_742_U117 ( .IN1(P2_N5008), .IN2(P2_lt_742_n148), 
        .QN(P2_lt_742_n147) );
  NAND2X0 P2_lt_742_U116 ( .IN1(P2_lt_742_n146), .IN2(P2_lt_742_n147), 
        .QN(P2_lt_742_n145) );
  NOR2X0 P2_lt_742_U115 ( .QN(P2_lt_742_n141), .IN1(P2_lt_742_n144), 
        .IN2(P2_lt_742_n145) );
  NOR2X0 P2_lt_742_U114 ( .QN(P2_lt_742_n142), .IN1(P2_N5009), 
        .IN2(P2_lt_742_n143) );
  NOR2X0 P2_lt_742_U113 ( .QN(P2_lt_742_n139), .IN1(P2_lt_742_n141), 
        .IN2(P2_lt_742_n142) );
  INVX0 P2_lt_742_U112 ( .ZN(P2_lt_742_n138), .INP(P2_N5325) );
  OR2X1 P2_lt_742_U111 ( .IN2(P2_N5010), .IN1(P2_lt_742_n138), 
        .Q(P2_lt_742_n140) );
  NAND2X0 P2_lt_742_U110 ( .IN1(P2_lt_742_n139), .IN2(P2_lt_742_n140), 
        .QN(P2_lt_742_n136) );
  NAND2X0 P2_lt_742_U109 ( .IN1(P2_N5010), .IN2(P2_lt_742_n138), 
        .QN(P2_lt_742_n137) );
  NAND2X0 P2_lt_742_U108 ( .IN1(P2_lt_742_n136), .IN2(P2_lt_742_n137), 
        .QN(P2_lt_742_n135) );
  NOR2X0 P2_lt_742_U107 ( .QN(P2_lt_742_n131), .IN1(P2_lt_742_n134), 
        .IN2(P2_lt_742_n135) );
  NOR2X0 P2_lt_742_U106 ( .QN(P2_lt_742_n132), .IN1(P2_N5011), 
        .IN2(P2_lt_742_n133) );
  NOR2X0 P2_lt_742_U105 ( .QN(P2_lt_742_n129), .IN1(P2_lt_742_n131), 
        .IN2(P2_lt_742_n132) );
  INVX0 P2_lt_742_U104 ( .ZN(P2_lt_742_n128), .INP(P2_N5327) );
  OR2X1 P2_lt_742_U103 ( .IN2(P2_N5012), .IN1(P2_lt_742_n128), 
        .Q(P2_lt_742_n130) );
  NAND2X0 P2_lt_742_U102 ( .IN1(P2_lt_742_n129), .IN2(P2_lt_742_n130), 
        .QN(P2_lt_742_n126) );
  NAND2X0 P2_lt_742_U101 ( .IN1(P2_N5012), .IN2(P2_lt_742_n128), 
        .QN(P2_lt_742_n127) );
  NAND2X0 P2_lt_742_U100 ( .IN1(P2_lt_742_n126), .IN2(P2_lt_742_n127), 
        .QN(P2_lt_742_n125) );
  NOR2X0 P2_lt_742_U99 ( .QN(P2_lt_742_n121), .IN1(P2_lt_742_n124), 
        .IN2(P2_lt_742_n125) );
  NOR2X0 P2_lt_742_U98 ( .QN(P2_lt_742_n122), .IN1(P2_N5013), 
        .IN2(P2_lt_742_n123) );
  NOR2X0 P2_lt_742_U97 ( .QN(P2_lt_742_n119), .IN1(P2_lt_742_n121), 
        .IN2(P2_lt_742_n122) );
  INVX0 P2_lt_742_U96 ( .ZN(P2_lt_742_n118), .INP(P2_N5329) );
  OR2X1 P2_lt_742_U95 ( .IN2(P2_N5014), .IN1(P2_lt_742_n118), 
        .Q(P2_lt_742_n120) );
  NAND2X0 P2_lt_742_U94 ( .IN1(P2_lt_742_n119), .IN2(P2_lt_742_n120), 
        .QN(P2_lt_742_n116) );
  NAND2X0 P2_lt_742_U93 ( .IN1(P2_N5014), .IN2(P2_lt_742_n118), 
        .QN(P2_lt_742_n117) );
  NAND2X0 P2_lt_742_U92 ( .IN1(P2_lt_742_n116), .IN2(P2_lt_742_n117), 
        .QN(P2_lt_742_n115) );
  NOR2X0 P2_lt_742_U91 ( .QN(P2_lt_742_n112), .IN1(P2_lt_742_n114), 
        .IN2(P2_lt_742_n115) );
  INVX0 P2_lt_742_U90 ( .ZN(P2_lt_742_n108), .INP(P2_N5331) );
  NOR2X0 P2_lt_742_U89 ( .QN(P2_lt_742_n113), .IN1(P2_N5016), 
        .IN2(P2_lt_742_n108) );
  NOR2X0 P2_lt_742_U88 ( .QN(P2_lt_742_n109), .IN1(P2_lt_742_n112), 
        .IN2(P2_lt_742_n113) );
  NAND2X0 P2_lt_742_U87 ( .IN1(P2_N5330), .IN2(n7275), .QN(P2_lt_742_n110) );
  NAND2X0 P2_lt_742_U86 ( .IN1(P2_lt_742_n109), .IN2(P2_lt_742_n110), 
        .QN(P2_lt_742_n106) );
  NAND2X0 P2_lt_742_U85 ( .IN1(P2_N5016), .IN2(P2_lt_742_n108), 
        .QN(P2_lt_742_n107) );
  NAND2X0 P2_lt_742_U84 ( .IN1(P2_lt_742_n106), .IN2(P2_lt_742_n107), 
        .QN(P2_lt_742_n105) );
  NOR2X0 P2_lt_742_U83 ( .QN(P2_lt_742_n101), .IN1(P2_lt_742_n104), 
        .IN2(P2_lt_742_n105) );
  NOR2X0 P2_lt_742_U82 ( .QN(P2_lt_742_n102), .IN1(P2_N5017), 
        .IN2(P2_lt_742_n103) );
  NOR2X0 P2_lt_742_U81 ( .QN(P2_lt_742_n99), .IN1(P2_lt_742_n101), 
        .IN2(P2_lt_742_n102) );
  INVX0 P2_lt_742_U80 ( .ZN(P2_lt_742_n98), .INP(P2_N5333) );
  OR2X1 P2_lt_742_U79 ( .IN2(P2_N5018), .IN1(P2_lt_742_n98), 
        .Q(P2_lt_742_n100) );
  NAND2X0 P2_lt_742_U78 ( .IN1(P2_lt_742_n99), .IN2(P2_lt_742_n100), 
        .QN(P2_lt_742_n96) );
  NAND2X0 P2_lt_742_U77 ( .IN1(P2_N5018), .IN2(P2_lt_742_n98), 
        .QN(P2_lt_742_n97) );
  NAND2X0 P2_lt_742_U76 ( .IN1(P2_lt_742_n96), .IN2(P2_lt_742_n97), 
        .QN(P2_lt_742_n95) );
  NOR2X0 P2_lt_742_U75 ( .QN(P2_lt_742_n91), .IN1(P2_lt_742_n94), 
        .IN2(P2_lt_742_n95) );
  NOR2X0 P2_lt_742_U74 ( .QN(P2_lt_742_n92), .IN1(P2_N5019), 
        .IN2(P2_lt_742_n93) );
  NOR2X0 P2_lt_742_U73 ( .QN(P2_lt_742_n89), .IN1(P2_lt_742_n91), 
        .IN2(P2_lt_742_n92) );
  INVX0 P2_lt_742_U72 ( .ZN(P2_lt_742_n88), .INP(P2_N5335) );
  OR2X1 P2_lt_742_U71 ( .IN2(P2_N5020), .IN1(P2_lt_742_n88), .Q(P2_lt_742_n90)
         );
  NAND2X0 P2_lt_742_U70 ( .IN1(P2_lt_742_n89), .IN2(P2_lt_742_n90), 
        .QN(P2_lt_742_n86) );
  NAND2X0 P2_lt_742_U69 ( .IN1(P2_N5020), .IN2(P2_lt_742_n88), 
        .QN(P2_lt_742_n87) );
  NAND2X0 P2_lt_742_U68 ( .IN1(P2_lt_742_n86), .IN2(P2_lt_742_n87), 
        .QN(P2_lt_742_n85) );
  NOR2X0 P2_lt_742_U67 ( .QN(P2_lt_742_n81), .IN1(P2_lt_742_n84), 
        .IN2(P2_lt_742_n85) );
  NOR2X0 P2_lt_742_U66 ( .QN(P2_lt_742_n82), .IN1(P2_N5021), 
        .IN2(P2_lt_742_n83) );
  NOR2X0 P2_lt_742_U65 ( .QN(P2_lt_742_n79), .IN1(P2_lt_742_n81), 
        .IN2(P2_lt_742_n82) );
  INVX0 P2_lt_742_U64 ( .ZN(P2_lt_742_n78), .INP(P2_N5337) );
  OR2X1 P2_lt_742_U63 ( .IN2(P2_N5022), .IN1(P2_lt_742_n78), .Q(P2_lt_742_n80)
         );
  NAND2X0 P2_lt_742_U62 ( .IN1(P2_lt_742_n79), .IN2(P2_lt_742_n80), 
        .QN(P2_lt_742_n76) );
  NAND2X0 P2_lt_742_U61 ( .IN1(P2_N5022), .IN2(P2_lt_742_n78), 
        .QN(P2_lt_742_n77) );
  NAND2X0 P2_lt_742_U60 ( .IN1(P2_lt_742_n76), .IN2(P2_lt_742_n77), 
        .QN(P2_lt_742_n75) );
  NOR2X0 P2_lt_742_U59 ( .QN(P2_lt_742_n71), .IN1(P2_lt_742_n74), 
        .IN2(P2_lt_742_n75) );
  NOR2X0 P2_lt_742_U58 ( .QN(P2_lt_742_n72), .IN1(P2_N5023), 
        .IN2(P2_lt_742_n73) );
  NOR2X0 P2_lt_742_U57 ( .QN(P2_lt_742_n69), .IN1(P2_lt_742_n71), 
        .IN2(P2_lt_742_n72) );
  INVX0 P2_lt_742_U157 ( .ZN(P2_lt_742_n5), .INP(P2_N5352) );
  OR2X1 P2_lt_742_U156 ( .IN2(P2_N5037), .IN1(P2_lt_742_n5), .Q(P2_lt_742_n1)
         );
  INVX0 P2_lt_742_U155 ( .ZN(P2_lt_742_n13), .INP(P2_N5350) );
  AND2X1 P2_lt_742_U154 ( .IN1(P2_lt_742_n13), .IN2(P2_N5035), 
        .Q(P2_lt_742_n14) );
  INVX0 P2_lt_742_U153 ( .ZN(P2_lt_742_n23), .INP(P2_N5348) );
  AND2X1 P2_lt_742_U152 ( .IN1(P2_lt_742_n23), .IN2(P2_N5033), 
        .Q(P2_lt_742_n24) );
  INVX0 P2_lt_742_U151 ( .ZN(P2_lt_742_n33), .INP(P2_N5346) );
  AND2X1 P2_lt_742_U150 ( .IN1(P2_lt_742_n33), .IN2(P2_N5031), 
        .Q(P2_lt_742_n34) );
  NAND2X0 P2_add_918_U93 ( .IN1(P2_add_918_n91), .IN2(P2_add_918_n92), 
        .QN(P2_add_918_n90) );
  NOR2X0 P2_add_918_U92 ( .QN(P2_add_918_n88), .IN1(P2_add_918_n87), 
        .IN2(P2_add_918_n90) );
  AND2X1 P2_add_918_U91 ( .IN1(P2_add_918_n87), .IN2(P2_add_918_n90), 
        .Q(P2_add_918_n89) );
  NOR2X0 P2_add_918_U90 ( .QN(P2_N2872), .IN1(P2_add_918_n88), 
        .IN2(P2_add_918_n89) );
  NAND2X0 P2_add_918_U89 ( .IN1(n7237), .IN2(P2_add_918_n87), 
        .QN(P2_add_918_n84) );
  OR2X1 P2_add_918_U88 ( .IN2(n7237), .IN1(P2_add_918_n87), .Q(P2_add_918_n86)
         );
  NAND2X0 P2_add_918_U87 ( .IN1(P2_N2630), .IN2(P2_add_918_n86), 
        .QN(P2_add_918_n85) );
  NAND2X0 P2_add_918_U86 ( .IN1(P2_add_918_n84), .IN2(P2_add_918_n85), 
        .QN(P2_add_918_n77) );
  OR2X1 P2_add_918_U84 ( .IN2(P2_N2631), .IN1(n7229), .Q(P2_add_918_n81) );
  NAND2X0 P2_add_918_U83 ( .IN1(P2_N2631), .IN2(n7229), .QN(P2_add_918_n82) );
  NAND2X0 P2_add_918_U82 ( .IN1(P2_add_918_n81), .IN2(P2_add_918_n82), 
        .QN(P2_add_918_n80) );
  NOR2X0 P2_add_918_U81 ( .QN(P2_add_918_n78), .IN1(P2_add_918_n77), 
        .IN2(P2_add_918_n80) );
  AND2X1 P2_add_918_U80 ( .IN1(P2_add_918_n77), .IN2(P2_add_918_n80), 
        .Q(P2_add_918_n79) );
  NOR2X0 P2_add_918_U79 ( .QN(P2_N2873), .IN1(P2_add_918_n78), 
        .IN2(P2_add_918_n79) );
  NAND2X0 P2_add_918_U78 ( .IN1(P2_N5097), .IN2(P2_add_918_n77), 
        .QN(P2_add_918_n74) );
  OR2X1 P2_add_918_U77 ( .IN2(P2_N5097), .IN1(P2_add_918_n77), 
        .Q(P2_add_918_n76) );
  NAND2X0 P2_add_918_U76 ( .IN1(P2_N2631), .IN2(P2_add_918_n76), 
        .QN(P2_add_918_n75) );
  NAND2X0 P2_add_918_U75 ( .IN1(P2_add_918_n74), .IN2(P2_add_918_n75), 
        .QN(P2_add_918_n64) );
  OR2X1 P2_add_918_U73 ( .IN2(P2_N2632), .IN1(n7224), .Q(P2_add_918_n71) );
  NAND2X0 P2_add_918_U72 ( .IN1(P2_N2632), .IN2(n7224), .QN(P2_add_918_n72) );
  NAND2X0 P2_add_918_U71 ( .IN1(P2_add_918_n71), .IN2(P2_add_918_n72), 
        .QN(P2_add_918_n70) );
  NOR2X0 P2_add_918_U70 ( .QN(P2_add_918_n68), .IN1(P2_add_918_n64), 
        .IN2(P2_add_918_n70) );
  AND2X1 P2_add_918_U69 ( .IN1(P2_add_918_n64), .IN2(P2_add_918_n70), 
        .Q(P2_add_918_n69) );
  NOR2X0 P2_add_918_U68 ( .QN(P2_N2874), .IN1(P2_add_918_n68), 
        .IN2(P2_add_918_n69) );
  OR2X1 P2_add_918_U66 ( .IN2(P2_N2633), .IN1(n7222), .Q(P2_add_918_n65) );
  NAND2X0 P2_add_918_U65 ( .IN1(P2_N2633), .IN2(n7222), .QN(P2_add_918_n66) );
  NAND2X0 P2_add_918_U64 ( .IN1(P2_add_918_n65), .IN2(P2_add_918_n66), 
        .QN(P2_add_918_n60) );
  NAND2X0 P2_add_918_U63 ( .IN1(P2_N5098), .IN2(P2_add_918_n64), 
        .QN(P2_add_918_n61) );
  OR2X1 P2_add_918_U62 ( .IN2(P2_N5098), .IN1(P2_add_918_n64), 
        .Q(P2_add_918_n63) );
  NAND2X0 P2_add_918_U61 ( .IN1(P2_N2632), .IN2(P2_add_918_n63), 
        .QN(P2_add_918_n62) );
  NAND2X0 P2_add_918_U60 ( .IN1(P2_add_918_n61), .IN2(P2_add_918_n62), 
        .QN(P2_add_918_n59) );
  NOR2X0 P2_add_918_U59 ( .QN(P2_add_918_n57), .IN1(P2_add_918_n60), 
        .IN2(P2_add_918_n59) );
  AND2X1 P2_add_918_U58 ( .IN1(P2_add_918_n59), .IN2(P2_add_918_n60), 
        .Q(P2_add_918_n58) );
  NOR2X0 P2_add_918_U57 ( .QN(P2_N2875), .IN1(P2_add_918_n57), 
        .IN2(P2_add_918_n58) );
  OR2X1 P2_add_918_U55 ( .IN2(P2_N2607), .IN1(n7182), .Q(P2_add_918_n54) );
  NAND2X0 P2_add_918_U54 ( .IN1(P2_N2607), .IN2(n7182), .QN(P2_add_918_n55) );
  NAND2X0 P2_add_918_U53 ( .IN1(P2_add_918_n54), .IN2(P2_add_918_n55), 
        .QN(P2_add_918_n53) );
  NOR2X0 P2_add_918_U52 ( .QN(P2_add_918_n50), .IN1(P2_add_918_n52), 
        .IN2(P2_add_918_n53) );
  AND2X1 P2_add_918_U51 ( .IN1(P2_add_918_n52), .IN2(P2_add_918_n53), 
        .Q(P2_add_918_n51) );
  NOR2X0 P2_add_918_U50 ( .QN(P2_N2849), .IN1(P2_add_918_n50), 
        .IN2(P2_add_918_n51) );
  OR2X1 P2_add_918_U48 ( .IN2(P2_N2608), .IN1(n7178), .Q(P2_add_918_n47) );
  NAND2X0 P2_add_918_U47 ( .IN1(P2_N2608), .IN2(n7178), .QN(P2_add_918_n48) );
  NAND2X0 P2_add_918_U46 ( .IN1(P2_add_918_n47), .IN2(P2_add_918_n48), 
        .QN(P2_add_918_n46) );
  NOR2X0 P2_add_918_U45 ( .QN(P2_add_918_n43), .IN1(P2_add_918_n45), 
        .IN2(P2_add_918_n46) );
  AND2X1 P2_add_918_U44 ( .IN1(P2_add_918_n45), .IN2(P2_add_918_n46), 
        .Q(P2_add_918_n44) );
  NOR2X0 P2_add_918_U43 ( .QN(P2_N2850), .IN1(P2_add_918_n43), 
        .IN2(P2_add_918_n44) );
  OR2X1 P2_add_918_U41 ( .IN2(P2_N2609), .IN1(n7174), .Q(P2_add_918_n40) );
  NAND2X0 P2_add_918_U40 ( .IN1(P2_N2609), .IN2(n7174), .QN(P2_add_918_n41) );
  NAND2X0 P2_add_918_U39 ( .IN1(P2_add_918_n40), .IN2(P2_add_918_n41), 
        .QN(P2_add_918_n39) );
  NOR2X0 P2_add_918_U38 ( .QN(P2_add_918_n36), .IN1(P2_add_918_n38), 
        .IN2(P2_add_918_n39) );
  AND2X1 P2_add_918_U37 ( .IN1(P2_add_918_n38), .IN2(P2_add_918_n39), 
        .Q(P2_add_918_n37) );
  NOR2X0 P2_add_918_U36 ( .QN(P2_N2851), .IN1(P2_add_918_n36), 
        .IN2(P2_add_918_n37) );
  OR2X1 P2_add_918_U34 ( .IN2(P2_N2610), .IN1(n7166), .Q(P2_add_918_n33) );
  NAND2X0 P2_add_918_U33 ( .IN1(P2_N2610), .IN2(n7166), .QN(P2_add_918_n34) );
  NAND2X0 P2_add_918_U32 ( .IN1(P2_add_918_n33), .IN2(P2_add_918_n34), 
        .QN(P2_add_918_n32) );
  NOR2X0 P2_add_918_U31 ( .QN(P2_add_918_n29), .IN1(P2_add_918_n31), 
        .IN2(P2_add_918_n32) );
  AND2X1 P2_add_918_U30 ( .IN1(P2_add_918_n31), .IN2(P2_add_918_n32), 
        .Q(P2_add_918_n30) );
  NOR2X0 P2_add_918_U29 ( .QN(P2_N2852), .IN1(P2_add_918_n29), 
        .IN2(P2_add_918_n30) );
  OR2X1 P2_add_918_U27 ( .IN2(P2_N2611), .IN1(n7164), .Q(P2_add_918_n26) );
  NAND2X0 P2_add_918_U26 ( .IN1(P2_N2611), .IN2(n7164), .QN(P2_add_918_n27) );
  NAND2X0 P2_add_918_U25 ( .IN1(P2_add_918_n26), .IN2(P2_add_918_n27), 
        .QN(P2_add_918_n25) );
  NOR2X0 P2_add_918_U24 ( .QN(P2_add_918_n22), .IN1(P2_add_918_n24), 
        .IN2(P2_add_918_n25) );
  AND2X1 P2_add_918_U23 ( .IN1(P2_add_918_n24), .IN2(P2_add_918_n25), 
        .Q(P2_add_918_n23) );
  NOR2X0 P2_add_918_U22 ( .QN(P2_N2853), .IN1(P2_add_918_n22), 
        .IN2(P2_add_918_n23) );
  OR2X1 P2_add_918_U20 ( .IN2(P2_N2612), .IN1(n7157), .Q(P2_add_918_n19) );
  NAND2X0 P2_add_918_U19 ( .IN1(P2_N2612), .IN2(n7157), .QN(P2_add_918_n20) );
  NAND2X0 P2_add_918_U18 ( .IN1(P2_add_918_n19), .IN2(P2_add_918_n20), 
        .QN(P2_add_918_n18) );
  NOR2X0 P2_add_918_U17 ( .QN(P2_add_918_n15), .IN1(P2_add_918_n17), 
        .IN2(P2_add_918_n18) );
  AND2X1 P2_add_918_U16 ( .IN1(P2_add_918_n17), .IN2(P2_add_918_n18), 
        .Q(P2_add_918_n16) );
  NOR2X0 P2_add_918_U15 ( .QN(P2_N2854), .IN1(P2_add_918_n15), 
        .IN2(P2_add_918_n16) );
  OR2X1 P2_add_918_U13 ( .IN2(P2_N2613), .IN1(n7153), .Q(P2_add_918_n12) );
  NAND2X0 P2_add_918_U12 ( .IN1(P2_N2613), .IN2(n7153), .QN(P2_add_918_n13) );
  NAND2X0 P2_add_918_U11 ( .IN1(P2_add_918_n12), .IN2(P2_add_918_n13), 
        .QN(P2_add_918_n11) );
  NOR2X0 P2_add_918_U10 ( .QN(P2_add_918_n8), .IN1(P2_add_918_n10), 
        .IN2(P2_add_918_n11) );
  AND2X1 P2_add_918_U9 ( .IN1(P2_add_918_n10), .IN2(P2_add_918_n11), 
        .Q(P2_add_918_n9) );
  NOR2X0 P2_add_918_U8 ( .QN(P2_N2855), .IN1(P2_add_918_n8), 
        .IN2(P2_add_918_n9) );
  OR2X1 P2_add_918_U6 ( .IN2(P2_N2614), .IN1(n7149), .Q(P2_add_918_n5) );
  NAND2X0 P2_add_918_U5 ( .IN1(P2_N2614), .IN2(n7149), .QN(P2_add_918_n6) );
  NAND2X0 P2_add_918_U4 ( .IN1(P2_add_918_n5), .IN2(P2_add_918_n6), 
        .QN(P2_add_918_n4) );
  NOR2X0 P2_add_918_U3 ( .QN(P2_add_918_n1), .IN1(P2_add_918_n3), 
        .IN2(P2_add_918_n4) );
  AND2X1 P2_add_918_U2 ( .IN1(P2_add_918_n3), .IN2(P2_add_918_n4), 
        .Q(P2_add_918_n2) );
  NOR2X0 P2_add_918_U1 ( .QN(P2_N2856), .IN1(P2_add_918_n1), 
        .IN2(P2_add_918_n2) );
  NOR2X0 P2_add_918_U186 ( .QN(P2_add_918_n175), .IN1(P2_add_918_n174), 
        .IN2(P2_add_918_n177) );
  AND2X1 P2_add_918_U185 ( .IN1(P2_add_918_n174), .IN2(P2_add_918_n177), 
        .Q(P2_add_918_n176) );
  NOR2X0 P2_add_918_U184 ( .QN(P2_N2864), .IN1(P2_add_918_n175), 
        .IN2(P2_add_918_n176) );
  NAND2X0 P2_add_918_U183 ( .IN1(P2_N5088), .IN2(P2_add_918_n174), 
        .QN(P2_add_918_n171) );
  OR2X1 P2_add_918_U182 ( .IN2(P2_N5088), .IN1(P2_add_918_n174), 
        .Q(P2_add_918_n173) );
  NAND2X0 P2_add_918_U181 ( .IN1(P2_N2622), .IN2(P2_add_918_n173), 
        .QN(P2_add_918_n172) );
  NAND2X0 P2_add_918_U180 ( .IN1(P2_add_918_n171), .IN2(P2_add_918_n172), 
        .QN(P2_add_918_n164) );
  OR2X1 P2_add_918_U178 ( .IN2(P2_N2623), .IN1(n7188), .Q(P2_add_918_n168) );
  NAND2X0 P2_add_918_U177 ( .IN1(P2_N2623), .IN2(n7188), .QN(P2_add_918_n169)
         );
  NAND2X0 P2_add_918_U176 ( .IN1(P2_add_918_n168), .IN2(P2_add_918_n169), 
        .QN(P2_add_918_n167) );
  NOR2X0 P2_add_918_U175 ( .QN(P2_add_918_n165), .IN1(P2_add_918_n164), 
        .IN2(P2_add_918_n167) );
  AND2X1 P2_add_918_U174 ( .IN1(P2_add_918_n164), .IN2(P2_add_918_n167), 
        .Q(P2_add_918_n166) );
  NOR2X0 P2_add_918_U173 ( .QN(P2_N2865), .IN1(P2_add_918_n165), 
        .IN2(P2_add_918_n166) );
  NAND2X0 P2_add_918_U172 ( .IN1(n7187), .IN2(P2_add_918_n164), 
        .QN(P2_add_918_n161) );
  OR2X1 P2_add_918_U171 ( .IN2(n7187), .IN1(P2_add_918_n164), 
        .Q(P2_add_918_n163) );
  NAND2X0 P2_add_918_U170 ( .IN1(P2_N2623), .IN2(P2_add_918_n163), 
        .QN(P2_add_918_n162) );
  NAND2X0 P2_add_918_U169 ( .IN1(P2_add_918_n161), .IN2(P2_add_918_n162), 
        .QN(P2_add_918_n147) );
  OR2X1 P2_add_918_U167 ( .IN2(P2_N2624), .IN1(n7264), .Q(P2_add_918_n158) );
  NAND2X0 P2_add_918_U166 ( .IN1(P2_N2624), .IN2(n7264), .QN(P2_add_918_n159)
         );
  NAND2X0 P2_add_918_U165 ( .IN1(P2_add_918_n158), .IN2(P2_add_918_n159), 
        .QN(P2_add_918_n157) );
  NOR2X0 P2_add_918_U164 ( .QN(P2_add_918_n155), .IN1(P2_add_918_n147), 
        .IN2(P2_add_918_n157) );
  AND2X1 P2_add_918_U163 ( .IN1(P2_add_918_n147), .IN2(P2_add_918_n157), 
        .Q(P2_add_918_n156) );
  NOR2X0 P2_add_918_U162 ( .QN(P2_N2866), .IN1(P2_add_918_n155), 
        .IN2(P2_add_918_n156) );
  OR2X1 P2_add_918_U161 ( .IN2(P2_N2606), .IN1(n7186), .Q(P2_add_918_n152) );
  NAND2X0 P2_add_918_U160 ( .IN1(P2_N2606), .IN2(n7186), .QN(P2_add_918_n153)
         );
  NAND2X0 P2_add_918_U159 ( .IN1(P2_add_918_n152), .IN2(P2_add_918_n153), 
        .QN(P2_add_918_n150) );
  NAND2X0 P2_add_918_U158 ( .IN1(P2_add_918_n150), .IN2(P2_add_918_n151), 
        .QN(P2_add_918_n148) );
  OR2X1 P2_add_918_U157 ( .IN2(P2_add_918_n151), .IN1(P2_add_918_n150), 
        .Q(P2_add_918_n149) );
  NAND2X0 P2_add_918_U156 ( .IN1(P2_add_918_n148), .IN2(P2_add_918_n149), 
        .QN(P2_N2848) );
  NAND2X0 P2_add_918_U155 ( .IN1(n7263), .IN2(P2_add_918_n147), 
        .QN(P2_add_918_n144) );
  OR2X1 P2_add_918_U154 ( .IN2(n7263), .IN1(P2_add_918_n147), 
        .Q(P2_add_918_n146) );
  NAND2X0 P2_add_918_U153 ( .IN1(P2_N2624), .IN2(P2_add_918_n146), 
        .QN(P2_add_918_n145) );
  NAND2X0 P2_add_918_U152 ( .IN1(P2_add_918_n144), .IN2(P2_add_918_n145), 
        .QN(P2_add_918_n137) );
  OR2X1 P2_add_918_U150 ( .IN2(P2_N2625), .IN1(n7260), .Q(P2_add_918_n141) );
  NAND2X0 P2_add_918_U149 ( .IN1(P2_N2625), .IN2(n7260), .QN(P2_add_918_n142)
         );
  NAND2X0 P2_add_918_U148 ( .IN1(P2_add_918_n141), .IN2(P2_add_918_n142), 
        .QN(P2_add_918_n140) );
  NOR2X0 P2_add_918_U147 ( .QN(P2_add_918_n138), .IN1(P2_add_918_n137), 
        .IN2(P2_add_918_n140) );
  AND2X1 P2_add_918_U146 ( .IN1(P2_add_918_n137), .IN2(P2_add_918_n140), 
        .Q(P2_add_918_n139) );
  NOR2X0 P2_add_918_U145 ( .QN(P2_N2867), .IN1(P2_add_918_n138), 
        .IN2(P2_add_918_n139) );
  NAND2X0 P2_add_918_U144 ( .IN1(n7259), .IN2(P2_add_918_n137), 
        .QN(P2_add_918_n134) );
  OR2X1 P2_add_918_U143 ( .IN2(n7259), .IN1(P2_add_918_n137), 
        .Q(P2_add_918_n136) );
  NAND2X0 P2_add_918_U142 ( .IN1(P2_N2625), .IN2(P2_add_918_n136), 
        .QN(P2_add_918_n135) );
  NAND2X0 P2_add_918_U141 ( .IN1(P2_add_918_n134), .IN2(P2_add_918_n135), 
        .QN(P2_add_918_n127) );
  OR2X1 P2_add_918_U139 ( .IN2(P2_N2626), .IN1(n7253), .Q(P2_add_918_n131) );
  NAND2X0 P2_add_918_U138 ( .IN1(P2_N2626), .IN2(n7253), .QN(P2_add_918_n132)
         );
  NAND2X0 P2_add_918_U137 ( .IN1(P2_add_918_n131), .IN2(P2_add_918_n132), 
        .QN(P2_add_918_n130) );
  NOR2X0 P2_add_918_U136 ( .QN(P2_add_918_n128), .IN1(P2_add_918_n127), 
        .IN2(P2_add_918_n130) );
  AND2X1 P2_add_918_U135 ( .IN1(P2_add_918_n127), .IN2(P2_add_918_n130), 
        .Q(P2_add_918_n129) );
  NOR2X0 P2_add_918_U134 ( .QN(P2_N2868), .IN1(P2_add_918_n128), 
        .IN2(P2_add_918_n129) );
  NAND2X0 P2_add_918_U133 ( .IN1(n7252), .IN2(P2_add_918_n127), 
        .QN(P2_add_918_n124) );
  OR2X1 P2_add_918_U132 ( .IN2(n7252), .IN1(P2_add_918_n127), 
        .Q(P2_add_918_n126) );
  NAND2X0 P2_add_918_U131 ( .IN1(P2_N2626), .IN2(P2_add_918_n126), 
        .QN(P2_add_918_n125) );
  NAND2X0 P2_add_918_U130 ( .IN1(P2_add_918_n124), .IN2(P2_add_918_n125), 
        .QN(P2_add_918_n117) );
  OR2X1 P2_add_918_U128 ( .IN2(P2_N2627), .IN1(n7248), .Q(P2_add_918_n121) );
  NAND2X0 P2_add_918_U127 ( .IN1(P2_N2627), .IN2(n7248), .QN(P2_add_918_n122)
         );
  NAND2X0 P2_add_918_U126 ( .IN1(P2_add_918_n121), .IN2(P2_add_918_n122), 
        .QN(P2_add_918_n120) );
  NOR2X0 P2_add_918_U125 ( .QN(P2_add_918_n118), .IN1(P2_add_918_n117), 
        .IN2(P2_add_918_n120) );
  AND2X1 P2_add_918_U124 ( .IN1(P2_add_918_n117), .IN2(P2_add_918_n120), 
        .Q(P2_add_918_n119) );
  NOR2X0 P2_add_918_U123 ( .QN(P2_N2869), .IN1(P2_add_918_n118), 
        .IN2(P2_add_918_n119) );
  NAND2X0 P2_add_918_U122 ( .IN1(n7247), .IN2(P2_add_918_n117), 
        .QN(P2_add_918_n114) );
  OR2X1 P2_add_918_U121 ( .IN2(n7247), .IN1(P2_add_918_n117), 
        .Q(P2_add_918_n116) );
  NAND2X0 P2_add_918_U120 ( .IN1(P2_N2627), .IN2(P2_add_918_n116), 
        .QN(P2_add_918_n115) );
  NAND2X0 P2_add_918_U119 ( .IN1(P2_add_918_n114), .IN2(P2_add_918_n115), 
        .QN(P2_add_918_n107) );
  OR2X1 P2_add_918_U117 ( .IN2(P2_N2628), .IN1(n7243), .Q(P2_add_918_n111) );
  NAND2X0 P2_add_918_U116 ( .IN1(P2_N2628), .IN2(n7243), .QN(P2_add_918_n112)
         );
  NAND2X0 P2_add_918_U115 ( .IN1(P2_add_918_n111), .IN2(P2_add_918_n112), 
        .QN(P2_add_918_n110) );
  NOR2X0 P2_add_918_U114 ( .QN(P2_add_918_n108), .IN1(P2_add_918_n107), 
        .IN2(P2_add_918_n110) );
  AND2X1 P2_add_918_U113 ( .IN1(P2_add_918_n107), .IN2(P2_add_918_n110), 
        .Q(P2_add_918_n109) );
  NOR2X0 P2_add_918_U112 ( .QN(P2_N2870), .IN1(P2_add_918_n108), 
        .IN2(P2_add_918_n109) );
  NAND2X0 P2_add_918_U111 ( .IN1(P2_N5094), .IN2(P2_add_918_n107), 
        .QN(P2_add_918_n104) );
  OR2X1 P2_add_918_U110 ( .IN2(n7242), .IN1(P2_add_918_n107), 
        .Q(P2_add_918_n106) );
  NAND2X0 P2_add_918_U109 ( .IN1(P2_N2628), .IN2(P2_add_918_n106), 
        .QN(P2_add_918_n105) );
  NAND2X0 P2_add_918_U108 ( .IN1(P2_add_918_n104), .IN2(P2_add_918_n105), 
        .QN(P2_add_918_n97) );
  OR2X1 P2_add_918_U106 ( .IN2(P2_N2629), .IN1(n7239), .Q(P2_add_918_n101) );
  NAND2X0 P2_add_918_U105 ( .IN1(P2_N2629), .IN2(n7239), .QN(P2_add_918_n102)
         );
  NAND2X0 P2_add_918_U104 ( .IN1(P2_add_918_n101), .IN2(P2_add_918_n102), 
        .QN(P2_add_918_n100) );
  NOR2X0 P2_add_918_U103 ( .QN(P2_add_918_n98), .IN1(P2_add_918_n97), 
        .IN2(P2_add_918_n100) );
  AND2X1 P2_add_918_U102 ( .IN1(P2_add_918_n97), .IN2(P2_add_918_n100), 
        .Q(P2_add_918_n99) );
  NOR2X0 P2_add_918_U101 ( .QN(P2_N2871), .IN1(P2_add_918_n98), 
        .IN2(P2_add_918_n99) );
  NAND2X0 P2_add_918_U100 ( .IN1(n7238), .IN2(P2_add_918_n97), 
        .QN(P2_add_918_n94) );
  OR2X1 P2_add_918_U99 ( .IN2(n7238), .IN1(P2_add_918_n97), .Q(P2_add_918_n96)
         );
  NAND2X0 P2_add_918_U98 ( .IN1(P2_N2629), .IN2(P2_add_918_n96), 
        .QN(P2_add_918_n95) );
  NAND2X0 P2_add_918_U97 ( .IN1(P2_add_918_n94), .IN2(P2_add_918_n95), 
        .QN(P2_add_918_n87) );
  OR2X1 P2_add_918_U95 ( .IN2(P2_N2630), .IN1(n7234), .Q(P2_add_918_n91) );
  NAND2X0 P2_add_918_U94 ( .IN1(P2_N2630), .IN2(n7234), .QN(P2_add_918_n92) );
  NAND2X0 P2_add_918_U279 ( .IN1(n7158), .IN2(P2_add_918_n17), 
        .QN(P2_add_918_n257) );
  OR2X1 P2_add_918_U278 ( .IN2(n7158), .IN1(P2_add_918_n17), 
        .Q(P2_add_918_n259) );
  NAND2X0 P2_add_918_U277 ( .IN1(P2_N2612), .IN2(P2_add_918_n259), 
        .QN(P2_add_918_n258) );
  NAND2X0 P2_add_918_U276 ( .IN1(P2_add_918_n257), .IN2(P2_add_918_n258), 
        .QN(P2_add_918_n10) );
  NAND2X0 P2_add_918_U275 ( .IN1(P2_N5079), .IN2(P2_add_918_n10), 
        .QN(P2_add_918_n254) );
  OR2X1 P2_add_918_U274 ( .IN2(P2_N5079), .IN1(P2_add_918_n10), 
        .Q(P2_add_918_n256) );
  NAND2X0 P2_add_918_U273 ( .IN1(P2_N2613), .IN2(P2_add_918_n256), 
        .QN(P2_add_918_n255) );
  NAND2X0 P2_add_918_U272 ( .IN1(P2_add_918_n254), .IN2(P2_add_918_n255), 
        .QN(P2_add_918_n3) );
  NAND2X0 P2_add_918_U271 ( .IN1(P2_N5080), .IN2(P2_add_918_n3), 
        .QN(P2_add_918_n251) );
  OR2X1 P2_add_918_U270 ( .IN2(P2_N5080), .IN1(P2_add_918_n3), 
        .Q(P2_add_918_n253) );
  NAND2X0 P2_add_918_U269 ( .IN1(P2_N2614), .IN2(P2_add_918_n253), 
        .QN(P2_add_918_n252) );
  NAND2X0 P2_add_918_U268 ( .IN1(P2_add_918_n251), .IN2(P2_add_918_n252), 
        .QN(P2_add_918_n244) );
  OR2X1 P2_add_918_U266 ( .IN2(P2_N2615), .IN1(n7219), .Q(P2_add_918_n248) );
  NAND2X0 P2_add_918_U265 ( .IN1(P2_N2615), .IN2(n7219), .QN(P2_add_918_n249)
         );
  NAND2X0 P2_add_918_U264 ( .IN1(P2_add_918_n248), .IN2(P2_add_918_n249), 
        .QN(P2_add_918_n247) );
  NOR2X0 P2_add_918_U263 ( .QN(P2_add_918_n245), .IN1(P2_add_918_n244), 
        .IN2(P2_add_918_n247) );
  AND2X1 P2_add_918_U262 ( .IN1(P2_add_918_n244), .IN2(P2_add_918_n247), 
        .Q(P2_add_918_n246) );
  NOR2X0 P2_add_918_U261 ( .QN(P2_N2857), .IN1(P2_add_918_n245), 
        .IN2(P2_add_918_n246) );
  NAND2X0 P2_add_918_U260 ( .IN1(P2_N5081), .IN2(P2_add_918_n244), 
        .QN(P2_add_918_n241) );
  OR2X1 P2_add_918_U259 ( .IN2(P2_N5081), .IN1(P2_add_918_n244), 
        .Q(P2_add_918_n243) );
  NAND2X0 P2_add_918_U258 ( .IN1(P2_N2615), .IN2(P2_add_918_n243), 
        .QN(P2_add_918_n242) );
  NAND2X0 P2_add_918_U257 ( .IN1(P2_add_918_n241), .IN2(P2_add_918_n242), 
        .QN(P2_add_918_n234) );
  OR2X1 P2_add_918_U255 ( .IN2(P2_N2616), .IN1(n7214), .Q(P2_add_918_n238) );
  NAND2X0 P2_add_918_U254 ( .IN1(P2_N2616), .IN2(n7214), .QN(P2_add_918_n239)
         );
  NAND2X0 P2_add_918_U253 ( .IN1(P2_add_918_n238), .IN2(P2_add_918_n239), 
        .QN(P2_add_918_n237) );
  NOR2X0 P2_add_918_U252 ( .QN(P2_add_918_n235), .IN1(P2_add_918_n234), 
        .IN2(P2_add_918_n237) );
  AND2X1 P2_add_918_U251 ( .IN1(P2_add_918_n234), .IN2(P2_add_918_n237), 
        .Q(P2_add_918_n236) );
  NOR2X0 P2_add_918_U250 ( .QN(P2_N2858), .IN1(P2_add_918_n235), 
        .IN2(P2_add_918_n236) );
  NAND2X0 P2_add_918_U249 ( .IN1(n7216), .IN2(P2_add_918_n234), 
        .QN(P2_add_918_n231) );
  OR2X1 P2_add_918_U248 ( .IN2(n7216), .IN1(P2_add_918_n234), 
        .Q(P2_add_918_n233) );
  NAND2X0 P2_add_918_U247 ( .IN1(P2_N2616), .IN2(P2_add_918_n233), 
        .QN(P2_add_918_n232) );
  NAND2X0 P2_add_918_U246 ( .IN1(P2_add_918_n231), .IN2(P2_add_918_n232), 
        .QN(P2_add_918_n224) );
  OR2X1 P2_add_918_U244 ( .IN2(P2_N2617), .IN1(n7211), .Q(P2_add_918_n228) );
  NAND2X0 P2_add_918_U243 ( .IN1(P2_N2617), .IN2(n7211), .QN(P2_add_918_n229)
         );
  NAND2X0 P2_add_918_U242 ( .IN1(P2_add_918_n228), .IN2(P2_add_918_n229), 
        .QN(P2_add_918_n227) );
  NOR2X0 P2_add_918_U241 ( .QN(P2_add_918_n225), .IN1(P2_add_918_n224), 
        .IN2(P2_add_918_n227) );
  AND2X1 P2_add_918_U240 ( .IN1(P2_add_918_n224), .IN2(P2_add_918_n227), 
        .Q(P2_add_918_n226) );
  NOR2X0 P2_add_918_U239 ( .QN(P2_N2859), .IN1(P2_add_918_n225), 
        .IN2(P2_add_918_n226) );
  NAND2X0 P2_add_918_U238 ( .IN1(n7210), .IN2(P2_add_918_n224), 
        .QN(P2_add_918_n221) );
  OR2X1 P2_add_918_U237 ( .IN2(n7210), .IN1(P2_add_918_n224), 
        .Q(P2_add_918_n223) );
  NAND2X0 P2_add_918_U236 ( .IN1(P2_N2617), .IN2(P2_add_918_n223), 
        .QN(P2_add_918_n222) );
  NAND2X0 P2_add_918_U235 ( .IN1(P2_add_918_n221), .IN2(P2_add_918_n222), 
        .QN(P2_add_918_n214) );
  OR2X1 P2_add_918_U233 ( .IN2(P2_N2618), .IN1(n7208), .Q(P2_add_918_n218) );
  NAND2X0 P2_add_918_U232 ( .IN1(P2_N2618), .IN2(n7208), .QN(P2_add_918_n219)
         );
  NAND2X0 P2_add_918_U231 ( .IN1(P2_add_918_n218), .IN2(P2_add_918_n219), 
        .QN(P2_add_918_n217) );
  NOR2X0 P2_add_918_U230 ( .QN(P2_add_918_n215), .IN1(P2_add_918_n214), 
        .IN2(P2_add_918_n217) );
  AND2X1 P2_add_918_U229 ( .IN1(P2_add_918_n214), .IN2(P2_add_918_n217), 
        .Q(P2_add_918_n216) );
  NOR2X0 P2_add_918_U228 ( .QN(P2_N2860), .IN1(P2_add_918_n215), 
        .IN2(P2_add_918_n216) );
  NAND2X0 P2_add_918_U227 ( .IN1(P2_N5084), .IN2(P2_add_918_n214), 
        .QN(P2_add_918_n211) );
  OR2X1 P2_add_918_U226 ( .IN2(P2_N5084), .IN1(P2_add_918_n214), 
        .Q(P2_add_918_n213) );
  NAND2X0 P2_add_918_U225 ( .IN1(P2_N2618), .IN2(P2_add_918_n213), 
        .QN(P2_add_918_n212) );
  NAND2X0 P2_add_918_U224 ( .IN1(P2_add_918_n211), .IN2(P2_add_918_n212), 
        .QN(P2_add_918_n204) );
  OR2X1 P2_add_918_U222 ( .IN2(P2_N2619), .IN1(n7205), .Q(P2_add_918_n208) );
  NAND2X0 P2_add_918_U221 ( .IN1(P2_N2619), .IN2(n7205), .QN(P2_add_918_n209)
         );
  NAND2X0 P2_add_918_U220 ( .IN1(P2_add_918_n208), .IN2(P2_add_918_n209), 
        .QN(P2_add_918_n207) );
  NOR2X0 P2_add_918_U219 ( .QN(P2_add_918_n205), .IN1(P2_add_918_n204), 
        .IN2(P2_add_918_n207) );
  AND2X1 P2_add_918_U218 ( .IN1(P2_add_918_n204), .IN2(P2_add_918_n207), 
        .Q(P2_add_918_n206) );
  NOR2X0 P2_add_918_U217 ( .QN(P2_N2861), .IN1(P2_add_918_n205), 
        .IN2(P2_add_918_n206) );
  NAND2X0 P2_add_918_U216 ( .IN1(P2_N5085), .IN2(P2_add_918_n204), 
        .QN(P2_add_918_n201) );
  OR2X1 P2_add_918_U215 ( .IN2(P2_N5085), .IN1(P2_add_918_n204), 
        .Q(P2_add_918_n203) );
  NAND2X0 P2_add_918_U214 ( .IN1(P2_N2619), .IN2(P2_add_918_n203), 
        .QN(P2_add_918_n202) );
  NAND2X0 P2_add_918_U213 ( .IN1(P2_add_918_n201), .IN2(P2_add_918_n202), 
        .QN(P2_add_918_n194) );
  OR2X1 P2_add_918_U211 ( .IN2(P2_N2620), .IN1(n7201), .Q(P2_add_918_n198) );
  NAND2X0 P2_add_918_U210 ( .IN1(P2_N2620), .IN2(n7201), .QN(P2_add_918_n199)
         );
  NAND2X0 P2_add_918_U209 ( .IN1(P2_add_918_n198), .IN2(P2_add_918_n199), 
        .QN(P2_add_918_n197) );
  NOR2X0 P2_add_918_U208 ( .QN(P2_add_918_n195), .IN1(P2_add_918_n194), 
        .IN2(P2_add_918_n197) );
  AND2X1 P2_add_918_U207 ( .IN1(P2_add_918_n194), .IN2(P2_add_918_n197), 
        .Q(P2_add_918_n196) );
  NOR2X0 P2_add_918_U206 ( .QN(P2_N2862), .IN1(P2_add_918_n195), 
        .IN2(P2_add_918_n196) );
  NAND2X0 P2_add_918_U205 ( .IN1(n7202), .IN2(P2_add_918_n194), 
        .QN(P2_add_918_n191) );
  OR2X1 P2_add_918_U204 ( .IN2(n7202), .IN1(P2_add_918_n194), 
        .Q(P2_add_918_n193) );
  NAND2X0 P2_add_918_U203 ( .IN1(P2_N2620), .IN2(P2_add_918_n193), 
        .QN(P2_add_918_n192) );
  NAND2X0 P2_add_918_U202 ( .IN1(P2_add_918_n191), .IN2(P2_add_918_n192), 
        .QN(P2_add_918_n184) );
  OR2X1 P2_add_918_U200 ( .IN2(P2_N2621), .IN1(n7197), .Q(P2_add_918_n188) );
  NAND2X0 P2_add_918_U199 ( .IN1(P2_N2621), .IN2(n7197), .QN(P2_add_918_n189)
         );
  NAND2X0 P2_add_918_U198 ( .IN1(P2_add_918_n188), .IN2(P2_add_918_n189), 
        .QN(P2_add_918_n187) );
  NOR2X0 P2_add_918_U197 ( .QN(P2_add_918_n185), .IN1(P2_add_918_n184), 
        .IN2(P2_add_918_n187) );
  AND2X1 P2_add_918_U196 ( .IN1(P2_add_918_n184), .IN2(P2_add_918_n187), 
        .Q(P2_add_918_n186) );
  NOR2X0 P2_add_918_U195 ( .QN(P2_N2863), .IN1(P2_add_918_n185), 
        .IN2(P2_add_918_n186) );
  NAND2X0 P2_add_918_U194 ( .IN1(P2_N5087), .IN2(P2_add_918_n184), 
        .QN(P2_add_918_n181) );
  OR2X1 P2_add_918_U193 ( .IN2(P2_N5087), .IN1(P2_add_918_n184), 
        .Q(P2_add_918_n183) );
  NAND2X0 P2_add_918_U192 ( .IN1(P2_N2621), .IN2(P2_add_918_n183), 
        .QN(P2_add_918_n182) );
  NAND2X0 P2_add_918_U191 ( .IN1(P2_add_918_n181), .IN2(P2_add_918_n182), 
        .QN(P2_add_918_n174) );
  OR2X1 P2_add_918_U189 ( .IN2(P2_N2622), .IN1(n7195), .Q(P2_add_918_n178) );
  NAND2X0 P2_add_918_U188 ( .IN1(P2_N2622), .IN2(n7195), .QN(P2_add_918_n179)
         );
  NAND2X0 P2_add_918_U187 ( .IN1(P2_add_918_n178), .IN2(P2_add_918_n179), 
        .QN(P2_add_918_n177) );
  OR2X1 P2_add_918_U308 ( .IN2(P2_N2605), .IN1(n2919), .Q(P2_add_918_n278) );
  NAND2X0 P2_add_918_U307 ( .IN1(P2_N2605), .IN2(n2919), .QN(P2_add_918_n279)
         );
  NAND2X0 P2_add_918_U306 ( .IN1(P2_add_918_n278), .IN2(P2_add_918_n279), 
        .QN(P2_N2847) );
  NAND2X0 P2_add_918_U304 ( .IN1(P2_N2605), .IN2(n7035), .QN(P2_add_918_n151)
         );
  OR2X1 P2_add_918_U303 ( .IN2(P2_add_918_n151), .IN1(n7186), 
        .Q(P2_add_918_n275) );
  NAND2X0 P2_add_918_U302 ( .IN1(n7186), .IN2(P2_add_918_n151), 
        .QN(P2_add_918_n277) );
  NAND2X0 P2_add_918_U301 ( .IN1(P2_N2606), .IN2(P2_add_918_n277), 
        .QN(P2_add_918_n276) );
  NAND2X0 P2_add_918_U300 ( .IN1(P2_add_918_n275), .IN2(P2_add_918_n276), 
        .QN(P2_add_918_n52) );
  NAND2X0 P2_add_918_U299 ( .IN1(n7181), .IN2(P2_add_918_n52), 
        .QN(P2_add_918_n272) );
  OR2X1 P2_add_918_U298 ( .IN2(n7181), .IN1(P2_add_918_n52), 
        .Q(P2_add_918_n274) );
  NAND2X0 P2_add_918_U297 ( .IN1(P2_N2607), .IN2(P2_add_918_n274), 
        .QN(P2_add_918_n273) );
  NAND2X0 P2_add_918_U296 ( .IN1(P2_add_918_n272), .IN2(P2_add_918_n273), 
        .QN(P2_add_918_n45) );
  NAND2X0 P2_add_918_U295 ( .IN1(n7177), .IN2(P2_add_918_n45), 
        .QN(P2_add_918_n269) );
  OR2X1 P2_add_918_U294 ( .IN2(n7177), .IN1(P2_add_918_n45), 
        .Q(P2_add_918_n271) );
  NAND2X0 P2_add_918_U293 ( .IN1(P2_N2608), .IN2(P2_add_918_n271), 
        .QN(P2_add_918_n270) );
  NAND2X0 P2_add_918_U292 ( .IN1(P2_add_918_n269), .IN2(P2_add_918_n270), 
        .QN(P2_add_918_n38) );
  NAND2X0 P2_add_918_U291 ( .IN1(n7173), .IN2(P2_add_918_n38), 
        .QN(P2_add_918_n266) );
  OR2X1 P2_add_918_U290 ( .IN2(n7173), .IN1(P2_add_918_n38), 
        .Q(P2_add_918_n268) );
  NAND2X0 P2_add_918_U289 ( .IN1(P2_N2609), .IN2(P2_add_918_n268), 
        .QN(P2_add_918_n267) );
  NAND2X0 P2_add_918_U288 ( .IN1(P2_add_918_n266), .IN2(P2_add_918_n267), 
        .QN(P2_add_918_n31) );
  NAND2X0 P2_add_918_U287 ( .IN1(n7165), .IN2(P2_add_918_n31), 
        .QN(P2_add_918_n263) );
  OR2X1 P2_add_918_U286 ( .IN2(n7165), .IN1(P2_add_918_n31), 
        .Q(P2_add_918_n265) );
  NAND2X0 P2_add_918_U285 ( .IN1(P2_N2610), .IN2(P2_add_918_n265), 
        .QN(P2_add_918_n264) );
  NAND2X0 P2_add_918_U284 ( .IN1(P2_add_918_n263), .IN2(P2_add_918_n264), 
        .QN(P2_add_918_n24) );
  NAND2X0 P2_add_918_U283 ( .IN1(P2_N5077), .IN2(P2_add_918_n24), 
        .QN(P2_add_918_n260) );
  OR2X1 P2_add_918_U282 ( .IN2(P2_N5077), .IN1(P2_add_918_n24), 
        .Q(P2_add_918_n262) );
  NAND2X0 P2_add_918_U281 ( .IN1(P2_N2611), .IN2(P2_add_918_n262), 
        .QN(P2_add_918_n261) );
  NAND2X0 P2_add_918_U280 ( .IN1(P2_add_918_n260), .IN2(P2_add_918_n261), 
        .QN(P2_add_918_n17) );
  NAND2X0 P2_sub_938_U31 ( .IN1(P2_sub_938_n36), .IN2(P2_sub_938_n37), 
        .QN(P2_N3224) );
  NAND2X0 P2_sub_938_U30 ( .IN1(n7165), .IN2(P2_sub_938_n35), 
        .QN(P2_sub_938_n33) );
  OR2X1 P2_sub_938_U29 ( .IN2(n7165), .IN1(P2_sub_938_n35), .Q(P2_sub_938_n34)
         );
  NAND2X0 P2_sub_938_U28 ( .IN1(P2_sub_938_n33), .IN2(P2_sub_938_n34), 
        .QN(P2_sub_938_n31) );
  NAND2X0 P2_sub_938_U27 ( .IN1(P2_sub_938_n31), .IN2(P2_sub_938_n32), 
        .QN(P2_sub_938_n29) );
  OR2X1 P2_sub_938_U26 ( .IN2(P2_sub_938_n32), .IN1(P2_sub_938_n31), 
        .Q(P2_sub_938_n30) );
  NAND2X0 P2_sub_938_U25 ( .IN1(P2_sub_938_n29), .IN2(P2_sub_938_n30), 
        .QN(P2_N3225) );
  NAND2X0 P2_sub_938_U24 ( .IN1(P2_N5077), .IN2(P2_sub_938_n28), 
        .QN(P2_sub_938_n26) );
  OR2X1 P2_sub_938_U23 ( .IN2(P2_N5077), .IN1(P2_sub_938_n28), 
        .Q(P2_sub_938_n27) );
  NAND2X0 P2_sub_938_U22 ( .IN1(P2_sub_938_n26), .IN2(P2_sub_938_n27), 
        .QN(P2_sub_938_n24) );
  NAND2X0 P2_sub_938_U21 ( .IN1(P2_sub_938_n24), .IN2(P2_sub_938_n25), 
        .QN(P2_sub_938_n22) );
  OR2X1 P2_sub_938_U20 ( .IN2(P2_sub_938_n25), .IN1(P2_sub_938_n24), 
        .Q(P2_sub_938_n23) );
  NAND2X0 P2_sub_938_U19 ( .IN1(P2_sub_938_n22), .IN2(P2_sub_938_n23), 
        .QN(P2_N3226) );
  NAND2X0 P2_sub_938_U18 ( .IN1(P2_N5078), .IN2(P2_sub_938_n21), 
        .QN(P2_sub_938_n19) );
  OR2X1 P2_sub_938_U17 ( .IN2(P2_N5078), .IN1(P2_sub_938_n21), 
        .Q(P2_sub_938_n20) );
  NAND2X0 P2_sub_938_U16 ( .IN1(P2_sub_938_n19), .IN2(P2_sub_938_n20), 
        .QN(P2_sub_938_n17) );
  NAND2X0 P2_sub_938_U15 ( .IN1(P2_sub_938_n17), .IN2(P2_sub_938_n18), 
        .QN(P2_sub_938_n15) );
  OR2X1 P2_sub_938_U14 ( .IN2(P2_sub_938_n18), .IN1(P2_sub_938_n17), 
        .Q(P2_sub_938_n16) );
  NAND2X0 P2_sub_938_U13 ( .IN1(P2_sub_938_n15), .IN2(P2_sub_938_n16), 
        .QN(P2_N3227) );
  NAND2X0 P2_sub_938_U12 ( .IN1(P2_N5079), .IN2(P2_sub_938_n14), 
        .QN(P2_sub_938_n12) );
  OR2X1 P2_sub_938_U11 ( .IN2(P2_N5079), .IN1(P2_sub_938_n14), 
        .Q(P2_sub_938_n13) );
  NAND2X0 P2_sub_938_U10 ( .IN1(P2_sub_938_n12), .IN2(P2_sub_938_n13), 
        .QN(P2_sub_938_n10) );
  NAND2X0 P2_sub_938_U9 ( .IN1(P2_sub_938_n10), .IN2(P2_sub_938_n11), 
        .QN(P2_sub_938_n8) );
  OR2X1 P2_sub_938_U8 ( .IN2(P2_sub_938_n11), .IN1(P2_sub_938_n10), 
        .Q(P2_sub_938_n9) );
  NAND2X0 P2_sub_938_U7 ( .IN1(P2_sub_938_n8), .IN2(P2_sub_938_n9), 
        .QN(P2_N3228) );
  NAND2X0 P2_sub_938_U6 ( .IN1(n7151), .IN2(P2_sub_938_n7), .QN(P2_sub_938_n5)
         );
  OR2X1 P2_sub_938_U5 ( .IN2(n7151), .IN1(P2_sub_938_n7), .Q(P2_sub_938_n6) );
  NAND2X0 P2_sub_938_U4 ( .IN1(P2_sub_938_n5), .IN2(P2_sub_938_n6), 
        .QN(P2_sub_938_n3) );
  NAND2X0 P2_sub_938_U3 ( .IN1(P2_sub_938_n3), .IN2(P2_sub_938_n4), 
        .QN(P2_sub_938_n1) );
  OR2X1 P2_sub_938_U2 ( .IN2(P2_sub_938_n4), .IN1(P2_sub_938_n3), 
        .Q(P2_sub_938_n2) );
  NAND2X0 P2_sub_938_U1 ( .IN1(P2_sub_938_n1), .IN2(P2_sub_938_n2), 
        .QN(P2_N3229) );
  NAND2X0 P2_sub_938_U124 ( .IN1(n7247), .IN2(P2_sub_938_n115), 
        .QN(P2_sub_938_n127) );
  OR2X1 P2_sub_938_U123 ( .IN2(n7247), .IN1(P2_sub_938_n115), 
        .Q(P2_sub_938_n128) );
  NAND2X0 P2_sub_938_U122 ( .IN1(P2_sub_938_n127), .IN2(P2_sub_938_n128), 
        .QN(P2_sub_938_n121) );
  NAND2X0 P2_sub_938_U121 ( .IN1(P2_N5092), .IN2(P2_sub_938_n126), 
        .QN(P2_sub_938_n122) );
  OR2X1 P2_sub_938_U120 ( .IN2(P2_N5092), .IN1(P2_sub_938_n126), 
        .Q(P2_sub_938_n124) );
  NAND2X0 P2_sub_938_U119 ( .IN1(P2_sub_938_n124), .IN2(P2_sub_938_n125), 
        .QN(P2_sub_938_n123) );
  NAND2X0 P2_sub_938_U118 ( .IN1(P2_sub_938_n122), .IN2(P2_sub_938_n123), 
        .QN(P2_sub_938_n116) );
  NAND2X0 P2_sub_938_U117 ( .IN1(P2_sub_938_n121), .IN2(P2_sub_938_n116), 
        .QN(P2_sub_938_n119) );
  OR2X1 P2_sub_938_U116 ( .IN2(P2_sub_938_n116), .IN1(P2_sub_938_n121), 
        .Q(P2_sub_938_n120) );
  NAND2X0 P2_sub_938_U115 ( .IN1(P2_sub_938_n119), .IN2(P2_sub_938_n120), 
        .QN(P2_N3242) );
  INVX0 P2_sub_938_U114 ( .ZN(P2_sub_938_n105), .INP(P2_N3001) );
  NAND2X0 P2_sub_938_U113 ( .IN1(P2_N5094), .IN2(P2_sub_938_n105), 
        .QN(P2_sub_938_n117) );
  OR2X1 P2_sub_938_U112 ( .IN2(P2_N5094), .IN1(P2_sub_938_n105), 
        .Q(P2_sub_938_n118) );
  NAND2X0 P2_sub_938_U111 ( .IN1(P2_sub_938_n117), .IN2(P2_sub_938_n118), 
        .QN(P2_sub_938_n111) );
  NAND2X0 P2_sub_938_U110 ( .IN1(n7247), .IN2(P2_sub_938_n116), 
        .QN(P2_sub_938_n112) );
  OR2X1 P2_sub_938_U109 ( .IN2(n7247), .IN1(P2_sub_938_n116), 
        .Q(P2_sub_938_n114) );
  NAND2X0 P2_sub_938_U108 ( .IN1(P2_sub_938_n114), .IN2(P2_sub_938_n115), 
        .QN(P2_sub_938_n113) );
  NAND2X0 P2_sub_938_U107 ( .IN1(P2_sub_938_n112), .IN2(P2_sub_938_n113), 
        .QN(P2_sub_938_n106) );
  NAND2X0 P2_sub_938_U106 ( .IN1(P2_sub_938_n111), .IN2(P2_sub_938_n106), 
        .QN(P2_sub_938_n109) );
  OR2X1 P2_sub_938_U105 ( .IN2(P2_sub_938_n106), .IN1(P2_sub_938_n111), 
        .Q(P2_sub_938_n110) );
  NAND2X0 P2_sub_938_U104 ( .IN1(P2_sub_938_n109), .IN2(P2_sub_938_n110), 
        .QN(P2_N3243) );
  INVX0 P2_sub_938_U103 ( .ZN(P2_sub_938_n95), .INP(P2_N3002) );
  NAND2X0 P2_sub_938_U102 ( .IN1(P2_N5095), .IN2(P2_sub_938_n95), 
        .QN(P2_sub_938_n107) );
  OR2X1 P2_sub_938_U101 ( .IN2(P2_N5095), .IN1(P2_sub_938_n95), 
        .Q(P2_sub_938_n108) );
  NAND2X0 P2_sub_938_U100 ( .IN1(P2_sub_938_n107), .IN2(P2_sub_938_n108), 
        .QN(P2_sub_938_n101) );
  NAND2X0 P2_sub_938_U99 ( .IN1(P2_N5094), .IN2(P2_sub_938_n106), 
        .QN(P2_sub_938_n102) );
  OR2X1 P2_sub_938_U98 ( .IN2(P2_N5094), .IN1(P2_sub_938_n106), 
        .Q(P2_sub_938_n104) );
  NAND2X0 P2_sub_938_U97 ( .IN1(P2_sub_938_n104), .IN2(P2_sub_938_n105), 
        .QN(P2_sub_938_n103) );
  NAND2X0 P2_sub_938_U96 ( .IN1(P2_sub_938_n102), .IN2(P2_sub_938_n103), 
        .QN(P2_sub_938_n96) );
  NAND2X0 P2_sub_938_U95 ( .IN1(P2_sub_938_n101), .IN2(P2_sub_938_n96), 
        .QN(P2_sub_938_n99) );
  OR2X1 P2_sub_938_U94 ( .IN2(P2_sub_938_n96), .IN1(P2_sub_938_n101), 
        .Q(P2_sub_938_n100) );
  NAND2X0 P2_sub_938_U93 ( .IN1(P2_sub_938_n99), .IN2(P2_sub_938_n100), 
        .QN(P2_N3244) );
  INVX0 P2_sub_938_U92 ( .ZN(P2_sub_938_n85), .INP(P2_N3003) );
  NAND2X0 P2_sub_938_U91 ( .IN1(n7237), .IN2(P2_sub_938_n85), 
        .QN(P2_sub_938_n97) );
  OR2X1 P2_sub_938_U90 ( .IN2(n7237), .IN1(P2_sub_938_n85), .Q(P2_sub_938_n98)
         );
  NAND2X0 P2_sub_938_U89 ( .IN1(P2_sub_938_n97), .IN2(P2_sub_938_n98), 
        .QN(P2_sub_938_n91) );
  NAND2X0 P2_sub_938_U88 ( .IN1(P2_N5095), .IN2(P2_sub_938_n96), 
        .QN(P2_sub_938_n92) );
  OR2X1 P2_sub_938_U87 ( .IN2(P2_N5095), .IN1(P2_sub_938_n96), 
        .Q(P2_sub_938_n94) );
  NAND2X0 P2_sub_938_U86 ( .IN1(P2_sub_938_n94), .IN2(P2_sub_938_n95), 
        .QN(P2_sub_938_n93) );
  NAND2X0 P2_sub_938_U85 ( .IN1(P2_sub_938_n92), .IN2(P2_sub_938_n93), 
        .QN(P2_sub_938_n86) );
  NAND2X0 P2_sub_938_U84 ( .IN1(P2_sub_938_n91), .IN2(P2_sub_938_n86), 
        .QN(P2_sub_938_n89) );
  OR2X1 P2_sub_938_U83 ( .IN2(P2_sub_938_n86), .IN1(P2_sub_938_n91), 
        .Q(P2_sub_938_n90) );
  NAND2X0 P2_sub_938_U82 ( .IN1(P2_sub_938_n89), .IN2(P2_sub_938_n90), 
        .QN(P2_N3245) );
  INVX0 P2_sub_938_U81 ( .ZN(P2_sub_938_n75), .INP(P2_N3004) );
  NAND2X0 P2_sub_938_U80 ( .IN1(n7231), .IN2(P2_sub_938_n75), 
        .QN(P2_sub_938_n87) );
  OR2X1 P2_sub_938_U79 ( .IN2(n7231), .IN1(P2_sub_938_n75), .Q(P2_sub_938_n88)
         );
  NAND2X0 P2_sub_938_U78 ( .IN1(P2_sub_938_n87), .IN2(P2_sub_938_n88), 
        .QN(P2_sub_938_n81) );
  NAND2X0 P2_sub_938_U77 ( .IN1(n7237), .IN2(P2_sub_938_n86), 
        .QN(P2_sub_938_n82) );
  OR2X1 P2_sub_938_U76 ( .IN2(n7237), .IN1(P2_sub_938_n86), .Q(P2_sub_938_n84)
         );
  NAND2X0 P2_sub_938_U75 ( .IN1(P2_sub_938_n84), .IN2(P2_sub_938_n85), 
        .QN(P2_sub_938_n83) );
  NAND2X0 P2_sub_938_U74 ( .IN1(P2_sub_938_n82), .IN2(P2_sub_938_n83), 
        .QN(P2_sub_938_n76) );
  NAND2X0 P2_sub_938_U73 ( .IN1(P2_sub_938_n81), .IN2(P2_sub_938_n76), 
        .QN(P2_sub_938_n79) );
  OR2X1 P2_sub_938_U72 ( .IN2(P2_sub_938_n76), .IN1(P2_sub_938_n81), 
        .Q(P2_sub_938_n80) );
  NAND2X0 P2_sub_938_U71 ( .IN1(P2_sub_938_n79), .IN2(P2_sub_938_n80), 
        .QN(P2_N3246) );
  INVX0 P2_sub_938_U70 ( .ZN(P2_sub_938_n64), .INP(P2_N3005) );
  NAND2X0 P2_sub_938_U69 ( .IN1(P2_N5098), .IN2(P2_sub_938_n64), 
        .QN(P2_sub_938_n77) );
  OR2X1 P2_sub_938_U68 ( .IN2(P2_N5098), .IN1(P2_sub_938_n64), 
        .Q(P2_sub_938_n78) );
  NAND2X0 P2_sub_938_U67 ( .IN1(P2_sub_938_n77), .IN2(P2_sub_938_n78), 
        .QN(P2_sub_938_n71) );
  NAND2X0 P2_sub_938_U66 ( .IN1(n7231), .IN2(P2_sub_938_n76), 
        .QN(P2_sub_938_n72) );
  OR2X1 P2_sub_938_U65 ( .IN2(n7231), .IN1(P2_sub_938_n76), .Q(P2_sub_938_n74)
         );
  NAND2X0 P2_sub_938_U64 ( .IN1(P2_sub_938_n74), .IN2(P2_sub_938_n75), 
        .QN(P2_sub_938_n73) );
  NAND2X0 P2_sub_938_U63 ( .IN1(P2_sub_938_n72), .IN2(P2_sub_938_n73), 
        .QN(P2_sub_938_n65) );
  NAND2X0 P2_sub_938_U62 ( .IN1(P2_sub_938_n71), .IN2(P2_sub_938_n65), 
        .QN(P2_sub_938_n69) );
  OR2X1 P2_sub_938_U61 ( .IN2(P2_sub_938_n65), .IN1(P2_sub_938_n71), 
        .Q(P2_sub_938_n70) );
  NAND2X0 P2_sub_938_U60 ( .IN1(P2_sub_938_n69), .IN2(P2_sub_938_n70), 
        .QN(P2_N3247) );
  OR2X1 P2_sub_938_U58 ( .IN2(P2_N3006), .IN1(n7222), .Q(P2_sub_938_n66) );
  NAND2X0 P2_sub_938_U57 ( .IN1(P2_N3006), .IN2(n7222), .QN(P2_sub_938_n67) );
  NAND2X0 P2_sub_938_U56 ( .IN1(P2_sub_938_n66), .IN2(P2_sub_938_n67), 
        .QN(P2_sub_938_n60) );
  NAND2X0 P2_sub_938_U55 ( .IN1(P2_N5098), .IN2(P2_sub_938_n65), 
        .QN(P2_sub_938_n61) );
  OR2X1 P2_sub_938_U54 ( .IN2(P2_N5098), .IN1(P2_sub_938_n65), 
        .Q(P2_sub_938_n63) );
  NAND2X0 P2_sub_938_U53 ( .IN1(P2_sub_938_n63), .IN2(P2_sub_938_n64), 
        .QN(P2_sub_938_n62) );
  NAND2X0 P2_sub_938_U52 ( .IN1(P2_sub_938_n61), .IN2(P2_sub_938_n62), 
        .QN(P2_sub_938_n59) );
  NAND2X0 P2_sub_938_U51 ( .IN1(P2_sub_938_n60), .IN2(P2_sub_938_n59), 
        .QN(P2_sub_938_n57) );
  OR2X1 P2_sub_938_U50 ( .IN2(P2_sub_938_n60), .IN1(P2_sub_938_n59), 
        .Q(P2_sub_938_n58) );
  NAND2X0 P2_sub_938_U49 ( .IN1(P2_sub_938_n57), .IN2(P2_sub_938_n58), 
        .QN(P2_N3248) );
  NAND2X0 P2_sub_938_U48 ( .IN1(P2_N5073), .IN2(P2_sub_938_n56), 
        .QN(P2_sub_938_n54) );
  OR2X1 P2_sub_938_U47 ( .IN2(P2_N5073), .IN1(P2_sub_938_n56), 
        .Q(P2_sub_938_n55) );
  NAND2X0 P2_sub_938_U46 ( .IN1(P2_sub_938_n54), .IN2(P2_sub_938_n55), 
        .QN(P2_sub_938_n52) );
  NAND2X0 P2_sub_938_U45 ( .IN1(P2_sub_938_n52), .IN2(P2_sub_938_n53), 
        .QN(P2_sub_938_n50) );
  OR2X1 P2_sub_938_U44 ( .IN2(P2_sub_938_n53), .IN1(P2_sub_938_n52), 
        .Q(P2_sub_938_n51) );
  NAND2X0 P2_sub_938_U43 ( .IN1(P2_sub_938_n50), .IN2(P2_sub_938_n51), 
        .QN(P2_N3222) );
  NAND2X0 P2_sub_938_U42 ( .IN1(P2_N5074), .IN2(P2_sub_938_n49), 
        .QN(P2_sub_938_n47) );
  OR2X1 P2_sub_938_U41 ( .IN2(P2_N5074), .IN1(P2_sub_938_n49), 
        .Q(P2_sub_938_n48) );
  NAND2X0 P2_sub_938_U40 ( .IN1(P2_sub_938_n47), .IN2(P2_sub_938_n48), 
        .QN(P2_sub_938_n45) );
  NAND2X0 P2_sub_938_U39 ( .IN1(P2_sub_938_n45), .IN2(P2_sub_938_n46), 
        .QN(P2_sub_938_n43) );
  OR2X1 P2_sub_938_U38 ( .IN2(P2_sub_938_n46), .IN1(P2_sub_938_n45), 
        .Q(P2_sub_938_n44) );
  NAND2X0 P2_sub_938_U37 ( .IN1(P2_sub_938_n43), .IN2(P2_sub_938_n44), 
        .QN(P2_N3223) );
  NAND2X0 P2_sub_938_U36 ( .IN1(P2_N5075), .IN2(P2_sub_938_n42), 
        .QN(P2_sub_938_n40) );
  OR2X1 P2_sub_938_U35 ( .IN2(P2_N5075), .IN1(P2_sub_938_n42), 
        .Q(P2_sub_938_n41) );
  NAND2X0 P2_sub_938_U34 ( .IN1(P2_sub_938_n40), .IN2(P2_sub_938_n41), 
        .QN(P2_sub_938_n38) );
  NAND2X0 P2_sub_938_U33 ( .IN1(P2_sub_938_n38), .IN2(P2_sub_938_n39), 
        .QN(P2_sub_938_n36) );
  OR2X1 P2_sub_938_U32 ( .IN2(P2_sub_938_n39), .IN1(P2_sub_938_n38), 
        .Q(P2_sub_938_n37) );
  OR2X1 P2_sub_938_U217 ( .IN2(P2_N5085), .IN1(P2_sub_938_n203), 
        .Q(P2_sub_938_n216) );
  NAND2X0 P2_sub_938_U216 ( .IN1(P2_sub_938_n215), .IN2(P2_sub_938_n216), 
        .QN(P2_sub_938_n209) );
  NAND2X0 P2_sub_938_U215 ( .IN1(P2_N5084), .IN2(P2_sub_938_n214), 
        .QN(P2_sub_938_n210) );
  OR2X1 P2_sub_938_U214 ( .IN2(P2_N5084), .IN1(P2_sub_938_n214), 
        .Q(P2_sub_938_n212) );
  NAND2X0 P2_sub_938_U213 ( .IN1(P2_sub_938_n212), .IN2(P2_sub_938_n213), 
        .QN(P2_sub_938_n211) );
  NAND2X0 P2_sub_938_U212 ( .IN1(P2_sub_938_n210), .IN2(P2_sub_938_n211), 
        .QN(P2_sub_938_n204) );
  NAND2X0 P2_sub_938_U211 ( .IN1(P2_sub_938_n209), .IN2(P2_sub_938_n204), 
        .QN(P2_sub_938_n207) );
  OR2X1 P2_sub_938_U210 ( .IN2(P2_sub_938_n204), .IN1(P2_sub_938_n209), 
        .Q(P2_sub_938_n208) );
  NAND2X0 P2_sub_938_U209 ( .IN1(P2_sub_938_n207), .IN2(P2_sub_938_n208), 
        .QN(P2_N3234) );
  INVX0 P2_sub_938_U208 ( .ZN(P2_sub_938_n193), .INP(P2_N2993) );
  NAND2X0 P2_sub_938_U207 ( .IN1(P2_N5086), .IN2(P2_sub_938_n193), 
        .QN(P2_sub_938_n205) );
  OR2X1 P2_sub_938_U206 ( .IN2(P2_N5086), .IN1(P2_sub_938_n193), 
        .Q(P2_sub_938_n206) );
  NAND2X0 P2_sub_938_U205 ( .IN1(P2_sub_938_n205), .IN2(P2_sub_938_n206), 
        .QN(P2_sub_938_n199) );
  NAND2X0 P2_sub_938_U204 ( .IN1(P2_N5085), .IN2(P2_sub_938_n204), 
        .QN(P2_sub_938_n200) );
  OR2X1 P2_sub_938_U203 ( .IN2(P2_N5085), .IN1(P2_sub_938_n204), 
        .Q(P2_sub_938_n202) );
  NAND2X0 P2_sub_938_U202 ( .IN1(P2_sub_938_n202), .IN2(P2_sub_938_n203), 
        .QN(P2_sub_938_n201) );
  NAND2X0 P2_sub_938_U201 ( .IN1(P2_sub_938_n200), .IN2(P2_sub_938_n201), 
        .QN(P2_sub_938_n194) );
  NAND2X0 P2_sub_938_U200 ( .IN1(P2_sub_938_n199), .IN2(P2_sub_938_n194), 
        .QN(P2_sub_938_n197) );
  OR2X1 P2_sub_938_U199 ( .IN2(P2_sub_938_n194), .IN1(P2_sub_938_n199), 
        .Q(P2_sub_938_n198) );
  NAND2X0 P2_sub_938_U198 ( .IN1(P2_sub_938_n197), .IN2(P2_sub_938_n198), 
        .QN(P2_N3235) );
  INVX0 P2_sub_938_U197 ( .ZN(P2_sub_938_n183), .INP(P2_N2994) );
  NAND2X0 P2_sub_938_U196 ( .IN1(n7198), .IN2(P2_sub_938_n183), 
        .QN(P2_sub_938_n195) );
  OR2X1 P2_sub_938_U195 ( .IN2(P2_N5087), .IN1(P2_sub_938_n183), 
        .Q(P2_sub_938_n196) );
  NAND2X0 P2_sub_938_U194 ( .IN1(P2_sub_938_n195), .IN2(P2_sub_938_n196), 
        .QN(P2_sub_938_n189) );
  NAND2X0 P2_sub_938_U193 ( .IN1(P2_N5086), .IN2(P2_sub_938_n194), 
        .QN(P2_sub_938_n190) );
  OR2X1 P2_sub_938_U192 ( .IN2(P2_N5086), .IN1(P2_sub_938_n194), 
        .Q(P2_sub_938_n192) );
  NAND2X0 P2_sub_938_U191 ( .IN1(P2_sub_938_n192), .IN2(P2_sub_938_n193), 
        .QN(P2_sub_938_n191) );
  NAND2X0 P2_sub_938_U190 ( .IN1(P2_sub_938_n190), .IN2(P2_sub_938_n191), 
        .QN(P2_sub_938_n184) );
  NAND2X0 P2_sub_938_U189 ( .IN1(P2_sub_938_n189), .IN2(P2_sub_938_n184), 
        .QN(P2_sub_938_n187) );
  OR2X1 P2_sub_938_U188 ( .IN2(P2_sub_938_n184), .IN1(P2_sub_938_n189), 
        .Q(P2_sub_938_n188) );
  NAND2X0 P2_sub_938_U187 ( .IN1(P2_sub_938_n187), .IN2(P2_sub_938_n188), 
        .QN(P2_N3236) );
  INVX0 P2_sub_938_U186 ( .ZN(P2_sub_938_n173), .INP(P2_N2995) );
  NAND2X0 P2_sub_938_U185 ( .IN1(n7194), .IN2(P2_sub_938_n173), 
        .QN(P2_sub_938_n185) );
  OR2X1 P2_sub_938_U184 ( .IN2(n7194), .IN1(P2_sub_938_n173), 
        .Q(P2_sub_938_n186) );
  NAND2X0 P2_sub_938_U183 ( .IN1(P2_sub_938_n185), .IN2(P2_sub_938_n186), 
        .QN(P2_sub_938_n179) );
  NAND2X0 P2_sub_938_U182 ( .IN1(n7198), .IN2(P2_sub_938_n184), 
        .QN(P2_sub_938_n180) );
  OR2X1 P2_sub_938_U181 ( .IN2(n7198), .IN1(P2_sub_938_n184), 
        .Q(P2_sub_938_n182) );
  NAND2X0 P2_sub_938_U180 ( .IN1(P2_sub_938_n182), .IN2(P2_sub_938_n183), 
        .QN(P2_sub_938_n181) );
  NAND2X0 P2_sub_938_U179 ( .IN1(P2_sub_938_n180), .IN2(P2_sub_938_n181), 
        .QN(P2_sub_938_n174) );
  NAND2X0 P2_sub_938_U178 ( .IN1(P2_sub_938_n179), .IN2(P2_sub_938_n174), 
        .QN(P2_sub_938_n177) );
  OR2X1 P2_sub_938_U177 ( .IN2(P2_sub_938_n174), .IN1(P2_sub_938_n179), 
        .Q(P2_sub_938_n178) );
  NAND2X0 P2_sub_938_U176 ( .IN1(P2_sub_938_n177), .IN2(P2_sub_938_n178), 
        .QN(P2_N3237) );
  INVX0 P2_sub_938_U175 ( .ZN(P2_sub_938_n163), .INP(P2_N2996) );
  NAND2X0 P2_sub_938_U174 ( .IN1(n7187), .IN2(P2_sub_938_n163), 
        .QN(P2_sub_938_n175) );
  OR2X1 P2_sub_938_U173 ( .IN2(n7187), .IN1(P2_sub_938_n163), 
        .Q(P2_sub_938_n176) );
  NAND2X0 P2_sub_938_U172 ( .IN1(P2_sub_938_n175), .IN2(P2_sub_938_n176), 
        .QN(P2_sub_938_n169) );
  NAND2X0 P2_sub_938_U171 ( .IN1(n7194), .IN2(P2_sub_938_n174), 
        .QN(P2_sub_938_n170) );
  OR2X1 P2_sub_938_U170 ( .IN2(n7194), .IN1(P2_sub_938_n174), 
        .Q(P2_sub_938_n172) );
  NAND2X0 P2_sub_938_U169 ( .IN1(P2_sub_938_n172), .IN2(P2_sub_938_n173), 
        .QN(P2_sub_938_n171) );
  NAND2X0 P2_sub_938_U168 ( .IN1(P2_sub_938_n170), .IN2(P2_sub_938_n171), 
        .QN(P2_sub_938_n164) );
  NAND2X0 P2_sub_938_U167 ( .IN1(P2_sub_938_n169), .IN2(P2_sub_938_n164), 
        .QN(P2_sub_938_n167) );
  OR2X1 P2_sub_938_U166 ( .IN2(P2_sub_938_n164), .IN1(P2_sub_938_n169), 
        .Q(P2_sub_938_n168) );
  NAND2X0 P2_sub_938_U165 ( .IN1(P2_sub_938_n167), .IN2(P2_sub_938_n168), 
        .QN(P2_N3238) );
  INVX0 P2_sub_938_U164 ( .ZN(P2_sub_938_n145), .INP(P2_N2997) );
  NAND2X0 P2_sub_938_U163 ( .IN1(P2_N5090), .IN2(P2_sub_938_n145), 
        .QN(P2_sub_938_n165) );
  OR2X1 P2_sub_938_U162 ( .IN2(P2_N5090), .IN1(P2_sub_938_n145), 
        .Q(P2_sub_938_n166) );
  NAND2X0 P2_sub_938_U161 ( .IN1(P2_sub_938_n165), .IN2(P2_sub_938_n166), 
        .QN(P2_sub_938_n159) );
  NAND2X0 P2_sub_938_U160 ( .IN1(n7187), .IN2(P2_sub_938_n164), 
        .QN(P2_sub_938_n160) );
  OR2X1 P2_sub_938_U159 ( .IN2(n7187), .IN1(P2_sub_938_n164), 
        .Q(P2_sub_938_n162) );
  NAND2X0 P2_sub_938_U158 ( .IN1(P2_sub_938_n162), .IN2(P2_sub_938_n163), 
        .QN(P2_sub_938_n161) );
  NAND2X0 P2_sub_938_U157 ( .IN1(P2_sub_938_n160), .IN2(P2_sub_938_n161), 
        .QN(P2_sub_938_n146) );
  NAND2X0 P2_sub_938_U156 ( .IN1(P2_sub_938_n159), .IN2(P2_sub_938_n146), 
        .QN(P2_sub_938_n157) );
  OR2X1 P2_sub_938_U155 ( .IN2(P2_sub_938_n146), .IN1(P2_sub_938_n159), 
        .Q(P2_sub_938_n158) );
  NAND2X0 P2_sub_938_U154 ( .IN1(P2_sub_938_n157), .IN2(P2_sub_938_n158), 
        .QN(P2_N3239) );
  NAND2X0 P2_sub_938_U153 ( .IN1(P2_N5072), .IN2(P2_sub_938_n156), 
        .QN(P2_sub_938_n153) );
  NAND2X0 P2_sub_938_U152 ( .IN1(P2_N2979), .IN2(n7184), .QN(P2_sub_938_n154)
         );
  NAND2X0 P2_sub_938_U151 ( .IN1(P2_sub_938_n153), .IN2(P2_sub_938_n154), 
        .QN(P2_sub_938_n151) );
  NAND2X0 P2_sub_938_U150 ( .IN1(P2_sub_938_n151), .IN2(P2_sub_938_n152), 
        .QN(P2_sub_938_n149) );
  OR2X1 P2_sub_938_U149 ( .IN2(P2_sub_938_n152), .IN1(P2_sub_938_n151), 
        .Q(P2_sub_938_n150) );
  NAND2X0 P2_sub_938_U148 ( .IN1(P2_sub_938_n149), .IN2(P2_sub_938_n150), 
        .QN(P2_N3221) );
  INVX0 P2_sub_938_U147 ( .ZN(P2_sub_938_n135), .INP(P2_N2998) );
  NAND2X0 P2_sub_938_U146 ( .IN1(P2_N5091), .IN2(P2_sub_938_n135), 
        .QN(P2_sub_938_n147) );
  OR2X1 P2_sub_938_U145 ( .IN2(P2_N5091), .IN1(P2_sub_938_n135), 
        .Q(P2_sub_938_n148) );
  NAND2X0 P2_sub_938_U144 ( .IN1(P2_sub_938_n147), .IN2(P2_sub_938_n148), 
        .QN(P2_sub_938_n141) );
  NAND2X0 P2_sub_938_U143 ( .IN1(P2_N5090), .IN2(P2_sub_938_n146), 
        .QN(P2_sub_938_n142) );
  OR2X1 P2_sub_938_U142 ( .IN2(P2_N5090), .IN1(P2_sub_938_n146), 
        .Q(P2_sub_938_n144) );
  NAND2X0 P2_sub_938_U141 ( .IN1(P2_sub_938_n144), .IN2(P2_sub_938_n145), 
        .QN(P2_sub_938_n143) );
  NAND2X0 P2_sub_938_U140 ( .IN1(P2_sub_938_n142), .IN2(P2_sub_938_n143), 
        .QN(P2_sub_938_n136) );
  NAND2X0 P2_sub_938_U139 ( .IN1(P2_sub_938_n141), .IN2(P2_sub_938_n136), 
        .QN(P2_sub_938_n139) );
  OR2X1 P2_sub_938_U138 ( .IN2(P2_sub_938_n136), .IN1(P2_sub_938_n141), 
        .Q(P2_sub_938_n140) );
  NAND2X0 P2_sub_938_U137 ( .IN1(P2_sub_938_n139), .IN2(P2_sub_938_n140), 
        .QN(P2_N3240) );
  INVX0 P2_sub_938_U136 ( .ZN(P2_sub_938_n125), .INP(P2_N2999) );
  NAND2X0 P2_sub_938_U135 ( .IN1(P2_N5092), .IN2(P2_sub_938_n125), 
        .QN(P2_sub_938_n137) );
  OR2X1 P2_sub_938_U134 ( .IN2(P2_N5092), .IN1(P2_sub_938_n125), 
        .Q(P2_sub_938_n138) );
  NAND2X0 P2_sub_938_U133 ( .IN1(P2_sub_938_n137), .IN2(P2_sub_938_n138), 
        .QN(P2_sub_938_n131) );
  NAND2X0 P2_sub_938_U132 ( .IN1(P2_N5091), .IN2(P2_sub_938_n136), 
        .QN(P2_sub_938_n132) );
  OR2X1 P2_sub_938_U131 ( .IN2(P2_N5091), .IN1(P2_sub_938_n136), 
        .Q(P2_sub_938_n134) );
  NAND2X0 P2_sub_938_U130 ( .IN1(P2_sub_938_n134), .IN2(P2_sub_938_n135), 
        .QN(P2_sub_938_n133) );
  NAND2X0 P2_sub_938_U129 ( .IN1(P2_sub_938_n132), .IN2(P2_sub_938_n133), 
        .QN(P2_sub_938_n126) );
  NAND2X0 P2_sub_938_U128 ( .IN1(P2_sub_938_n131), .IN2(P2_sub_938_n126), 
        .QN(P2_sub_938_n129) );
  OR2X1 P2_sub_938_U127 ( .IN2(P2_sub_938_n126), .IN1(P2_sub_938_n131), 
        .Q(P2_sub_938_n130) );
  NAND2X0 P2_sub_938_U126 ( .IN1(P2_sub_938_n129), .IN2(P2_sub_938_n130), 
        .QN(P2_N3241) );
  INVX0 P2_sub_938_U125 ( .ZN(P2_sub_938_n115), .INP(P2_N3000) );
  INVX0 P2_sub_938_U310 ( .ZN(P2_sub_938_n281), .INP(P2_N2978) );
  NOR2X0 P2_sub_938_U309 ( .QN(P2_sub_938_n277), .IN1(P2_sub_938_n281), 
        .IN2(n7035) );
  INVX0 P2_sub_938_U308 ( .ZN(P2_sub_938_n152), .INP(P2_sub_938_n277) );
  NAND2X0 P2_sub_938_U307 ( .IN1(n7035), .IN2(P2_sub_938_n281), 
        .QN(P2_sub_938_n280) );
  NAND2X0 P2_sub_938_U306 ( .IN1(P2_sub_938_n152), .IN2(P2_sub_938_n280), 
        .QN(P2_N3220) );
  INVX0 P2_sub_938_U305 ( .ZN(P2_sub_938_n243), .INP(P2_N2988) );
  NAND2X0 P2_sub_938_U304 ( .IN1(P2_N5081), .IN2(P2_sub_938_n243), 
        .QN(P2_sub_938_n278) );
  OR2X1 P2_sub_938_U303 ( .IN2(P2_N5081), .IN1(P2_sub_938_n243), 
        .Q(P2_sub_938_n279) );
  NAND2X0 P2_sub_938_U302 ( .IN1(P2_sub_938_n278), .IN2(P2_sub_938_n279), 
        .QN(P2_sub_938_n249) );
  NAND2X0 P2_sub_938_U301 ( .IN1(P2_N5072), .IN2(P2_sub_938_n152), 
        .QN(P2_sub_938_n274) );
  NAND2X0 P2_sub_938_U299 ( .IN1(P2_sub_938_n277), .IN2(n7184), 
        .QN(P2_sub_938_n276) );
  INVX0 P2_sub_938_U298 ( .ZN(P2_sub_938_n156), .INP(P2_N2979) );
  NAND2X0 P2_sub_938_U297 ( .IN1(P2_sub_938_n276), .IN2(P2_sub_938_n156), 
        .QN(P2_sub_938_n275) );
  NAND2X0 P2_sub_938_U296 ( .IN1(P2_sub_938_n274), .IN2(P2_sub_938_n275), 
        .QN(P2_sub_938_n53) );
  NAND2X0 P2_sub_938_U295 ( .IN1(P2_N5073), .IN2(P2_sub_938_n53), 
        .QN(P2_sub_938_n271) );
  OR2X1 P2_sub_938_U294 ( .IN2(P2_N5073), .IN1(P2_sub_938_n53), 
        .Q(P2_sub_938_n273) );
  INVX0 P2_sub_938_U293 ( .ZN(P2_sub_938_n56), .INP(P2_N2980) );
  NAND2X0 P2_sub_938_U292 ( .IN1(P2_sub_938_n273), .IN2(P2_sub_938_n56), 
        .QN(P2_sub_938_n272) );
  NAND2X0 P2_sub_938_U291 ( .IN1(P2_sub_938_n271), .IN2(P2_sub_938_n272), 
        .QN(P2_sub_938_n46) );
  NAND2X0 P2_sub_938_U290 ( .IN1(P2_N5074), .IN2(P2_sub_938_n46), 
        .QN(P2_sub_938_n268) );
  OR2X1 P2_sub_938_U289 ( .IN2(P2_N5074), .IN1(P2_sub_938_n46), 
        .Q(P2_sub_938_n270) );
  INVX0 P2_sub_938_U288 ( .ZN(P2_sub_938_n49), .INP(P2_N2981) );
  NAND2X0 P2_sub_938_U287 ( .IN1(P2_sub_938_n270), .IN2(P2_sub_938_n49), 
        .QN(P2_sub_938_n269) );
  NAND2X0 P2_sub_938_U286 ( .IN1(P2_sub_938_n268), .IN2(P2_sub_938_n269), 
        .QN(P2_sub_938_n39) );
  NAND2X0 P2_sub_938_U285 ( .IN1(P2_N5075), .IN2(P2_sub_938_n39), 
        .QN(P2_sub_938_n265) );
  OR2X1 P2_sub_938_U284 ( .IN2(P2_N5075), .IN1(P2_sub_938_n39), 
        .Q(P2_sub_938_n267) );
  INVX0 P2_sub_938_U283 ( .ZN(P2_sub_938_n42), .INP(P2_N2982) );
  NAND2X0 P2_sub_938_U282 ( .IN1(P2_sub_938_n267), .IN2(P2_sub_938_n42), 
        .QN(P2_sub_938_n266) );
  NAND2X0 P2_sub_938_U281 ( .IN1(P2_sub_938_n265), .IN2(P2_sub_938_n266), 
        .QN(P2_sub_938_n32) );
  NAND2X0 P2_sub_938_U280 ( .IN1(n7165), .IN2(P2_sub_938_n32), 
        .QN(P2_sub_938_n262) );
  OR2X1 P2_sub_938_U279 ( .IN2(n7165), .IN1(P2_sub_938_n32), 
        .Q(P2_sub_938_n264) );
  INVX0 P2_sub_938_U278 ( .ZN(P2_sub_938_n35), .INP(P2_N2983) );
  NAND2X0 P2_sub_938_U277 ( .IN1(P2_sub_938_n264), .IN2(P2_sub_938_n35), 
        .QN(P2_sub_938_n263) );
  NAND2X0 P2_sub_938_U276 ( .IN1(P2_sub_938_n262), .IN2(P2_sub_938_n263), 
        .QN(P2_sub_938_n25) );
  NAND2X0 P2_sub_938_U275 ( .IN1(P2_N5077), .IN2(P2_sub_938_n25), 
        .QN(P2_sub_938_n259) );
  OR2X1 P2_sub_938_U274 ( .IN2(P2_N5077), .IN1(P2_sub_938_n25), 
        .Q(P2_sub_938_n261) );
  INVX0 P2_sub_938_U273 ( .ZN(P2_sub_938_n28), .INP(P2_N2984) );
  NAND2X0 P2_sub_938_U272 ( .IN1(P2_sub_938_n261), .IN2(P2_sub_938_n28), 
        .QN(P2_sub_938_n260) );
  NAND2X0 P2_sub_938_U271 ( .IN1(P2_sub_938_n259), .IN2(P2_sub_938_n260), 
        .QN(P2_sub_938_n18) );
  NAND2X0 P2_sub_938_U270 ( .IN1(P2_N5078), .IN2(P2_sub_938_n18), 
        .QN(P2_sub_938_n256) );
  OR2X1 P2_sub_938_U269 ( .IN2(P2_N5078), .IN1(P2_sub_938_n18), 
        .Q(P2_sub_938_n258) );
  INVX0 P2_sub_938_U268 ( .ZN(P2_sub_938_n21), .INP(P2_N2985) );
  NAND2X0 P2_sub_938_U267 ( .IN1(P2_sub_938_n258), .IN2(P2_sub_938_n21), 
        .QN(P2_sub_938_n257) );
  NAND2X0 P2_sub_938_U266 ( .IN1(P2_sub_938_n256), .IN2(P2_sub_938_n257), 
        .QN(P2_sub_938_n11) );
  NAND2X0 P2_sub_938_U265 ( .IN1(P2_N5079), .IN2(P2_sub_938_n11), 
        .QN(P2_sub_938_n253) );
  OR2X1 P2_sub_938_U264 ( .IN2(P2_N5079), .IN1(P2_sub_938_n11), 
        .Q(P2_sub_938_n255) );
  INVX0 P2_sub_938_U263 ( .ZN(P2_sub_938_n14), .INP(P2_N2986) );
  NAND2X0 P2_sub_938_U262 ( .IN1(P2_sub_938_n255), .IN2(P2_sub_938_n14), 
        .QN(P2_sub_938_n254) );
  NAND2X0 P2_sub_938_U261 ( .IN1(P2_sub_938_n253), .IN2(P2_sub_938_n254), 
        .QN(P2_sub_938_n4) );
  NAND2X0 P2_sub_938_U260 ( .IN1(n7151), .IN2(P2_sub_938_n4), 
        .QN(P2_sub_938_n250) );
  OR2X1 P2_sub_938_U259 ( .IN2(n7151), .IN1(P2_sub_938_n4), 
        .Q(P2_sub_938_n252) );
  INVX0 P2_sub_938_U258 ( .ZN(P2_sub_938_n7), .INP(P2_N2987) );
  NAND2X0 P2_sub_938_U257 ( .IN1(P2_sub_938_n252), .IN2(P2_sub_938_n7), 
        .QN(P2_sub_938_n251) );
  NAND2X0 P2_sub_938_U256 ( .IN1(P2_sub_938_n250), .IN2(P2_sub_938_n251), 
        .QN(P2_sub_938_n244) );
  NAND2X0 P2_sub_938_U255 ( .IN1(P2_sub_938_n249), .IN2(P2_sub_938_n244), 
        .QN(P2_sub_938_n247) );
  OR2X1 P2_sub_938_U254 ( .IN2(P2_sub_938_n244), .IN1(P2_sub_938_n249), 
        .Q(P2_sub_938_n248) );
  NAND2X0 P2_sub_938_U253 ( .IN1(P2_sub_938_n247), .IN2(P2_sub_938_n248), 
        .QN(P2_N3230) );
  INVX0 P2_sub_938_U252 ( .ZN(P2_sub_938_n233), .INP(P2_N2989) );
  NAND2X0 P2_sub_938_U251 ( .IN1(P2_N5082), .IN2(P2_sub_938_n233), 
        .QN(P2_sub_938_n245) );
  OR2X1 P2_sub_938_U250 ( .IN2(P2_N5082), .IN1(P2_sub_938_n233), 
        .Q(P2_sub_938_n246) );
  NAND2X0 P2_sub_938_U249 ( .IN1(P2_sub_938_n245), .IN2(P2_sub_938_n246), 
        .QN(P2_sub_938_n239) );
  NAND2X0 P2_sub_938_U248 ( .IN1(P2_N5081), .IN2(P2_sub_938_n244), 
        .QN(P2_sub_938_n240) );
  OR2X1 P2_sub_938_U247 ( .IN2(P2_N5081), .IN1(P2_sub_938_n244), 
        .Q(P2_sub_938_n242) );
  NAND2X0 P2_sub_938_U246 ( .IN1(P2_sub_938_n242), .IN2(P2_sub_938_n243), 
        .QN(P2_sub_938_n241) );
  NAND2X0 P2_sub_938_U245 ( .IN1(P2_sub_938_n240), .IN2(P2_sub_938_n241), 
        .QN(P2_sub_938_n234) );
  NAND2X0 P2_sub_938_U244 ( .IN1(P2_sub_938_n239), .IN2(P2_sub_938_n234), 
        .QN(P2_sub_938_n237) );
  OR2X1 P2_sub_938_U243 ( .IN2(P2_sub_938_n234), .IN1(P2_sub_938_n239), 
        .Q(P2_sub_938_n238) );
  NAND2X0 P2_sub_938_U242 ( .IN1(P2_sub_938_n237), .IN2(P2_sub_938_n238), 
        .QN(P2_N3231) );
  INVX0 P2_sub_938_U241 ( .ZN(P2_sub_938_n223), .INP(P2_N2990) );
  NAND2X0 P2_sub_938_U240 ( .IN1(P2_N5083), .IN2(P2_sub_938_n223), 
        .QN(P2_sub_938_n235) );
  OR2X1 P2_sub_938_U239 ( .IN2(P2_N5083), .IN1(P2_sub_938_n223), 
        .Q(P2_sub_938_n236) );
  NAND2X0 P2_sub_938_U238 ( .IN1(P2_sub_938_n235), .IN2(P2_sub_938_n236), 
        .QN(P2_sub_938_n229) );
  NAND2X0 P2_sub_938_U237 ( .IN1(P2_N5082), .IN2(P2_sub_938_n234), 
        .QN(P2_sub_938_n230) );
  OR2X1 P2_sub_938_U236 ( .IN2(P2_N5082), .IN1(P2_sub_938_n234), 
        .Q(P2_sub_938_n232) );
  NAND2X0 P2_sub_938_U235 ( .IN1(P2_sub_938_n232), .IN2(P2_sub_938_n233), 
        .QN(P2_sub_938_n231) );
  NAND2X0 P2_sub_938_U234 ( .IN1(P2_sub_938_n230), .IN2(P2_sub_938_n231), 
        .QN(P2_sub_938_n224) );
  NAND2X0 P2_sub_938_U233 ( .IN1(P2_sub_938_n229), .IN2(P2_sub_938_n224), 
        .QN(P2_sub_938_n227) );
  OR2X1 P2_sub_938_U232 ( .IN2(P2_sub_938_n224), .IN1(P2_sub_938_n229), 
        .Q(P2_sub_938_n228) );
  NAND2X0 P2_sub_938_U231 ( .IN1(P2_sub_938_n227), .IN2(P2_sub_938_n228), 
        .QN(P2_N3232) );
  INVX0 P2_sub_938_U230 ( .ZN(P2_sub_938_n213), .INP(P2_N2991) );
  NAND2X0 P2_sub_938_U229 ( .IN1(P2_N5084), .IN2(P2_sub_938_n213), 
        .QN(P2_sub_938_n225) );
  OR2X1 P2_sub_938_U228 ( .IN2(P2_N5084), .IN1(P2_sub_938_n213), 
        .Q(P2_sub_938_n226) );
  NAND2X0 P2_sub_938_U227 ( .IN1(P2_sub_938_n225), .IN2(P2_sub_938_n226), 
        .QN(P2_sub_938_n219) );
  NAND2X0 P2_sub_938_U226 ( .IN1(P2_N5083), .IN2(P2_sub_938_n224), 
        .QN(P2_sub_938_n220) );
  OR2X1 P2_sub_938_U225 ( .IN2(P2_N5083), .IN1(P2_sub_938_n224), 
        .Q(P2_sub_938_n222) );
  NAND2X0 P2_sub_938_U224 ( .IN1(P2_sub_938_n222), .IN2(P2_sub_938_n223), 
        .QN(P2_sub_938_n221) );
  NAND2X0 P2_sub_938_U223 ( .IN1(P2_sub_938_n220), .IN2(P2_sub_938_n221), 
        .QN(P2_sub_938_n214) );
  NAND2X0 P2_sub_938_U222 ( .IN1(P2_sub_938_n219), .IN2(P2_sub_938_n214), 
        .QN(P2_sub_938_n217) );
  OR2X1 P2_sub_938_U221 ( .IN2(P2_sub_938_n214), .IN1(P2_sub_938_n219), 
        .Q(P2_sub_938_n218) );
  NAND2X0 P2_sub_938_U220 ( .IN1(P2_sub_938_n217), .IN2(P2_sub_938_n218), 
        .QN(P2_N3233) );
  INVX0 P2_sub_938_U219 ( .ZN(P2_sub_938_n203), .INP(P2_N2992) );
  NAND2X0 P2_sub_938_U218 ( .IN1(P2_N5085), .IN2(P2_sub_938_n203), 
        .QN(P2_sub_938_n215) );
  NAND2X0 P2_add_958_U61 ( .IN1(P2_N3378), .IN2(P2_add_958_n63), 
        .QN(P2_add_958_n62) );
  NAND2X0 P2_add_958_U60 ( .IN1(P2_add_958_n61), .IN2(P2_add_958_n62), 
        .QN(P2_add_958_n59) );
  NOR2X0 P2_add_958_U59 ( .QN(P2_add_958_n57), .IN1(P2_add_958_n60), 
        .IN2(P2_add_958_n59) );
  AND2X1 P2_add_958_U58 ( .IN1(P2_add_958_n59), .IN2(P2_add_958_n60), 
        .Q(P2_add_958_n58) );
  NOR2X0 P2_add_958_U57 ( .QN(P2_N3621), .IN1(P2_add_958_n57), 
        .IN2(P2_add_958_n58) );
  OR2X1 P2_add_958_U55 ( .IN2(P2_N3353), .IN1(n7182), .Q(P2_add_958_n54) );
  NAND2X0 P2_add_958_U54 ( .IN1(P2_N3353), .IN2(n7182), .QN(P2_add_958_n55) );
  NAND2X0 P2_add_958_U53 ( .IN1(P2_add_958_n54), .IN2(P2_add_958_n55), 
        .QN(P2_add_958_n53) );
  NOR2X0 P2_add_958_U52 ( .QN(P2_add_958_n50), .IN1(P2_add_958_n52), 
        .IN2(P2_add_958_n53) );
  AND2X1 P2_add_958_U51 ( .IN1(P2_add_958_n52), .IN2(P2_add_958_n53), 
        .Q(P2_add_958_n51) );
  NOR2X0 P2_add_958_U50 ( .QN(P2_N3595), .IN1(P2_add_958_n50), 
        .IN2(P2_add_958_n51) );
  OR2X1 P2_add_958_U48 ( .IN2(P2_N3354), .IN1(n7178), .Q(P2_add_958_n47) );
  NAND2X0 P2_add_958_U47 ( .IN1(P2_N3354), .IN2(n7178), .QN(P2_add_958_n48) );
  NAND2X0 P2_add_958_U46 ( .IN1(P2_add_958_n47), .IN2(P2_add_958_n48), 
        .QN(P2_add_958_n46) );
  NOR2X0 P2_add_958_U45 ( .QN(P2_add_958_n43), .IN1(P2_add_958_n45), 
        .IN2(P2_add_958_n46) );
  AND2X1 P2_add_958_U44 ( .IN1(P2_add_958_n45), .IN2(P2_add_958_n46), 
        .Q(P2_add_958_n44) );
  NOR2X0 P2_add_958_U43 ( .QN(P2_N3596), .IN1(P2_add_958_n43), 
        .IN2(P2_add_958_n44) );
  OR2X1 P2_add_958_U41 ( .IN2(P2_N3355), .IN1(n7174), .Q(P2_add_958_n40) );
  NAND2X0 P2_add_958_U40 ( .IN1(P2_N3355), .IN2(n7174), .QN(P2_add_958_n41) );
  NAND2X0 P2_add_958_U39 ( .IN1(P2_add_958_n40), .IN2(P2_add_958_n41), 
        .QN(P2_add_958_n39) );
  NOR2X0 P2_add_958_U38 ( .QN(P2_add_958_n36), .IN1(P2_add_958_n38), 
        .IN2(P2_add_958_n39) );
  AND2X1 P2_add_958_U37 ( .IN1(P2_add_958_n38), .IN2(P2_add_958_n39), 
        .Q(P2_add_958_n37) );
  NOR2X0 P2_add_958_U36 ( .QN(P2_N3597), .IN1(P2_add_958_n36), 
        .IN2(P2_add_958_n37) );
  OR2X1 P2_add_958_U34 ( .IN2(P2_N3356), .IN1(n7166), .Q(P2_add_958_n33) );
  NAND2X0 P2_add_958_U33 ( .IN1(P2_N3356), .IN2(n7166), .QN(P2_add_958_n34) );
  NAND2X0 P2_add_958_U32 ( .IN1(P2_add_958_n33), .IN2(P2_add_958_n34), 
        .QN(P2_add_958_n32) );
  NOR2X0 P2_add_958_U31 ( .QN(P2_add_958_n29), .IN1(P2_add_958_n31), 
        .IN2(P2_add_958_n32) );
  AND2X1 P2_add_958_U30 ( .IN1(P2_add_958_n31), .IN2(P2_add_958_n32), 
        .Q(P2_add_958_n30) );
  NOR2X0 P2_add_958_U29 ( .QN(P2_N3598), .IN1(P2_add_958_n29), 
        .IN2(P2_add_958_n30) );
  OR2X1 P2_add_958_U27 ( .IN2(P2_N3357), .IN1(n7164), .Q(P2_add_958_n26) );
  NAND2X0 P2_add_958_U26 ( .IN1(P2_N3357), .IN2(n7164), .QN(P2_add_958_n27) );
  NAND2X0 P2_add_958_U25 ( .IN1(P2_add_958_n26), .IN2(P2_add_958_n27), 
        .QN(P2_add_958_n25) );
  NOR2X0 P2_add_958_U24 ( .QN(P2_add_958_n22), .IN1(P2_add_958_n24), 
        .IN2(P2_add_958_n25) );
  AND2X1 P2_add_958_U23 ( .IN1(P2_add_958_n24), .IN2(P2_add_958_n25), 
        .Q(P2_add_958_n23) );
  NOR2X0 P2_add_958_U22 ( .QN(P2_N3599), .IN1(P2_add_958_n22), 
        .IN2(P2_add_958_n23) );
  OR2X1 P2_add_958_U20 ( .IN2(P2_N3358), .IN1(n7157), .Q(P2_add_958_n19) );
  NAND2X0 P2_add_958_U19 ( .IN1(P2_N3358), .IN2(n7157), .QN(P2_add_958_n20) );
  NAND2X0 P2_add_958_U18 ( .IN1(P2_add_958_n19), .IN2(P2_add_958_n20), 
        .QN(P2_add_958_n18) );
  NOR2X0 P2_add_958_U17 ( .QN(P2_add_958_n15), .IN1(P2_add_958_n17), 
        .IN2(P2_add_958_n18) );
  AND2X1 P2_add_958_U16 ( .IN1(P2_add_958_n17), .IN2(P2_add_958_n18), 
        .Q(P2_add_958_n16) );
  NOR2X0 P2_add_958_U15 ( .QN(P2_N3600), .IN1(P2_add_958_n15), 
        .IN2(P2_add_958_n16) );
  OR2X1 P2_add_958_U13 ( .IN2(P2_N3359), .IN1(n7153), .Q(P2_add_958_n12) );
  NAND2X0 P2_add_958_U12 ( .IN1(P2_N3359), .IN2(n7153), .QN(P2_add_958_n13) );
  NAND2X0 P2_add_958_U11 ( .IN1(P2_add_958_n12), .IN2(P2_add_958_n13), 
        .QN(P2_add_958_n11) );
  NOR2X0 P2_add_958_U10 ( .QN(P2_add_958_n8), .IN1(P2_add_958_n10), 
        .IN2(P2_add_958_n11) );
  AND2X1 P2_add_958_U9 ( .IN1(P2_add_958_n10), .IN2(P2_add_958_n11), 
        .Q(P2_add_958_n9) );
  NOR2X0 P2_add_958_U8 ( .QN(P2_N3601), .IN1(P2_add_958_n8), 
        .IN2(P2_add_958_n9) );
  OR2X1 P2_add_958_U6 ( .IN2(P2_N3360), .IN1(n7149), .Q(P2_add_958_n5) );
  NAND2X0 P2_add_958_U5 ( .IN1(P2_N3360), .IN2(n7149), .QN(P2_add_958_n6) );
  NAND2X0 P2_add_958_U4 ( .IN1(P2_add_958_n5), .IN2(P2_add_958_n6), 
        .QN(P2_add_958_n4) );
  NOR2X0 P2_add_958_U3 ( .QN(P2_add_958_n1), .IN1(P2_add_958_n3), 
        .IN2(P2_add_958_n4) );
  AND2X1 P2_add_958_U2 ( .IN1(P2_add_958_n3), .IN2(P2_add_958_n4), 
        .Q(P2_add_958_n2) );
  NOR2X0 P2_add_958_U1 ( .QN(P2_N3602), .IN1(P2_add_958_n1), 
        .IN2(P2_add_958_n2) );
  OR2X1 P2_add_958_U154 ( .IN2(P2_N5090), .IN1(P2_add_958_n147), 
        .Q(P2_add_958_n146) );
  NAND2X0 P2_add_958_U153 ( .IN1(P2_N3370), .IN2(P2_add_958_n146), 
        .QN(P2_add_958_n145) );
  NAND2X0 P2_add_958_U152 ( .IN1(P2_add_958_n144), .IN2(P2_add_958_n145), 
        .QN(P2_add_958_n137) );
  OR2X1 P2_add_958_U150 ( .IN2(P2_N3371), .IN1(n7260), .Q(P2_add_958_n141) );
  NAND2X0 P2_add_958_U149 ( .IN1(P2_N3371), .IN2(n7260), .QN(P2_add_958_n142)
         );
  NAND2X0 P2_add_958_U148 ( .IN1(P2_add_958_n141), .IN2(P2_add_958_n142), 
        .QN(P2_add_958_n140) );
  NOR2X0 P2_add_958_U147 ( .QN(P2_add_958_n138), .IN1(P2_add_958_n137), 
        .IN2(P2_add_958_n140) );
  AND2X1 P2_add_958_U146 ( .IN1(P2_add_958_n137), .IN2(P2_add_958_n140), 
        .Q(P2_add_958_n139) );
  NOR2X0 P2_add_958_U145 ( .QN(P2_N3613), .IN1(P2_add_958_n138), 
        .IN2(P2_add_958_n139) );
  NAND2X0 P2_add_958_U144 ( .IN1(P2_N5091), .IN2(P2_add_958_n137), 
        .QN(P2_add_958_n134) );
  OR2X1 P2_add_958_U143 ( .IN2(P2_N5091), .IN1(P2_add_958_n137), 
        .Q(P2_add_958_n136) );
  NAND2X0 P2_add_958_U142 ( .IN1(P2_N3371), .IN2(P2_add_958_n136), 
        .QN(P2_add_958_n135) );
  NAND2X0 P2_add_958_U141 ( .IN1(P2_add_958_n134), .IN2(P2_add_958_n135), 
        .QN(P2_add_958_n127) );
  OR2X1 P2_add_958_U139 ( .IN2(P2_N3372), .IN1(n7253), .Q(P2_add_958_n131) );
  NAND2X0 P2_add_958_U138 ( .IN1(P2_N3372), .IN2(n7253), .QN(P2_add_958_n132)
         );
  NAND2X0 P2_add_958_U137 ( .IN1(P2_add_958_n131), .IN2(P2_add_958_n132), 
        .QN(P2_add_958_n130) );
  NOR2X0 P2_add_958_U136 ( .QN(P2_add_958_n128), .IN1(P2_add_958_n127), 
        .IN2(P2_add_958_n130) );
  AND2X1 P2_add_958_U135 ( .IN1(P2_add_958_n127), .IN2(P2_add_958_n130), 
        .Q(P2_add_958_n129) );
  NOR2X0 P2_add_958_U134 ( .QN(P2_N3614), .IN1(P2_add_958_n128), 
        .IN2(P2_add_958_n129) );
  NAND2X0 P2_add_958_U133 ( .IN1(n7252), .IN2(P2_add_958_n127), 
        .QN(P2_add_958_n124) );
  OR2X1 P2_add_958_U132 ( .IN2(n7252), .IN1(P2_add_958_n127), 
        .Q(P2_add_958_n126) );
  NAND2X0 P2_add_958_U131 ( .IN1(P2_N3372), .IN2(P2_add_958_n126), 
        .QN(P2_add_958_n125) );
  NAND2X0 P2_add_958_U130 ( .IN1(P2_add_958_n124), .IN2(P2_add_958_n125), 
        .QN(P2_add_958_n117) );
  OR2X1 P2_add_958_U128 ( .IN2(P2_N3373), .IN1(n7248), .Q(P2_add_958_n121) );
  NAND2X0 P2_add_958_U127 ( .IN1(P2_N3373), .IN2(n7248), .QN(P2_add_958_n122)
         );
  NAND2X0 P2_add_958_U126 ( .IN1(P2_add_958_n121), .IN2(P2_add_958_n122), 
        .QN(P2_add_958_n120) );
  NOR2X0 P2_add_958_U125 ( .QN(P2_add_958_n118), .IN1(P2_add_958_n117), 
        .IN2(P2_add_958_n120) );
  AND2X1 P2_add_958_U124 ( .IN1(P2_add_958_n117), .IN2(P2_add_958_n120), 
        .Q(P2_add_958_n119) );
  NOR2X0 P2_add_958_U123 ( .QN(P2_N3615), .IN1(P2_add_958_n118), 
        .IN2(P2_add_958_n119) );
  NAND2X0 P2_add_958_U122 ( .IN1(P2_N5093), .IN2(P2_add_958_n117), 
        .QN(P2_add_958_n114) );
  OR2X1 P2_add_958_U121 ( .IN2(P2_N5093), .IN1(P2_add_958_n117), 
        .Q(P2_add_958_n116) );
  NAND2X0 P2_add_958_U120 ( .IN1(P2_N3373), .IN2(P2_add_958_n116), 
        .QN(P2_add_958_n115) );
  NAND2X0 P2_add_958_U119 ( .IN1(P2_add_958_n114), .IN2(P2_add_958_n115), 
        .QN(P2_add_958_n107) );
  OR2X1 P2_add_958_U117 ( .IN2(P2_N3374), .IN1(n7243), .Q(P2_add_958_n111) );
  NAND2X0 P2_add_958_U116 ( .IN1(P2_N3374), .IN2(n7243), .QN(P2_add_958_n112)
         );
  NAND2X0 P2_add_958_U115 ( .IN1(P2_add_958_n111), .IN2(P2_add_958_n112), 
        .QN(P2_add_958_n110) );
  NOR2X0 P2_add_958_U114 ( .QN(P2_add_958_n108), .IN1(P2_add_958_n107), 
        .IN2(P2_add_958_n110) );
  AND2X1 P2_add_958_U113 ( .IN1(P2_add_958_n107), .IN2(P2_add_958_n110), 
        .Q(P2_add_958_n109) );
  NOR2X0 P2_add_958_U112 ( .QN(P2_N3616), .IN1(P2_add_958_n108), 
        .IN2(P2_add_958_n109) );
  NAND2X0 P2_add_958_U111 ( .IN1(n7242), .IN2(P2_add_958_n107), 
        .QN(P2_add_958_n104) );
  OR2X1 P2_add_958_U110 ( .IN2(n7242), .IN1(P2_add_958_n107), 
        .Q(P2_add_958_n106) );
  NAND2X0 P2_add_958_U109 ( .IN1(P2_N3374), .IN2(P2_add_958_n106), 
        .QN(P2_add_958_n105) );
  NAND2X0 P2_add_958_U108 ( .IN1(P2_add_958_n104), .IN2(P2_add_958_n105), 
        .QN(P2_add_958_n97) );
  OR2X1 P2_add_958_U106 ( .IN2(P2_N3375), .IN1(n7239), .Q(P2_add_958_n101) );
  NAND2X0 P2_add_958_U105 ( .IN1(P2_N3375), .IN2(n7239), .QN(P2_add_958_n102)
         );
  NAND2X0 P2_add_958_U104 ( .IN1(P2_add_958_n101), .IN2(P2_add_958_n102), 
        .QN(P2_add_958_n100) );
  NOR2X0 P2_add_958_U103 ( .QN(P2_add_958_n98), .IN1(P2_add_958_n97), 
        .IN2(P2_add_958_n100) );
  AND2X1 P2_add_958_U102 ( .IN1(P2_add_958_n97), .IN2(P2_add_958_n100), 
        .Q(P2_add_958_n99) );
  NOR2X0 P2_add_958_U101 ( .QN(P2_N3617), .IN1(P2_add_958_n98), 
        .IN2(P2_add_958_n99) );
  NAND2X0 P2_add_958_U100 ( .IN1(P2_N5095), .IN2(P2_add_958_n97), 
        .QN(P2_add_958_n94) );
  OR2X1 P2_add_958_U99 ( .IN2(P2_N5095), .IN1(P2_add_958_n97), 
        .Q(P2_add_958_n96) );
  NAND2X0 P2_add_958_U98 ( .IN1(P2_N3375), .IN2(P2_add_958_n96), 
        .QN(P2_add_958_n95) );
  NAND2X0 P2_add_958_U97 ( .IN1(P2_add_958_n94), .IN2(P2_add_958_n95), 
        .QN(P2_add_958_n87) );
  OR2X1 P2_add_958_U95 ( .IN2(P2_N3376), .IN1(n7234), .Q(P2_add_958_n91) );
  NAND2X0 P2_add_958_U94 ( .IN1(P2_N3376), .IN2(n7234), .QN(P2_add_958_n92) );
  NAND2X0 P2_add_958_U93 ( .IN1(P2_add_958_n91), .IN2(P2_add_958_n92), 
        .QN(P2_add_958_n90) );
  NOR2X0 P2_add_958_U92 ( .QN(P2_add_958_n88), .IN1(P2_add_958_n87), 
        .IN2(P2_add_958_n90) );
  AND2X1 P2_add_958_U91 ( .IN1(P2_add_958_n87), .IN2(P2_add_958_n90), 
        .Q(P2_add_958_n89) );
  NOR2X0 P2_add_958_U90 ( .QN(P2_N3618), .IN1(P2_add_958_n88), 
        .IN2(P2_add_958_n89) );
  NAND2X0 P2_add_958_U89 ( .IN1(n7237), .IN2(P2_add_958_n87), 
        .QN(P2_add_958_n84) );
  OR2X1 P2_add_958_U88 ( .IN2(n7237), .IN1(P2_add_958_n87), .Q(P2_add_958_n86)
         );
  NAND2X0 P2_add_958_U87 ( .IN1(P2_N3376), .IN2(P2_add_958_n86), 
        .QN(P2_add_958_n85) );
  NAND2X0 P2_add_958_U86 ( .IN1(P2_add_958_n84), .IN2(P2_add_958_n85), 
        .QN(P2_add_958_n77) );
  OR2X1 P2_add_958_U84 ( .IN2(P2_N3377), .IN1(n7229), .Q(P2_add_958_n81) );
  NAND2X0 P2_add_958_U83 ( .IN1(P2_N3377), .IN2(n7229), .QN(P2_add_958_n82) );
  NAND2X0 P2_add_958_U82 ( .IN1(P2_add_958_n81), .IN2(P2_add_958_n82), 
        .QN(P2_add_958_n80) );
  NOR2X0 P2_add_958_U81 ( .QN(P2_add_958_n78), .IN1(P2_add_958_n77), 
        .IN2(P2_add_958_n80) );
  AND2X1 P2_add_958_U80 ( .IN1(P2_add_958_n77), .IN2(P2_add_958_n80), 
        .Q(P2_add_958_n79) );
  NOR2X0 P2_add_958_U79 ( .QN(P2_N3619), .IN1(P2_add_958_n78), 
        .IN2(P2_add_958_n79) );
  NAND2X0 P2_add_958_U78 ( .IN1(n7231), .IN2(P2_add_958_n77), 
        .QN(P2_add_958_n74) );
  OR2X1 P2_add_958_U77 ( .IN2(n7231), .IN1(P2_add_958_n77), .Q(P2_add_958_n76)
         );
  NAND2X0 P2_add_958_U76 ( .IN1(P2_N3377), .IN2(P2_add_958_n76), 
        .QN(P2_add_958_n75) );
  NAND2X0 P2_add_958_U75 ( .IN1(P2_add_958_n74), .IN2(P2_add_958_n75), 
        .QN(P2_add_958_n64) );
  OR2X1 P2_add_958_U73 ( .IN2(P2_N3378), .IN1(n7224), .Q(P2_add_958_n71) );
  NAND2X0 P2_add_958_U72 ( .IN1(P2_N3378), .IN2(n7224), .QN(P2_add_958_n72) );
  NAND2X0 P2_add_958_U71 ( .IN1(P2_add_958_n71), .IN2(P2_add_958_n72), 
        .QN(P2_add_958_n70) );
  NOR2X0 P2_add_958_U70 ( .QN(P2_add_958_n68), .IN1(P2_add_958_n64), 
        .IN2(P2_add_958_n70) );
  AND2X1 P2_add_958_U69 ( .IN1(P2_add_958_n64), .IN2(P2_add_958_n70), 
        .Q(P2_add_958_n69) );
  NOR2X0 P2_add_958_U68 ( .QN(P2_N3620), .IN1(P2_add_958_n68), 
        .IN2(P2_add_958_n69) );
  OR2X1 P2_add_958_U66 ( .IN2(P2_N3379), .IN1(n7222), .Q(P2_add_958_n65) );
  NAND2X0 P2_add_958_U65 ( .IN1(P2_N3379), .IN2(n7222), .QN(P2_add_958_n66) );
  NAND2X0 P2_add_958_U64 ( .IN1(P2_add_958_n65), .IN2(P2_add_958_n66), 
        .QN(P2_add_958_n60) );
  NAND2X0 P2_add_958_U63 ( .IN1(P2_N5098), .IN2(P2_add_958_n64), 
        .QN(P2_add_958_n61) );
  OR2X1 P2_add_958_U62 ( .IN2(P2_N5098), .IN1(P2_add_958_n64), 
        .Q(P2_add_958_n63) );
  NAND2X0 P2_add_958_U247 ( .IN1(P2_N3362), .IN2(P2_add_958_n233), 
        .QN(P2_add_958_n232) );
  NAND2X0 P2_add_958_U246 ( .IN1(P2_add_958_n231), .IN2(P2_add_958_n232), 
        .QN(P2_add_958_n224) );
  OR2X1 P2_add_958_U244 ( .IN2(P2_N3363), .IN1(n7211), .Q(P2_add_958_n228) );
  NAND2X0 P2_add_958_U243 ( .IN1(P2_N3363), .IN2(n7211), .QN(P2_add_958_n229)
         );
  NAND2X0 P2_add_958_U242 ( .IN1(P2_add_958_n228), .IN2(P2_add_958_n229), 
        .QN(P2_add_958_n227) );
  NOR2X0 P2_add_958_U241 ( .QN(P2_add_958_n225), .IN1(P2_add_958_n224), 
        .IN2(P2_add_958_n227) );
  AND2X1 P2_add_958_U240 ( .IN1(P2_add_958_n224), .IN2(P2_add_958_n227), 
        .Q(P2_add_958_n226) );
  NOR2X0 P2_add_958_U239 ( .QN(P2_N3605), .IN1(P2_add_958_n225), 
        .IN2(P2_add_958_n226) );
  NAND2X0 P2_add_958_U238 ( .IN1(n7210), .IN2(P2_add_958_n224), 
        .QN(P2_add_958_n221) );
  OR2X1 P2_add_958_U237 ( .IN2(n7210), .IN1(P2_add_958_n224), 
        .Q(P2_add_958_n223) );
  NAND2X0 P2_add_958_U236 ( .IN1(P2_N3363), .IN2(P2_add_958_n223), 
        .QN(P2_add_958_n222) );
  NAND2X0 P2_add_958_U235 ( .IN1(P2_add_958_n221), .IN2(P2_add_958_n222), 
        .QN(P2_add_958_n214) );
  OR2X1 P2_add_958_U233 ( .IN2(P2_N3364), .IN1(n7208), .Q(P2_add_958_n218) );
  NAND2X0 P2_add_958_U232 ( .IN1(P2_N3364), .IN2(n7208), .QN(P2_add_958_n219)
         );
  NAND2X0 P2_add_958_U231 ( .IN1(P2_add_958_n218), .IN2(P2_add_958_n219), 
        .QN(P2_add_958_n217) );
  NOR2X0 P2_add_958_U230 ( .QN(P2_add_958_n215), .IN1(P2_add_958_n214), 
        .IN2(P2_add_958_n217) );
  AND2X1 P2_add_958_U229 ( .IN1(P2_add_958_n214), .IN2(P2_add_958_n217), 
        .Q(P2_add_958_n216) );
  NOR2X0 P2_add_958_U228 ( .QN(P2_N3606), .IN1(P2_add_958_n215), 
        .IN2(P2_add_958_n216) );
  NAND2X0 P2_add_958_U227 ( .IN1(P2_N5084), .IN2(P2_add_958_n214), 
        .QN(P2_add_958_n211) );
  OR2X1 P2_add_958_U226 ( .IN2(P2_N5084), .IN1(P2_add_958_n214), 
        .Q(P2_add_958_n213) );
  NAND2X0 P2_add_958_U225 ( .IN1(P2_N3364), .IN2(P2_add_958_n213), 
        .QN(P2_add_958_n212) );
  NAND2X0 P2_add_958_U224 ( .IN1(P2_add_958_n211), .IN2(P2_add_958_n212), 
        .QN(P2_add_958_n204) );
  OR2X1 P2_add_958_U222 ( .IN2(P2_N3365), .IN1(n7205), .Q(P2_add_958_n208) );
  NAND2X0 P2_add_958_U221 ( .IN1(P2_N3365), .IN2(n7205), .QN(P2_add_958_n209)
         );
  NAND2X0 P2_add_958_U220 ( .IN1(P2_add_958_n208), .IN2(P2_add_958_n209), 
        .QN(P2_add_958_n207) );
  NOR2X0 P2_add_958_U219 ( .QN(P2_add_958_n205), .IN1(P2_add_958_n204), 
        .IN2(P2_add_958_n207) );
  AND2X1 P2_add_958_U218 ( .IN1(P2_add_958_n204), .IN2(P2_add_958_n207), 
        .Q(P2_add_958_n206) );
  NOR2X0 P2_add_958_U217 ( .QN(P2_N3607), .IN1(P2_add_958_n205), 
        .IN2(P2_add_958_n206) );
  NAND2X0 P2_add_958_U216 ( .IN1(P2_N5085), .IN2(P2_add_958_n204), 
        .QN(P2_add_958_n201) );
  OR2X1 P2_add_958_U215 ( .IN2(P2_N5085), .IN1(P2_add_958_n204), 
        .Q(P2_add_958_n203) );
  NAND2X0 P2_add_958_U214 ( .IN1(P2_N3365), .IN2(P2_add_958_n203), 
        .QN(P2_add_958_n202) );
  NAND2X0 P2_add_958_U213 ( .IN1(P2_add_958_n201), .IN2(P2_add_958_n202), 
        .QN(P2_add_958_n194) );
  OR2X1 P2_add_958_U211 ( .IN2(P2_N3366), .IN1(n7201), .Q(P2_add_958_n198) );
  NAND2X0 P2_add_958_U210 ( .IN1(P2_N3366), .IN2(n7201), .QN(P2_add_958_n199)
         );
  NAND2X0 P2_add_958_U209 ( .IN1(P2_add_958_n198), .IN2(P2_add_958_n199), 
        .QN(P2_add_958_n197) );
  NOR2X0 P2_add_958_U208 ( .QN(P2_add_958_n195), .IN1(P2_add_958_n194), 
        .IN2(P2_add_958_n197) );
  AND2X1 P2_add_958_U207 ( .IN1(P2_add_958_n194), .IN2(P2_add_958_n197), 
        .Q(P2_add_958_n196) );
  NOR2X0 P2_add_958_U206 ( .QN(P2_N3608), .IN1(P2_add_958_n195), 
        .IN2(P2_add_958_n196) );
  NAND2X0 P2_add_958_U205 ( .IN1(P2_N5086), .IN2(P2_add_958_n194), 
        .QN(P2_add_958_n191) );
  OR2X1 P2_add_958_U204 ( .IN2(P2_N5086), .IN1(P2_add_958_n194), 
        .Q(P2_add_958_n193) );
  NAND2X0 P2_add_958_U203 ( .IN1(P2_N3366), .IN2(P2_add_958_n193), 
        .QN(P2_add_958_n192) );
  NAND2X0 P2_add_958_U202 ( .IN1(P2_add_958_n191), .IN2(P2_add_958_n192), 
        .QN(P2_add_958_n184) );
  OR2X1 P2_add_958_U200 ( .IN2(P2_N3367), .IN1(n7197), .Q(P2_add_958_n188) );
  NAND2X0 P2_add_958_U199 ( .IN1(P2_N3367), .IN2(n7197), .QN(P2_add_958_n189)
         );
  NAND2X0 P2_add_958_U198 ( .IN1(P2_add_958_n188), .IN2(P2_add_958_n189), 
        .QN(P2_add_958_n187) );
  NOR2X0 P2_add_958_U197 ( .QN(P2_add_958_n185), .IN1(P2_add_958_n184), 
        .IN2(P2_add_958_n187) );
  AND2X1 P2_add_958_U196 ( .IN1(P2_add_958_n184), .IN2(P2_add_958_n187), 
        .Q(P2_add_958_n186) );
  NOR2X0 P2_add_958_U195 ( .QN(P2_N3609), .IN1(P2_add_958_n185), 
        .IN2(P2_add_958_n186) );
  NAND2X0 P2_add_958_U194 ( .IN1(n7198), .IN2(P2_add_958_n184), 
        .QN(P2_add_958_n181) );
  OR2X1 P2_add_958_U193 ( .IN2(n7198), .IN1(P2_add_958_n184), 
        .Q(P2_add_958_n183) );
  NAND2X0 P2_add_958_U192 ( .IN1(P2_N3367), .IN2(P2_add_958_n183), 
        .QN(P2_add_958_n182) );
  NAND2X0 P2_add_958_U191 ( .IN1(P2_add_958_n181), .IN2(P2_add_958_n182), 
        .QN(P2_add_958_n174) );
  OR2X1 P2_add_958_U189 ( .IN2(P2_N3368), .IN1(n7195), .Q(P2_add_958_n178) );
  NAND2X0 P2_add_958_U188 ( .IN1(P2_N3368), .IN2(n7195), .QN(P2_add_958_n179)
         );
  NAND2X0 P2_add_958_U187 ( .IN1(P2_add_958_n178), .IN2(P2_add_958_n179), 
        .QN(P2_add_958_n177) );
  NOR2X0 P2_add_958_U186 ( .QN(P2_add_958_n175), .IN1(P2_add_958_n174), 
        .IN2(P2_add_958_n177) );
  AND2X1 P2_add_958_U185 ( .IN1(P2_add_958_n174), .IN2(P2_add_958_n177), 
        .Q(P2_add_958_n176) );
  NOR2X0 P2_add_958_U184 ( .QN(P2_N3610), .IN1(P2_add_958_n175), 
        .IN2(P2_add_958_n176) );
  NAND2X0 P2_add_958_U183 ( .IN1(n7194), .IN2(P2_add_958_n174), 
        .QN(P2_add_958_n171) );
  OR2X1 P2_add_958_U182 ( .IN2(n7194), .IN1(P2_add_958_n174), 
        .Q(P2_add_958_n173) );
  NAND2X0 P2_add_958_U181 ( .IN1(P2_N3368), .IN2(P2_add_958_n173), 
        .QN(P2_add_958_n172) );
  NAND2X0 P2_add_958_U180 ( .IN1(P2_add_958_n171), .IN2(P2_add_958_n172), 
        .QN(P2_add_958_n164) );
  OR2X1 P2_add_958_U178 ( .IN2(P2_N3369), .IN1(n7188), .Q(P2_add_958_n168) );
  NAND2X0 P2_add_958_U177 ( .IN1(P2_N3369), .IN2(n7188), .QN(P2_add_958_n169)
         );
  NAND2X0 P2_add_958_U176 ( .IN1(P2_add_958_n168), .IN2(P2_add_958_n169), 
        .QN(P2_add_958_n167) );
  NOR2X0 P2_add_958_U175 ( .QN(P2_add_958_n165), .IN1(P2_add_958_n164), 
        .IN2(P2_add_958_n167) );
  AND2X1 P2_add_958_U174 ( .IN1(P2_add_958_n164), .IN2(P2_add_958_n167), 
        .Q(P2_add_958_n166) );
  NOR2X0 P2_add_958_U173 ( .QN(P2_N3611), .IN1(P2_add_958_n165), 
        .IN2(P2_add_958_n166) );
  NAND2X0 P2_add_958_U172 ( .IN1(P2_N5089), .IN2(P2_add_958_n164), 
        .QN(P2_add_958_n161) );
  OR2X1 P2_add_958_U171 ( .IN2(P2_N5089), .IN1(P2_add_958_n164), 
        .Q(P2_add_958_n163) );
  NAND2X0 P2_add_958_U170 ( .IN1(P2_N3369), .IN2(P2_add_958_n163), 
        .QN(P2_add_958_n162) );
  NAND2X0 P2_add_958_U169 ( .IN1(P2_add_958_n161), .IN2(P2_add_958_n162), 
        .QN(P2_add_958_n147) );
  OR2X1 P2_add_958_U167 ( .IN2(P2_N3370), .IN1(n7264), .Q(P2_add_958_n158) );
  NAND2X0 P2_add_958_U166 ( .IN1(P2_N3370), .IN2(n7264), .QN(P2_add_958_n159)
         );
  NAND2X0 P2_add_958_U165 ( .IN1(P2_add_958_n158), .IN2(P2_add_958_n159), 
        .QN(P2_add_958_n157) );
  NOR2X0 P2_add_958_U164 ( .QN(P2_add_958_n155), .IN1(P2_add_958_n147), 
        .IN2(P2_add_958_n157) );
  AND2X1 P2_add_958_U163 ( .IN1(P2_add_958_n147), .IN2(P2_add_958_n157), 
        .Q(P2_add_958_n156) );
  NOR2X0 P2_add_958_U162 ( .QN(P2_N3612), .IN1(P2_add_958_n155), 
        .IN2(P2_add_958_n156) );
  OR2X1 P2_add_958_U161 ( .IN2(P2_N3352), .IN1(n7184), .Q(P2_add_958_n152) );
  NAND2X0 P2_add_958_U160 ( .IN1(P2_N3352), .IN2(n7184), .QN(P2_add_958_n153)
         );
  NAND2X0 P2_add_958_U159 ( .IN1(P2_add_958_n152), .IN2(P2_add_958_n153), 
        .QN(P2_add_958_n150) );
  NAND2X0 P2_add_958_U158 ( .IN1(P2_add_958_n150), .IN2(P2_add_958_n151), 
        .QN(P2_add_958_n148) );
  OR2X1 P2_add_958_U157 ( .IN2(P2_add_958_n151), .IN1(P2_add_958_n150), 
        .Q(P2_add_958_n149) );
  NAND2X0 P2_add_958_U156 ( .IN1(P2_add_958_n148), .IN2(P2_add_958_n149), 
        .QN(P2_N3594) );
  NAND2X0 P2_add_958_U155 ( .IN1(P2_N5090), .IN2(P2_add_958_n147), 
        .QN(P2_add_958_n144) );
  OR2X1 P2_add_958_U308 ( .IN2(P2_N3351), .IN1(n2919), .Q(P2_add_958_n278) );
  NAND2X0 P2_add_958_U307 ( .IN1(P2_N3351), .IN2(n2919), .QN(P2_add_958_n279)
         );
  NAND2X0 P2_add_958_U306 ( .IN1(P2_add_958_n278), .IN2(P2_add_958_n279), 
        .QN(P2_N3593) );
  NAND2X0 P2_add_958_U304 ( .IN1(P2_N3351), .IN2(n7035), .QN(P2_add_958_n151)
         );
  OR2X1 P2_add_958_U303 ( .IN2(P2_add_958_n151), .IN1(n7184), 
        .Q(P2_add_958_n275) );
  NAND2X0 P2_add_958_U302 ( .IN1(n7184), .IN2(P2_add_958_n151), 
        .QN(P2_add_958_n277) );
  NAND2X0 P2_add_958_U301 ( .IN1(P2_N3352), .IN2(P2_add_958_n277), 
        .QN(P2_add_958_n276) );
  NAND2X0 P2_add_958_U300 ( .IN1(P2_add_958_n275), .IN2(P2_add_958_n276), 
        .QN(P2_add_958_n52) );
  NAND2X0 P2_add_958_U299 ( .IN1(P2_N5073), .IN2(P2_add_958_n52), 
        .QN(P2_add_958_n272) );
  OR2X1 P2_add_958_U298 ( .IN2(P2_N5073), .IN1(P2_add_958_n52), 
        .Q(P2_add_958_n274) );
  NAND2X0 P2_add_958_U297 ( .IN1(P2_N3353), .IN2(P2_add_958_n274), 
        .QN(P2_add_958_n273) );
  NAND2X0 P2_add_958_U296 ( .IN1(P2_add_958_n272), .IN2(P2_add_958_n273), 
        .QN(P2_add_958_n45) );
  NAND2X0 P2_add_958_U295 ( .IN1(P2_N5074), .IN2(P2_add_958_n45), 
        .QN(P2_add_958_n269) );
  OR2X1 P2_add_958_U294 ( .IN2(P2_N5074), .IN1(P2_add_958_n45), 
        .Q(P2_add_958_n271) );
  NAND2X0 P2_add_958_U293 ( .IN1(P2_N3354), .IN2(P2_add_958_n271), 
        .QN(P2_add_958_n270) );
  NAND2X0 P2_add_958_U292 ( .IN1(P2_add_958_n269), .IN2(P2_add_958_n270), 
        .QN(P2_add_958_n38) );
  NAND2X0 P2_add_958_U291 ( .IN1(P2_N5075), .IN2(P2_add_958_n38), 
        .QN(P2_add_958_n266) );
  OR2X1 P2_add_958_U290 ( .IN2(P2_N5075), .IN1(P2_add_958_n38), 
        .Q(P2_add_958_n268) );
  NAND2X0 P2_add_958_U289 ( .IN1(P2_N3355), .IN2(P2_add_958_n268), 
        .QN(P2_add_958_n267) );
  NAND2X0 P2_add_958_U288 ( .IN1(P2_add_958_n266), .IN2(P2_add_958_n267), 
        .QN(P2_add_958_n31) );
  NAND2X0 P2_add_958_U287 ( .IN1(n7165), .IN2(P2_add_958_n31), 
        .QN(P2_add_958_n263) );
  OR2X1 P2_add_958_U286 ( .IN2(n7165), .IN1(P2_add_958_n31), 
        .Q(P2_add_958_n265) );
  NAND2X0 P2_add_958_U285 ( .IN1(P2_N3356), .IN2(P2_add_958_n265), 
        .QN(P2_add_958_n264) );
  NAND2X0 P2_add_958_U284 ( .IN1(P2_add_958_n263), .IN2(P2_add_958_n264), 
        .QN(P2_add_958_n24) );
  NAND2X0 P2_add_958_U283 ( .IN1(P2_N5077), .IN2(P2_add_958_n24), 
        .QN(P2_add_958_n260) );
  OR2X1 P2_add_958_U282 ( .IN2(P2_N5077), .IN1(P2_add_958_n24), 
        .Q(P2_add_958_n262) );
  NAND2X0 P2_add_958_U281 ( .IN1(P2_N3357), .IN2(P2_add_958_n262), 
        .QN(P2_add_958_n261) );
  NAND2X0 P2_add_958_U280 ( .IN1(P2_add_958_n260), .IN2(P2_add_958_n261), 
        .QN(P2_add_958_n17) );
  NAND2X0 P2_add_958_U279 ( .IN1(n7158), .IN2(P2_add_958_n17), 
        .QN(P2_add_958_n257) );
  OR2X1 P2_add_958_U278 ( .IN2(n7158), .IN1(P2_add_958_n17), 
        .Q(P2_add_958_n259) );
  NAND2X0 P2_add_958_U277 ( .IN1(P2_N3358), .IN2(P2_add_958_n259), 
        .QN(P2_add_958_n258) );
  NAND2X0 P2_add_958_U276 ( .IN1(P2_add_958_n257), .IN2(P2_add_958_n258), 
        .QN(P2_add_958_n10) );
  NAND2X0 P2_add_958_U275 ( .IN1(P2_N5079), .IN2(P2_add_958_n10), 
        .QN(P2_add_958_n254) );
  OR2X1 P2_add_958_U274 ( .IN2(P2_N5079), .IN1(P2_add_958_n10), 
        .Q(P2_add_958_n256) );
  NAND2X0 P2_add_958_U273 ( .IN1(P2_N3359), .IN2(P2_add_958_n256), 
        .QN(P2_add_958_n255) );
  NAND2X0 P2_add_958_U272 ( .IN1(P2_add_958_n254), .IN2(P2_add_958_n255), 
        .QN(P2_add_958_n3) );
  NAND2X0 P2_add_958_U271 ( .IN1(P2_N5080), .IN2(P2_add_958_n3), 
        .QN(P2_add_958_n251) );
  OR2X1 P2_add_958_U270 ( .IN2(P2_N5080), .IN1(P2_add_958_n3), 
        .Q(P2_add_958_n253) );
  NAND2X0 P2_add_958_U269 ( .IN1(P2_N3360), .IN2(P2_add_958_n253), 
        .QN(P2_add_958_n252) );
  NAND2X0 P2_add_958_U268 ( .IN1(P2_add_958_n251), .IN2(P2_add_958_n252), 
        .QN(P2_add_958_n244) );
  OR2X1 P2_add_958_U266 ( .IN2(P2_N3361), .IN1(n7219), .Q(P2_add_958_n248) );
  NAND2X0 P2_add_958_U265 ( .IN1(P2_N3361), .IN2(n7219), .QN(P2_add_958_n249)
         );
  NAND2X0 P2_add_958_U264 ( .IN1(P2_add_958_n248), .IN2(P2_add_958_n249), 
        .QN(P2_add_958_n247) );
  NOR2X0 P2_add_958_U263 ( .QN(P2_add_958_n245), .IN1(P2_add_958_n244), 
        .IN2(P2_add_958_n247) );
  AND2X1 P2_add_958_U262 ( .IN1(P2_add_958_n244), .IN2(P2_add_958_n247), 
        .Q(P2_add_958_n246) );
  NOR2X0 P2_add_958_U261 ( .QN(P2_N3603), .IN1(P2_add_958_n245), 
        .IN2(P2_add_958_n246) );
  NAND2X0 P2_add_958_U260 ( .IN1(P2_N5081), .IN2(P2_add_958_n244), 
        .QN(P2_add_958_n241) );
  OR2X1 P2_add_958_U259 ( .IN2(P2_N5081), .IN1(P2_add_958_n244), 
        .Q(P2_add_958_n243) );
  NAND2X0 P2_add_958_U258 ( .IN1(P2_N3361), .IN2(P2_add_958_n243), 
        .QN(P2_add_958_n242) );
  NAND2X0 P2_add_958_U257 ( .IN1(P2_add_958_n241), .IN2(P2_add_958_n242), 
        .QN(P2_add_958_n234) );
  OR2X1 P2_add_958_U255 ( .IN2(P2_N3362), .IN1(n7214), .Q(P2_add_958_n238) );
  NAND2X0 P2_add_958_U254 ( .IN1(P2_N3362), .IN2(n7214), .QN(P2_add_958_n239)
         );
  NAND2X0 P2_add_958_U253 ( .IN1(P2_add_958_n238), .IN2(P2_add_958_n239), 
        .QN(P2_add_958_n237) );
  NOR2X0 P2_add_958_U252 ( .QN(P2_add_958_n235), .IN1(P2_add_958_n234), 
        .IN2(P2_add_958_n237) );
  AND2X1 P2_add_958_U251 ( .IN1(P2_add_958_n234), .IN2(P2_add_958_n237), 
        .Q(P2_add_958_n236) );
  NOR2X0 P2_add_958_U250 ( .QN(P2_N3604), .IN1(P2_add_958_n235), 
        .IN2(P2_add_958_n236) );
  NAND2X0 P2_add_958_U249 ( .IN1(n7216), .IN2(P2_add_958_n234), 
        .QN(P2_add_958_n231) );
  OR2X1 P2_add_958_U248 ( .IN2(n7216), .IN1(P2_add_958_n234), 
        .Q(P2_add_958_n233) );
  INVX0 P2_sub_978_U92 ( .ZN(P2_sub_978_n85), .INP(P2_N3749) );
  NAND2X0 P2_sub_978_U91 ( .IN1(n7237), .IN2(P2_sub_978_n85), 
        .QN(P2_sub_978_n97) );
  OR2X1 P2_sub_978_U90 ( .IN2(n7237), .IN1(P2_sub_978_n85), .Q(P2_sub_978_n98)
         );
  NAND2X0 P2_sub_978_U89 ( .IN1(P2_sub_978_n97), .IN2(P2_sub_978_n98), 
        .QN(P2_sub_978_n91) );
  NAND2X0 P2_sub_978_U88 ( .IN1(n7238), .IN2(P2_sub_978_n96), 
        .QN(P2_sub_978_n92) );
  OR2X1 P2_sub_978_U87 ( .IN2(n7238), .IN1(P2_sub_978_n96), .Q(P2_sub_978_n94)
         );
  NAND2X0 P2_sub_978_U86 ( .IN1(P2_sub_978_n94), .IN2(P2_sub_978_n95), 
        .QN(P2_sub_978_n93) );
  NAND2X0 P2_sub_978_U85 ( .IN1(P2_sub_978_n92), .IN2(P2_sub_978_n93), 
        .QN(P2_sub_978_n86) );
  NAND2X0 P2_sub_978_U84 ( .IN1(P2_sub_978_n91), .IN2(P2_sub_978_n86), 
        .QN(P2_sub_978_n89) );
  OR2X1 P2_sub_978_U83 ( .IN2(P2_sub_978_n86), .IN1(P2_sub_978_n91), 
        .Q(P2_sub_978_n90) );
  NAND2X0 P2_sub_978_U82 ( .IN1(P2_sub_978_n89), .IN2(P2_sub_978_n90), 
        .QN(P2_N3991) );
  INVX0 P2_sub_978_U81 ( .ZN(P2_sub_978_n75), .INP(P2_N3750) );
  NAND2X0 P2_sub_978_U80 ( .IN1(n7231), .IN2(P2_sub_978_n75), 
        .QN(P2_sub_978_n87) );
  OR2X1 P2_sub_978_U79 ( .IN2(n7231), .IN1(P2_sub_978_n75), .Q(P2_sub_978_n88)
         );
  NAND2X0 P2_sub_978_U78 ( .IN1(P2_sub_978_n87), .IN2(P2_sub_978_n88), 
        .QN(P2_sub_978_n81) );
  NAND2X0 P2_sub_978_U77 ( .IN1(n7237), .IN2(P2_sub_978_n86), 
        .QN(P2_sub_978_n82) );
  OR2X1 P2_sub_978_U76 ( .IN2(n7237), .IN1(P2_sub_978_n86), .Q(P2_sub_978_n84)
         );
  NAND2X0 P2_sub_978_U75 ( .IN1(P2_sub_978_n84), .IN2(P2_sub_978_n85), 
        .QN(P2_sub_978_n83) );
  NAND2X0 P2_sub_978_U74 ( .IN1(P2_sub_978_n82), .IN2(P2_sub_978_n83), 
        .QN(P2_sub_978_n76) );
  NAND2X0 P2_sub_978_U73 ( .IN1(P2_sub_978_n81), .IN2(P2_sub_978_n76), 
        .QN(P2_sub_978_n79) );
  OR2X1 P2_sub_978_U72 ( .IN2(P2_sub_978_n76), .IN1(P2_sub_978_n81), 
        .Q(P2_sub_978_n80) );
  NAND2X0 P2_sub_978_U71 ( .IN1(P2_sub_978_n79), .IN2(P2_sub_978_n80), 
        .QN(P2_N3992) );
  INVX0 P2_sub_978_U70 ( .ZN(P2_sub_978_n64), .INP(P2_N3751) );
  NAND2X0 P2_sub_978_U69 ( .IN1(P2_N5098), .IN2(P2_sub_978_n64), 
        .QN(P2_sub_978_n77) );
  OR2X1 P2_sub_978_U68 ( .IN2(P2_N5098), .IN1(P2_sub_978_n64), 
        .Q(P2_sub_978_n78) );
  NAND2X0 P2_sub_978_U67 ( .IN1(P2_sub_978_n77), .IN2(P2_sub_978_n78), 
        .QN(P2_sub_978_n71) );
  NAND2X0 P2_sub_978_U66 ( .IN1(n7231), .IN2(P2_sub_978_n76), 
        .QN(P2_sub_978_n72) );
  OR2X1 P2_sub_978_U65 ( .IN2(n7231), .IN1(P2_sub_978_n76), .Q(P2_sub_978_n74)
         );
  NAND2X0 P2_sub_978_U64 ( .IN1(P2_sub_978_n74), .IN2(P2_sub_978_n75), 
        .QN(P2_sub_978_n73) );
  NAND2X0 P2_sub_978_U63 ( .IN1(P2_sub_978_n72), .IN2(P2_sub_978_n73), 
        .QN(P2_sub_978_n65) );
  NAND2X0 P2_sub_978_U62 ( .IN1(P2_sub_978_n71), .IN2(P2_sub_978_n65), 
        .QN(P2_sub_978_n69) );
  OR2X1 P2_sub_978_U61 ( .IN2(P2_sub_978_n65), .IN1(P2_sub_978_n71), 
        .Q(P2_sub_978_n70) );
  NAND2X0 P2_sub_978_U60 ( .IN1(P2_sub_978_n69), .IN2(P2_sub_978_n70), 
        .QN(P2_N3993) );
  OR2X1 P2_sub_978_U58 ( .IN2(P2_N3752), .IN1(n7222), .Q(P2_sub_978_n66) );
  NAND2X0 P2_sub_978_U57 ( .IN1(P2_N3752), .IN2(n7222), .QN(P2_sub_978_n67) );
  NAND2X0 P2_sub_978_U56 ( .IN1(P2_sub_978_n66), .IN2(P2_sub_978_n67), 
        .QN(P2_sub_978_n60) );
  NAND2X0 P2_sub_978_U55 ( .IN1(P2_N5098), .IN2(P2_sub_978_n65), 
        .QN(P2_sub_978_n61) );
  OR2X1 P2_sub_978_U54 ( .IN2(P2_N5098), .IN1(P2_sub_978_n65), 
        .Q(P2_sub_978_n63) );
  NAND2X0 P2_sub_978_U53 ( .IN1(P2_sub_978_n63), .IN2(P2_sub_978_n64), 
        .QN(P2_sub_978_n62) );
  NAND2X0 P2_sub_978_U52 ( .IN1(P2_sub_978_n61), .IN2(P2_sub_978_n62), 
        .QN(P2_sub_978_n59) );
  NAND2X0 P2_sub_978_U51 ( .IN1(P2_sub_978_n60), .IN2(P2_sub_978_n59), 
        .QN(P2_sub_978_n57) );
  OR2X1 P2_sub_978_U50 ( .IN2(P2_sub_978_n60), .IN1(P2_sub_978_n59), 
        .Q(P2_sub_978_n58) );
  NAND2X0 P2_sub_978_U49 ( .IN1(P2_sub_978_n57), .IN2(P2_sub_978_n58), 
        .QN(P2_N3994) );
  NAND2X0 P2_sub_978_U48 ( .IN1(n7181), .IN2(P2_sub_978_n56), 
        .QN(P2_sub_978_n54) );
  OR2X1 P2_sub_978_U47 ( .IN2(n7181), .IN1(P2_sub_978_n56), .Q(P2_sub_978_n55)
         );
  NAND2X0 P2_sub_978_U46 ( .IN1(P2_sub_978_n54), .IN2(P2_sub_978_n55), 
        .QN(P2_sub_978_n52) );
  NAND2X0 P2_sub_978_U45 ( .IN1(P2_sub_978_n52), .IN2(P2_sub_978_n53), 
        .QN(P2_sub_978_n50) );
  OR2X1 P2_sub_978_U44 ( .IN2(P2_sub_978_n53), .IN1(P2_sub_978_n52), 
        .Q(P2_sub_978_n51) );
  NAND2X0 P2_sub_978_U43 ( .IN1(P2_sub_978_n50), .IN2(P2_sub_978_n51), 
        .QN(P2_N3968) );
  NAND2X0 P2_sub_978_U42 ( .IN1(n7177), .IN2(P2_sub_978_n49), 
        .QN(P2_sub_978_n47) );
  OR2X1 P2_sub_978_U41 ( .IN2(n7177), .IN1(P2_sub_978_n49), .Q(P2_sub_978_n48)
         );
  NAND2X0 P2_sub_978_U40 ( .IN1(P2_sub_978_n47), .IN2(P2_sub_978_n48), 
        .QN(P2_sub_978_n45) );
  NAND2X0 P2_sub_978_U39 ( .IN1(P2_sub_978_n45), .IN2(P2_sub_978_n46), 
        .QN(P2_sub_978_n43) );
  OR2X1 P2_sub_978_U38 ( .IN2(P2_sub_978_n46), .IN1(P2_sub_978_n45), 
        .Q(P2_sub_978_n44) );
  NAND2X0 P2_sub_978_U37 ( .IN1(P2_sub_978_n43), .IN2(P2_sub_978_n44), 
        .QN(P2_N3969) );
  NAND2X0 P2_sub_978_U36 ( .IN1(n7173), .IN2(P2_sub_978_n42), 
        .QN(P2_sub_978_n40) );
  OR2X1 P2_sub_978_U35 ( .IN2(n7173), .IN1(P2_sub_978_n42), .Q(P2_sub_978_n41)
         );
  NAND2X0 P2_sub_978_U34 ( .IN1(P2_sub_978_n40), .IN2(P2_sub_978_n41), 
        .QN(P2_sub_978_n38) );
  NAND2X0 P2_sub_978_U33 ( .IN1(P2_sub_978_n38), .IN2(P2_sub_978_n39), 
        .QN(P2_sub_978_n36) );
  OR2X1 P2_sub_978_U32 ( .IN2(P2_sub_978_n39), .IN1(P2_sub_978_n38), 
        .Q(P2_sub_978_n37) );
  NAND2X0 P2_sub_978_U31 ( .IN1(P2_sub_978_n36), .IN2(P2_sub_978_n37), 
        .QN(P2_N3970) );
  NAND2X0 P2_sub_978_U30 ( .IN1(P2_N5076), .IN2(P2_sub_978_n35), 
        .QN(P2_sub_978_n33) );
  OR2X1 P2_sub_978_U29 ( .IN2(P2_N5076), .IN1(P2_sub_978_n35), 
        .Q(P2_sub_978_n34) );
  NAND2X0 P2_sub_978_U28 ( .IN1(P2_sub_978_n33), .IN2(P2_sub_978_n34), 
        .QN(P2_sub_978_n31) );
  NAND2X0 P2_sub_978_U27 ( .IN1(P2_sub_978_n31), .IN2(P2_sub_978_n32), 
        .QN(P2_sub_978_n29) );
  OR2X1 P2_sub_978_U26 ( .IN2(P2_sub_978_n32), .IN1(P2_sub_978_n31), 
        .Q(P2_sub_978_n30) );
  NAND2X0 P2_sub_978_U25 ( .IN1(P2_sub_978_n29), .IN2(P2_sub_978_n30), 
        .QN(P2_N3971) );
  NAND2X0 P2_sub_978_U24 ( .IN1(P2_N5077), .IN2(P2_sub_978_n28), 
        .QN(P2_sub_978_n26) );
  OR2X1 P2_sub_978_U23 ( .IN2(P2_N5077), .IN1(P2_sub_978_n28), 
        .Q(P2_sub_978_n27) );
  NAND2X0 P2_sub_978_U22 ( .IN1(P2_sub_978_n26), .IN2(P2_sub_978_n27), 
        .QN(P2_sub_978_n24) );
  NAND2X0 P2_sub_978_U21 ( .IN1(P2_sub_978_n24), .IN2(P2_sub_978_n25), 
        .QN(P2_sub_978_n22) );
  OR2X1 P2_sub_978_U20 ( .IN2(P2_sub_978_n25), .IN1(P2_sub_978_n24), 
        .Q(P2_sub_978_n23) );
  NAND2X0 P2_sub_978_U19 ( .IN1(P2_sub_978_n22), .IN2(P2_sub_978_n23), 
        .QN(P2_N3972) );
  NAND2X0 P2_sub_978_U18 ( .IN1(n7158), .IN2(P2_sub_978_n21), 
        .QN(P2_sub_978_n19) );
  OR2X1 P2_sub_978_U17 ( .IN2(n7158), .IN1(P2_sub_978_n21), .Q(P2_sub_978_n20)
         );
  NAND2X0 P2_sub_978_U16 ( .IN1(P2_sub_978_n19), .IN2(P2_sub_978_n20), 
        .QN(P2_sub_978_n17) );
  NAND2X0 P2_sub_978_U15 ( .IN1(P2_sub_978_n17), .IN2(P2_sub_978_n18), 
        .QN(P2_sub_978_n15) );
  OR2X1 P2_sub_978_U14 ( .IN2(P2_sub_978_n18), .IN1(P2_sub_978_n17), 
        .Q(P2_sub_978_n16) );
  NAND2X0 P2_sub_978_U13 ( .IN1(P2_sub_978_n15), .IN2(P2_sub_978_n16), 
        .QN(P2_N3973) );
  NAND2X0 P2_sub_978_U12 ( .IN1(n7154), .IN2(P2_sub_978_n14), 
        .QN(P2_sub_978_n12) );
  OR2X1 P2_sub_978_U11 ( .IN2(n7154), .IN1(P2_sub_978_n14), .Q(P2_sub_978_n13)
         );
  NAND2X0 P2_sub_978_U10 ( .IN1(P2_sub_978_n12), .IN2(P2_sub_978_n13), 
        .QN(P2_sub_978_n10) );
  NAND2X0 P2_sub_978_U9 ( .IN1(P2_sub_978_n10), .IN2(P2_sub_978_n11), 
        .QN(P2_sub_978_n8) );
  OR2X1 P2_sub_978_U8 ( .IN2(P2_sub_978_n11), .IN1(P2_sub_978_n10), 
        .Q(P2_sub_978_n9) );
  NAND2X0 P2_sub_978_U7 ( .IN1(P2_sub_978_n8), .IN2(P2_sub_978_n9), 
        .QN(P2_N3974) );
  NAND2X0 P2_sub_978_U6 ( .IN1(n7151), .IN2(P2_sub_978_n7), .QN(P2_sub_978_n5)
         );
  OR2X1 P2_sub_978_U5 ( .IN2(n7151), .IN1(P2_sub_978_n7), .Q(P2_sub_978_n6) );
  NAND2X0 P2_sub_978_U4 ( .IN1(P2_sub_978_n5), .IN2(P2_sub_978_n6), 
        .QN(P2_sub_978_n3) );
  NAND2X0 P2_sub_978_U3 ( .IN1(P2_sub_978_n3), .IN2(P2_sub_978_n4), 
        .QN(P2_sub_978_n1) );
  OR2X1 P2_sub_978_U2 ( .IN2(P2_sub_978_n4), .IN1(P2_sub_978_n3), 
        .Q(P2_sub_978_n2) );
  NAND2X0 P2_sub_978_U1 ( .IN1(P2_sub_978_n1), .IN2(P2_sub_978_n2), 
        .QN(P2_N3975) );
  NAND2X0 P2_sub_978_U185 ( .IN1(n7194), .IN2(P2_sub_978_n173), 
        .QN(P2_sub_978_n185) );
  OR2X1 P2_sub_978_U184 ( .IN2(n7194), .IN1(P2_sub_978_n173), 
        .Q(P2_sub_978_n186) );
  NAND2X0 P2_sub_978_U183 ( .IN1(P2_sub_978_n185), .IN2(P2_sub_978_n186), 
        .QN(P2_sub_978_n179) );
  NAND2X0 P2_sub_978_U182 ( .IN1(P2_N5087), .IN2(P2_sub_978_n184), 
        .QN(P2_sub_978_n180) );
  OR2X1 P2_sub_978_U181 ( .IN2(P2_N5087), .IN1(P2_sub_978_n184), 
        .Q(P2_sub_978_n182) );
  NAND2X0 P2_sub_978_U180 ( .IN1(P2_sub_978_n182), .IN2(P2_sub_978_n183), 
        .QN(P2_sub_978_n181) );
  NAND2X0 P2_sub_978_U179 ( .IN1(P2_sub_978_n180), .IN2(P2_sub_978_n181), 
        .QN(P2_sub_978_n174) );
  NAND2X0 P2_sub_978_U178 ( .IN1(P2_sub_978_n179), .IN2(P2_sub_978_n174), 
        .QN(P2_sub_978_n177) );
  OR2X1 P2_sub_978_U177 ( .IN2(P2_sub_978_n174), .IN1(P2_sub_978_n179), 
        .Q(P2_sub_978_n178) );
  NAND2X0 P2_sub_978_U176 ( .IN1(P2_sub_978_n177), .IN2(P2_sub_978_n178), 
        .QN(P2_N3983) );
  INVX0 P2_sub_978_U175 ( .ZN(P2_sub_978_n163), .INP(P2_N3742) );
  NAND2X0 P2_sub_978_U174 ( .IN1(n7187), .IN2(P2_sub_978_n163), 
        .QN(P2_sub_978_n175) );
  OR2X1 P2_sub_978_U173 ( .IN2(n7187), .IN1(P2_sub_978_n163), 
        .Q(P2_sub_978_n176) );
  NAND2X0 P2_sub_978_U172 ( .IN1(P2_sub_978_n175), .IN2(P2_sub_978_n176), 
        .QN(P2_sub_978_n169) );
  NAND2X0 P2_sub_978_U171 ( .IN1(n7194), .IN2(P2_sub_978_n174), 
        .QN(P2_sub_978_n170) );
  OR2X1 P2_sub_978_U170 ( .IN2(n7194), .IN1(P2_sub_978_n174), 
        .Q(P2_sub_978_n172) );
  NAND2X0 P2_sub_978_U169 ( .IN1(P2_sub_978_n172), .IN2(P2_sub_978_n173), 
        .QN(P2_sub_978_n171) );
  NAND2X0 P2_sub_978_U168 ( .IN1(P2_sub_978_n170), .IN2(P2_sub_978_n171), 
        .QN(P2_sub_978_n164) );
  NAND2X0 P2_sub_978_U167 ( .IN1(P2_sub_978_n169), .IN2(P2_sub_978_n164), 
        .QN(P2_sub_978_n167) );
  OR2X1 P2_sub_978_U166 ( .IN2(P2_sub_978_n164), .IN1(P2_sub_978_n169), 
        .Q(P2_sub_978_n168) );
  NAND2X0 P2_sub_978_U165 ( .IN1(P2_sub_978_n167), .IN2(P2_sub_978_n168), 
        .QN(P2_N3984) );
  INVX0 P2_sub_978_U164 ( .ZN(P2_sub_978_n145), .INP(P2_N3743) );
  NAND2X0 P2_sub_978_U163 ( .IN1(n7263), .IN2(P2_sub_978_n145), 
        .QN(P2_sub_978_n165) );
  OR2X1 P2_sub_978_U162 ( .IN2(n7263), .IN1(P2_sub_978_n145), 
        .Q(P2_sub_978_n166) );
  NAND2X0 P2_sub_978_U161 ( .IN1(P2_sub_978_n165), .IN2(P2_sub_978_n166), 
        .QN(P2_sub_978_n159) );
  NAND2X0 P2_sub_978_U160 ( .IN1(n7187), .IN2(P2_sub_978_n164), 
        .QN(P2_sub_978_n160) );
  OR2X1 P2_sub_978_U159 ( .IN2(n7187), .IN1(P2_sub_978_n164), 
        .Q(P2_sub_978_n162) );
  NAND2X0 P2_sub_978_U158 ( .IN1(P2_sub_978_n162), .IN2(P2_sub_978_n163), 
        .QN(P2_sub_978_n161) );
  NAND2X0 P2_sub_978_U157 ( .IN1(P2_sub_978_n160), .IN2(P2_sub_978_n161), 
        .QN(P2_sub_978_n146) );
  NAND2X0 P2_sub_978_U156 ( .IN1(P2_sub_978_n159), .IN2(P2_sub_978_n146), 
        .QN(P2_sub_978_n157) );
  OR2X1 P2_sub_978_U155 ( .IN2(P2_sub_978_n146), .IN1(P2_sub_978_n159), 
        .Q(P2_sub_978_n158) );
  NAND2X0 P2_sub_978_U154 ( .IN1(P2_sub_978_n157), .IN2(P2_sub_978_n158), 
        .QN(P2_N3985) );
  NAND2X0 P2_sub_978_U153 ( .IN1(P2_N5072), .IN2(P2_sub_978_n156), 
        .QN(P2_sub_978_n153) );
  NAND2X0 P2_sub_978_U152 ( .IN1(P2_N3725), .IN2(n7184), .QN(P2_sub_978_n154)
         );
  NAND2X0 P2_sub_978_U151 ( .IN1(P2_sub_978_n153), .IN2(P2_sub_978_n154), 
        .QN(P2_sub_978_n151) );
  NAND2X0 P2_sub_978_U150 ( .IN1(P2_sub_978_n151), .IN2(P2_sub_978_n152), 
        .QN(P2_sub_978_n149) );
  OR2X1 P2_sub_978_U149 ( .IN2(P2_sub_978_n152), .IN1(P2_sub_978_n151), 
        .Q(P2_sub_978_n150) );
  NAND2X0 P2_sub_978_U148 ( .IN1(P2_sub_978_n149), .IN2(P2_sub_978_n150), 
        .QN(P2_N3967) );
  INVX0 P2_sub_978_U147 ( .ZN(P2_sub_978_n135), .INP(P2_N3744) );
  NAND2X0 P2_sub_978_U146 ( .IN1(n7259), .IN2(P2_sub_978_n135), 
        .QN(P2_sub_978_n147) );
  OR2X1 P2_sub_978_U145 ( .IN2(n7259), .IN1(P2_sub_978_n135), 
        .Q(P2_sub_978_n148) );
  NAND2X0 P2_sub_978_U144 ( .IN1(P2_sub_978_n147), .IN2(P2_sub_978_n148), 
        .QN(P2_sub_978_n141) );
  NAND2X0 P2_sub_978_U143 ( .IN1(n7263), .IN2(P2_sub_978_n146), 
        .QN(P2_sub_978_n142) );
  OR2X1 P2_sub_978_U142 ( .IN2(n7263), .IN1(P2_sub_978_n146), 
        .Q(P2_sub_978_n144) );
  NAND2X0 P2_sub_978_U141 ( .IN1(P2_sub_978_n144), .IN2(P2_sub_978_n145), 
        .QN(P2_sub_978_n143) );
  NAND2X0 P2_sub_978_U140 ( .IN1(P2_sub_978_n142), .IN2(P2_sub_978_n143), 
        .QN(P2_sub_978_n136) );
  NAND2X0 P2_sub_978_U139 ( .IN1(P2_sub_978_n141), .IN2(P2_sub_978_n136), 
        .QN(P2_sub_978_n139) );
  OR2X1 P2_sub_978_U138 ( .IN2(P2_sub_978_n136), .IN1(P2_sub_978_n141), 
        .Q(P2_sub_978_n140) );
  NAND2X0 P2_sub_978_U137 ( .IN1(P2_sub_978_n139), .IN2(P2_sub_978_n140), 
        .QN(P2_N3986) );
  INVX0 P2_sub_978_U136 ( .ZN(P2_sub_978_n125), .INP(P2_N3745) );
  NAND2X0 P2_sub_978_U135 ( .IN1(n7252), .IN2(P2_sub_978_n125), 
        .QN(P2_sub_978_n137) );
  OR2X1 P2_sub_978_U134 ( .IN2(n7252), .IN1(P2_sub_978_n125), 
        .Q(P2_sub_978_n138) );
  NAND2X0 P2_sub_978_U133 ( .IN1(P2_sub_978_n137), .IN2(P2_sub_978_n138), 
        .QN(P2_sub_978_n131) );
  NAND2X0 P2_sub_978_U132 ( .IN1(n7259), .IN2(P2_sub_978_n136), 
        .QN(P2_sub_978_n132) );
  OR2X1 P2_sub_978_U131 ( .IN2(n7259), .IN1(P2_sub_978_n136), 
        .Q(P2_sub_978_n134) );
  NAND2X0 P2_sub_978_U130 ( .IN1(P2_sub_978_n134), .IN2(P2_sub_978_n135), 
        .QN(P2_sub_978_n133) );
  NAND2X0 P2_sub_978_U129 ( .IN1(P2_sub_978_n132), .IN2(P2_sub_978_n133), 
        .QN(P2_sub_978_n126) );
  NAND2X0 P2_sub_978_U128 ( .IN1(P2_sub_978_n131), .IN2(P2_sub_978_n126), 
        .QN(P2_sub_978_n129) );
  OR2X1 P2_sub_978_U127 ( .IN2(P2_sub_978_n126), .IN1(P2_sub_978_n131), 
        .Q(P2_sub_978_n130) );
  NAND2X0 P2_sub_978_U126 ( .IN1(P2_sub_978_n129), .IN2(P2_sub_978_n130), 
        .QN(P2_N3987) );
  INVX0 P2_sub_978_U125 ( .ZN(P2_sub_978_n115), .INP(P2_N3746) );
  NAND2X0 P2_sub_978_U124 ( .IN1(n7247), .IN2(P2_sub_978_n115), 
        .QN(P2_sub_978_n127) );
  OR2X1 P2_sub_978_U123 ( .IN2(n7247), .IN1(P2_sub_978_n115), 
        .Q(P2_sub_978_n128) );
  NAND2X0 P2_sub_978_U122 ( .IN1(P2_sub_978_n127), .IN2(P2_sub_978_n128), 
        .QN(P2_sub_978_n121) );
  NAND2X0 P2_sub_978_U121 ( .IN1(n7252), .IN2(P2_sub_978_n126), 
        .QN(P2_sub_978_n122) );
  OR2X1 P2_sub_978_U120 ( .IN2(n7252), .IN1(P2_sub_978_n126), 
        .Q(P2_sub_978_n124) );
  NAND2X0 P2_sub_978_U119 ( .IN1(P2_sub_978_n124), .IN2(P2_sub_978_n125), 
        .QN(P2_sub_978_n123) );
  NAND2X0 P2_sub_978_U118 ( .IN1(P2_sub_978_n122), .IN2(P2_sub_978_n123), 
        .QN(P2_sub_978_n116) );
  NAND2X0 P2_sub_978_U117 ( .IN1(P2_sub_978_n121), .IN2(P2_sub_978_n116), 
        .QN(P2_sub_978_n119) );
  OR2X1 P2_sub_978_U116 ( .IN2(P2_sub_978_n116), .IN1(P2_sub_978_n121), 
        .Q(P2_sub_978_n120) );
  NAND2X0 P2_sub_978_U115 ( .IN1(P2_sub_978_n119), .IN2(P2_sub_978_n120), 
        .QN(P2_N3988) );
  INVX0 P2_sub_978_U114 ( .ZN(P2_sub_978_n105), .INP(P2_N3747) );
  NAND2X0 P2_sub_978_U113 ( .IN1(n7242), .IN2(P2_sub_978_n105), 
        .QN(P2_sub_978_n117) );
  OR2X1 P2_sub_978_U112 ( .IN2(n7242), .IN1(P2_sub_978_n105), 
        .Q(P2_sub_978_n118) );
  NAND2X0 P2_sub_978_U111 ( .IN1(P2_sub_978_n117), .IN2(P2_sub_978_n118), 
        .QN(P2_sub_978_n111) );
  NAND2X0 P2_sub_978_U110 ( .IN1(n7247), .IN2(P2_sub_978_n116), 
        .QN(P2_sub_978_n112) );
  OR2X1 P2_sub_978_U109 ( .IN2(n7247), .IN1(P2_sub_978_n116), 
        .Q(P2_sub_978_n114) );
  NAND2X0 P2_sub_978_U108 ( .IN1(P2_sub_978_n114), .IN2(P2_sub_978_n115), 
        .QN(P2_sub_978_n113) );
  NAND2X0 P2_sub_978_U107 ( .IN1(P2_sub_978_n112), .IN2(P2_sub_978_n113), 
        .QN(P2_sub_978_n106) );
  NAND2X0 P2_sub_978_U106 ( .IN1(P2_sub_978_n111), .IN2(P2_sub_978_n106), 
        .QN(P2_sub_978_n109) );
  OR2X1 P2_sub_978_U105 ( .IN2(P2_sub_978_n106), .IN1(P2_sub_978_n111), 
        .Q(P2_sub_978_n110) );
  NAND2X0 P2_sub_978_U104 ( .IN1(P2_sub_978_n109), .IN2(P2_sub_978_n110), 
        .QN(P2_N3989) );
  INVX0 P2_sub_978_U103 ( .ZN(P2_sub_978_n95), .INP(P2_N3748) );
  NAND2X0 P2_sub_978_U102 ( .IN1(n7238), .IN2(P2_sub_978_n95), 
        .QN(P2_sub_978_n107) );
  OR2X1 P2_sub_978_U101 ( .IN2(n7238), .IN1(P2_sub_978_n95), 
        .Q(P2_sub_978_n108) );
  NAND2X0 P2_sub_978_U100 ( .IN1(P2_sub_978_n107), .IN2(P2_sub_978_n108), 
        .QN(P2_sub_978_n101) );
  NAND2X0 P2_sub_978_U99 ( .IN1(n7242), .IN2(P2_sub_978_n106), 
        .QN(P2_sub_978_n102) );
  OR2X1 P2_sub_978_U98 ( .IN2(n7242), .IN1(P2_sub_978_n106), 
        .Q(P2_sub_978_n104) );
  NAND2X0 P2_sub_978_U97 ( .IN1(P2_sub_978_n104), .IN2(P2_sub_978_n105), 
        .QN(P2_sub_978_n103) );
  NAND2X0 P2_sub_978_U96 ( .IN1(P2_sub_978_n102), .IN2(P2_sub_978_n103), 
        .QN(P2_sub_978_n96) );
  NAND2X0 P2_sub_978_U95 ( .IN1(P2_sub_978_n101), .IN2(P2_sub_978_n96), 
        .QN(P2_sub_978_n99) );
  OR2X1 P2_sub_978_U94 ( .IN2(P2_sub_978_n96), .IN1(P2_sub_978_n101), 
        .Q(P2_sub_978_n100) );
  NAND2X0 P2_sub_978_U93 ( .IN1(P2_sub_978_n99), .IN2(P2_sub_978_n100), 
        .QN(P2_N3990) );
  INVX0 P2_sub_978_U278 ( .ZN(P2_sub_978_n35), .INP(P2_N3729) );
  NAND2X0 P2_sub_978_U277 ( .IN1(P2_sub_978_n264), .IN2(P2_sub_978_n35), 
        .QN(P2_sub_978_n263) );
  NAND2X0 P2_sub_978_U276 ( .IN1(P2_sub_978_n262), .IN2(P2_sub_978_n263), 
        .QN(P2_sub_978_n25) );
  NAND2X0 P2_sub_978_U275 ( .IN1(P2_N5077), .IN2(P2_sub_978_n25), 
        .QN(P2_sub_978_n259) );
  OR2X1 P2_sub_978_U274 ( .IN2(P2_N5077), .IN1(P2_sub_978_n25), 
        .Q(P2_sub_978_n261) );
  INVX0 P2_sub_978_U273 ( .ZN(P2_sub_978_n28), .INP(P2_N3730) );
  NAND2X0 P2_sub_978_U272 ( .IN1(P2_sub_978_n261), .IN2(P2_sub_978_n28), 
        .QN(P2_sub_978_n260) );
  NAND2X0 P2_sub_978_U271 ( .IN1(P2_sub_978_n259), .IN2(P2_sub_978_n260), 
        .QN(P2_sub_978_n18) );
  NAND2X0 P2_sub_978_U270 ( .IN1(n7158), .IN2(P2_sub_978_n18), 
        .QN(P2_sub_978_n256) );
  OR2X1 P2_sub_978_U269 ( .IN2(n7158), .IN1(P2_sub_978_n18), 
        .Q(P2_sub_978_n258) );
  INVX0 P2_sub_978_U268 ( .ZN(P2_sub_978_n21), .INP(P2_N3731) );
  NAND2X0 P2_sub_978_U267 ( .IN1(P2_sub_978_n258), .IN2(P2_sub_978_n21), 
        .QN(P2_sub_978_n257) );
  NAND2X0 P2_sub_978_U266 ( .IN1(P2_sub_978_n256), .IN2(P2_sub_978_n257), 
        .QN(P2_sub_978_n11) );
  NAND2X0 P2_sub_978_U265 ( .IN1(n7154), .IN2(P2_sub_978_n11), 
        .QN(P2_sub_978_n253) );
  OR2X1 P2_sub_978_U264 ( .IN2(n7154), .IN1(P2_sub_978_n11), 
        .Q(P2_sub_978_n255) );
  INVX0 P2_sub_978_U263 ( .ZN(P2_sub_978_n14), .INP(P2_N3732) );
  NAND2X0 P2_sub_978_U262 ( .IN1(P2_sub_978_n255), .IN2(P2_sub_978_n14), 
        .QN(P2_sub_978_n254) );
  NAND2X0 P2_sub_978_U261 ( .IN1(P2_sub_978_n253), .IN2(P2_sub_978_n254), 
        .QN(P2_sub_978_n4) );
  NAND2X0 P2_sub_978_U260 ( .IN1(n7151), .IN2(P2_sub_978_n4), 
        .QN(P2_sub_978_n250) );
  OR2X1 P2_sub_978_U259 ( .IN2(n7151), .IN1(P2_sub_978_n4), 
        .Q(P2_sub_978_n252) );
  INVX0 P2_sub_978_U258 ( .ZN(P2_sub_978_n7), .INP(P2_N3733) );
  NAND2X0 P2_sub_978_U257 ( .IN1(P2_sub_978_n252), .IN2(P2_sub_978_n7), 
        .QN(P2_sub_978_n251) );
  NAND2X0 P2_sub_978_U256 ( .IN1(P2_sub_978_n250), .IN2(P2_sub_978_n251), 
        .QN(P2_sub_978_n244) );
  NAND2X0 P2_sub_978_U255 ( .IN1(P2_sub_978_n249), .IN2(P2_sub_978_n244), 
        .QN(P2_sub_978_n247) );
  OR2X1 P2_sub_978_U254 ( .IN2(P2_sub_978_n244), .IN1(P2_sub_978_n249), 
        .Q(P2_sub_978_n248) );
  NAND2X0 P2_sub_978_U253 ( .IN1(P2_sub_978_n247), .IN2(P2_sub_978_n248), 
        .QN(P2_N3976) );
  INVX0 P2_sub_978_U252 ( .ZN(P2_sub_978_n233), .INP(P2_N3735) );
  NAND2X0 P2_sub_978_U251 ( .IN1(n7216), .IN2(P2_sub_978_n233), 
        .QN(P2_sub_978_n245) );
  OR2X1 P2_sub_978_U250 ( .IN2(n7216), .IN1(P2_sub_978_n233), 
        .Q(P2_sub_978_n246) );
  NAND2X0 P2_sub_978_U249 ( .IN1(P2_sub_978_n245), .IN2(P2_sub_978_n246), 
        .QN(P2_sub_978_n239) );
  NAND2X0 P2_sub_978_U248 ( .IN1(P2_N5081), .IN2(P2_sub_978_n244), 
        .QN(P2_sub_978_n240) );
  OR2X1 P2_sub_978_U247 ( .IN2(P2_N5081), .IN1(P2_sub_978_n244), 
        .Q(P2_sub_978_n242) );
  NAND2X0 P2_sub_978_U246 ( .IN1(P2_sub_978_n242), .IN2(P2_sub_978_n243), 
        .QN(P2_sub_978_n241) );
  NAND2X0 P2_sub_978_U245 ( .IN1(P2_sub_978_n240), .IN2(P2_sub_978_n241), 
        .QN(P2_sub_978_n234) );
  NAND2X0 P2_sub_978_U244 ( .IN1(P2_sub_978_n239), .IN2(P2_sub_978_n234), 
        .QN(P2_sub_978_n237) );
  OR2X1 P2_sub_978_U243 ( .IN2(P2_sub_978_n234), .IN1(P2_sub_978_n239), 
        .Q(P2_sub_978_n238) );
  NAND2X0 P2_sub_978_U242 ( .IN1(P2_sub_978_n237), .IN2(P2_sub_978_n238), 
        .QN(P2_N3977) );
  INVX0 P2_sub_978_U241 ( .ZN(P2_sub_978_n223), .INP(P2_N3736) );
  NAND2X0 P2_sub_978_U240 ( .IN1(n7210), .IN2(P2_sub_978_n223), 
        .QN(P2_sub_978_n235) );
  OR2X1 P2_sub_978_U239 ( .IN2(n7210), .IN1(P2_sub_978_n223), 
        .Q(P2_sub_978_n236) );
  NAND2X0 P2_sub_978_U238 ( .IN1(P2_sub_978_n235), .IN2(P2_sub_978_n236), 
        .QN(P2_sub_978_n229) );
  NAND2X0 P2_sub_978_U237 ( .IN1(n7216), .IN2(P2_sub_978_n234), 
        .QN(P2_sub_978_n230) );
  OR2X1 P2_sub_978_U236 ( .IN2(n7216), .IN1(P2_sub_978_n234), 
        .Q(P2_sub_978_n232) );
  NAND2X0 P2_sub_978_U235 ( .IN1(P2_sub_978_n232), .IN2(P2_sub_978_n233), 
        .QN(P2_sub_978_n231) );
  NAND2X0 P2_sub_978_U234 ( .IN1(P2_sub_978_n230), .IN2(P2_sub_978_n231), 
        .QN(P2_sub_978_n224) );
  NAND2X0 P2_sub_978_U233 ( .IN1(P2_sub_978_n229), .IN2(P2_sub_978_n224), 
        .QN(P2_sub_978_n227) );
  OR2X1 P2_sub_978_U232 ( .IN2(P2_sub_978_n224), .IN1(P2_sub_978_n229), 
        .Q(P2_sub_978_n228) );
  NAND2X0 P2_sub_978_U231 ( .IN1(P2_sub_978_n227), .IN2(P2_sub_978_n228), 
        .QN(P2_N3978) );
  INVX0 P2_sub_978_U230 ( .ZN(P2_sub_978_n213), .INP(P2_N3737) );
  NAND2X0 P2_sub_978_U229 ( .IN1(n7209), .IN2(P2_sub_978_n213), 
        .QN(P2_sub_978_n225) );
  OR2X1 P2_sub_978_U228 ( .IN2(n7209), .IN1(P2_sub_978_n213), 
        .Q(P2_sub_978_n226) );
  NAND2X0 P2_sub_978_U227 ( .IN1(P2_sub_978_n225), .IN2(P2_sub_978_n226), 
        .QN(P2_sub_978_n219) );
  NAND2X0 P2_sub_978_U226 ( .IN1(n7210), .IN2(P2_sub_978_n224), 
        .QN(P2_sub_978_n220) );
  OR2X1 P2_sub_978_U225 ( .IN2(n7210), .IN1(P2_sub_978_n224), 
        .Q(P2_sub_978_n222) );
  NAND2X0 P2_sub_978_U224 ( .IN1(P2_sub_978_n222), .IN2(P2_sub_978_n223), 
        .QN(P2_sub_978_n221) );
  NAND2X0 P2_sub_978_U223 ( .IN1(P2_sub_978_n220), .IN2(P2_sub_978_n221), 
        .QN(P2_sub_978_n214) );
  NAND2X0 P2_sub_978_U222 ( .IN1(P2_sub_978_n219), .IN2(P2_sub_978_n214), 
        .QN(P2_sub_978_n217) );
  OR2X1 P2_sub_978_U221 ( .IN2(P2_sub_978_n214), .IN1(P2_sub_978_n219), 
        .Q(P2_sub_978_n218) );
  NAND2X0 P2_sub_978_U220 ( .IN1(P2_sub_978_n217), .IN2(P2_sub_978_n218), 
        .QN(P2_N3979) );
  INVX0 P2_sub_978_U219 ( .ZN(P2_sub_978_n203), .INP(P2_N3738) );
  NAND2X0 P2_sub_978_U218 ( .IN1(n7206), .IN2(P2_sub_978_n203), 
        .QN(P2_sub_978_n215) );
  OR2X1 P2_sub_978_U217 ( .IN2(n7206), .IN1(P2_sub_978_n203), 
        .Q(P2_sub_978_n216) );
  NAND2X0 P2_sub_978_U216 ( .IN1(P2_sub_978_n215), .IN2(P2_sub_978_n216), 
        .QN(P2_sub_978_n209) );
  NAND2X0 P2_sub_978_U215 ( .IN1(n7209), .IN2(P2_sub_978_n214), 
        .QN(P2_sub_978_n210) );
  OR2X1 P2_sub_978_U214 ( .IN2(n7209), .IN1(P2_sub_978_n214), 
        .Q(P2_sub_978_n212) );
  NAND2X0 P2_sub_978_U213 ( .IN1(P2_sub_978_n212), .IN2(P2_sub_978_n213), 
        .QN(P2_sub_978_n211) );
  NAND2X0 P2_sub_978_U212 ( .IN1(P2_sub_978_n210), .IN2(P2_sub_978_n211), 
        .QN(P2_sub_978_n204) );
  NAND2X0 P2_sub_978_U211 ( .IN1(P2_sub_978_n209), .IN2(P2_sub_978_n204), 
        .QN(P2_sub_978_n207) );
  OR2X1 P2_sub_978_U210 ( .IN2(P2_sub_978_n204), .IN1(P2_sub_978_n209), 
        .Q(P2_sub_978_n208) );
  NAND2X0 P2_sub_978_U209 ( .IN1(P2_sub_978_n207), .IN2(P2_sub_978_n208), 
        .QN(P2_N3980) );
  INVX0 P2_sub_978_U208 ( .ZN(P2_sub_978_n193), .INP(P2_N3739) );
  NAND2X0 P2_sub_978_U207 ( .IN1(n7202), .IN2(P2_sub_978_n193), 
        .QN(P2_sub_978_n205) );
  OR2X1 P2_sub_978_U206 ( .IN2(n7202), .IN1(P2_sub_978_n193), 
        .Q(P2_sub_978_n206) );
  NAND2X0 P2_sub_978_U205 ( .IN1(P2_sub_978_n205), .IN2(P2_sub_978_n206), 
        .QN(P2_sub_978_n199) );
  NAND2X0 P2_sub_978_U204 ( .IN1(n7206), .IN2(P2_sub_978_n204), 
        .QN(P2_sub_978_n200) );
  OR2X1 P2_sub_978_U203 ( .IN2(n7206), .IN1(P2_sub_978_n204), 
        .Q(P2_sub_978_n202) );
  NAND2X0 P2_sub_978_U202 ( .IN1(P2_sub_978_n202), .IN2(P2_sub_978_n203), 
        .QN(P2_sub_978_n201) );
  NAND2X0 P2_sub_978_U201 ( .IN1(P2_sub_978_n200), .IN2(P2_sub_978_n201), 
        .QN(P2_sub_978_n194) );
  NAND2X0 P2_sub_978_U200 ( .IN1(P2_sub_978_n199), .IN2(P2_sub_978_n194), 
        .QN(P2_sub_978_n197) );
  OR2X1 P2_sub_978_U199 ( .IN2(P2_sub_978_n194), .IN1(P2_sub_978_n199), 
        .Q(P2_sub_978_n198) );
  NAND2X0 P2_sub_978_U198 ( .IN1(P2_sub_978_n197), .IN2(P2_sub_978_n198), 
        .QN(P2_N3981) );
  INVX0 P2_sub_978_U197 ( .ZN(P2_sub_978_n183), .INP(P2_N3740) );
  NAND2X0 P2_sub_978_U196 ( .IN1(P2_N5087), .IN2(P2_sub_978_n183), 
        .QN(P2_sub_978_n195) );
  OR2X1 P2_sub_978_U195 ( .IN2(P2_N5087), .IN1(P2_sub_978_n183), 
        .Q(P2_sub_978_n196) );
  NAND2X0 P2_sub_978_U194 ( .IN1(P2_sub_978_n195), .IN2(P2_sub_978_n196), 
        .QN(P2_sub_978_n189) );
  NAND2X0 P2_sub_978_U193 ( .IN1(n7202), .IN2(P2_sub_978_n194), 
        .QN(P2_sub_978_n190) );
  OR2X1 P2_sub_978_U192 ( .IN2(n7202), .IN1(P2_sub_978_n194), 
        .Q(P2_sub_978_n192) );
  NAND2X0 P2_sub_978_U191 ( .IN1(P2_sub_978_n192), .IN2(P2_sub_978_n193), 
        .QN(P2_sub_978_n191) );
  NAND2X0 P2_sub_978_U190 ( .IN1(P2_sub_978_n190), .IN2(P2_sub_978_n191), 
        .QN(P2_sub_978_n184) );
  NAND2X0 P2_sub_978_U189 ( .IN1(P2_sub_978_n189), .IN2(P2_sub_978_n184), 
        .QN(P2_sub_978_n187) );
  OR2X1 P2_sub_978_U188 ( .IN2(P2_sub_978_n184), .IN1(P2_sub_978_n189), 
        .Q(P2_sub_978_n188) );
  NAND2X0 P2_sub_978_U187 ( .IN1(P2_sub_978_n187), .IN2(P2_sub_978_n188), 
        .QN(P2_N3982) );
  INVX0 P2_sub_978_U186 ( .ZN(P2_sub_978_n173), .INP(P2_N3741) );
  INVX0 P2_sub_978_U310 ( .ZN(P2_sub_978_n281), .INP(P2_N3724) );
  NOR2X0 P2_sub_978_U309 ( .QN(P2_sub_978_n277), .IN1(P2_sub_978_n281), 
        .IN2(n7035) );
  INVX0 P2_sub_978_U308 ( .ZN(P2_sub_978_n152), .INP(P2_sub_978_n277) );
  NAND2X0 P2_sub_978_U307 ( .IN1(n7035), .IN2(P2_sub_978_n281), 
        .QN(P2_sub_978_n280) );
  NAND2X0 P2_sub_978_U306 ( .IN1(P2_sub_978_n152), .IN2(P2_sub_978_n280), 
        .QN(P2_N3966) );
  INVX0 P2_sub_978_U305 ( .ZN(P2_sub_978_n243), .INP(P2_N3734) );
  NAND2X0 P2_sub_978_U304 ( .IN1(P2_N5081), .IN2(P2_sub_978_n243), 
        .QN(P2_sub_978_n278) );
  OR2X1 P2_sub_978_U303 ( .IN2(P2_N5081), .IN1(P2_sub_978_n243), 
        .Q(P2_sub_978_n279) );
  NAND2X0 P2_sub_978_U302 ( .IN1(P2_sub_978_n278), .IN2(P2_sub_978_n279), 
        .QN(P2_sub_978_n249) );
  NAND2X0 P2_sub_978_U301 ( .IN1(P2_N5072), .IN2(P2_sub_978_n152), 
        .QN(P2_sub_978_n274) );
  NAND2X0 P2_sub_978_U299 ( .IN1(P2_sub_978_n277), .IN2(n7184), 
        .QN(P2_sub_978_n276) );
  INVX0 P2_sub_978_U298 ( .ZN(P2_sub_978_n156), .INP(P2_N3725) );
  NAND2X0 P2_sub_978_U297 ( .IN1(P2_sub_978_n276), .IN2(P2_sub_978_n156), 
        .QN(P2_sub_978_n275) );
  NAND2X0 P2_sub_978_U296 ( .IN1(P2_sub_978_n274), .IN2(P2_sub_978_n275), 
        .QN(P2_sub_978_n53) );
  NAND2X0 P2_sub_978_U295 ( .IN1(n7181), .IN2(P2_sub_978_n53), 
        .QN(P2_sub_978_n271) );
  OR2X1 P2_sub_978_U294 ( .IN2(n7181), .IN1(P2_sub_978_n53), 
        .Q(P2_sub_978_n273) );
  INVX0 P2_sub_978_U293 ( .ZN(P2_sub_978_n56), .INP(P2_N3726) );
  NAND2X0 P2_sub_978_U292 ( .IN1(P2_sub_978_n273), .IN2(P2_sub_978_n56), 
        .QN(P2_sub_978_n272) );
  NAND2X0 P2_sub_978_U291 ( .IN1(P2_sub_978_n271), .IN2(P2_sub_978_n272), 
        .QN(P2_sub_978_n46) );
  NAND2X0 P2_sub_978_U290 ( .IN1(n7177), .IN2(P2_sub_978_n46), 
        .QN(P2_sub_978_n268) );
  OR2X1 P2_sub_978_U289 ( .IN2(n7177), .IN1(P2_sub_978_n46), 
        .Q(P2_sub_978_n270) );
  INVX0 P2_sub_978_U288 ( .ZN(P2_sub_978_n49), .INP(P2_N3727) );
  NAND2X0 P2_sub_978_U287 ( .IN1(P2_sub_978_n270), .IN2(P2_sub_978_n49), 
        .QN(P2_sub_978_n269) );
  NAND2X0 P2_sub_978_U286 ( .IN1(P2_sub_978_n268), .IN2(P2_sub_978_n269), 
        .QN(P2_sub_978_n39) );
  NAND2X0 P2_sub_978_U285 ( .IN1(n7173), .IN2(P2_sub_978_n39), 
        .QN(P2_sub_978_n265) );
  OR2X1 P2_sub_978_U284 ( .IN2(n7173), .IN1(P2_sub_978_n39), 
        .Q(P2_sub_978_n267) );
  INVX0 P2_sub_978_U283 ( .ZN(P2_sub_978_n42), .INP(P2_N3728) );
  NAND2X0 P2_sub_978_U282 ( .IN1(P2_sub_978_n267), .IN2(P2_sub_978_n42), 
        .QN(P2_sub_978_n266) );
  NAND2X0 P2_sub_978_U281 ( .IN1(P2_sub_978_n265), .IN2(P2_sub_978_n266), 
        .QN(P2_sub_978_n32) );
  NAND2X0 P2_sub_978_U280 ( .IN1(P2_N5076), .IN2(P2_sub_978_n32), 
        .QN(P2_sub_978_n262) );
  OR2X1 P2_sub_978_U279 ( .IN2(P2_N5076), .IN1(P2_sub_978_n32), 
        .Q(P2_sub_978_n264) );
  NOR2X0 P2_add_998_U29 ( .QN(P2_N4254), .IN1(P2_add_998_n29), 
        .IN2(P2_add_998_n30) );
  OR2X1 P2_add_998_U27 ( .IN2(P2_N4103), .IN1(n7164), .Q(P2_add_998_n26) );
  NAND2X0 P2_add_998_U26 ( .IN1(P2_N4103), .IN2(n7164), .QN(P2_add_998_n27) );
  NAND2X0 P2_add_998_U25 ( .IN1(P2_add_998_n26), .IN2(P2_add_998_n27), 
        .QN(P2_add_998_n25) );
  NOR2X0 P2_add_998_U24 ( .QN(P2_add_998_n22), .IN1(P2_add_998_n24), 
        .IN2(P2_add_998_n25) );
  AND2X1 P2_add_998_U23 ( .IN1(P2_add_998_n24), .IN2(P2_add_998_n25), 
        .Q(P2_add_998_n23) );
  NOR2X0 P2_add_998_U22 ( .QN(P2_N4255), .IN1(P2_add_998_n22), 
        .IN2(P2_add_998_n23) );
  OR2X1 P2_add_998_U20 ( .IN2(P2_N4104), .IN1(P2_add_998_n49), 
        .Q(P2_add_998_n19) );
  NAND2X0 P2_add_998_U19 ( .IN1(P2_N4104), .IN2(P2_add_998_n49), 
        .QN(P2_add_998_n20) );
  NAND2X0 P2_add_998_U18 ( .IN1(P2_add_998_n19), .IN2(P2_add_998_n20), 
        .QN(P2_add_998_n18) );
  NOR2X0 P2_add_998_U17 ( .QN(P2_add_998_n15), .IN1(P2_add_998_n17), 
        .IN2(P2_add_998_n18) );
  AND2X1 P2_add_998_U16 ( .IN1(P2_add_998_n17), .IN2(P2_add_998_n18), 
        .Q(P2_add_998_n16) );
  NOR2X0 P2_add_998_U15 ( .QN(P2_N4256), .IN1(P2_add_998_n15), 
        .IN2(P2_add_998_n16) );
  OR2X1 P2_add_998_U13 ( .IN2(P2_N4105), .IN1(n7153), .Q(P2_add_998_n12) );
  NAND2X0 P2_add_998_U12 ( .IN1(P2_N4105), .IN2(n7153), .QN(P2_add_998_n13) );
  NAND2X0 P2_add_998_U11 ( .IN1(P2_add_998_n12), .IN2(P2_add_998_n13), 
        .QN(P2_add_998_n11) );
  NOR2X0 P2_add_998_U10 ( .QN(P2_add_998_n8), .IN1(P2_add_998_n10), 
        .IN2(P2_add_998_n11) );
  AND2X1 P2_add_998_U9 ( .IN1(P2_add_998_n10), .IN2(P2_add_998_n11), 
        .Q(P2_add_998_n9) );
  NOR2X0 P2_add_998_U8 ( .QN(P2_N4257), .IN1(P2_add_998_n8), 
        .IN2(P2_add_998_n9) );
  OR2X1 P2_add_998_U6 ( .IN2(P2_N4106), .IN1(n7149), .Q(P2_add_998_n5) );
  NAND2X0 P2_add_998_U5 ( .IN1(P2_N4106), .IN2(n7149), .QN(P2_add_998_n6) );
  NAND2X0 P2_add_998_U4 ( .IN1(P2_add_998_n5), .IN2(P2_add_998_n6), 
        .QN(P2_add_998_n4) );
  NOR2X0 P2_add_998_U3 ( .QN(P2_add_998_n1), .IN1(P2_add_998_n3), 
        .IN2(P2_add_998_n4) );
  AND2X1 P2_add_998_U2 ( .IN1(P2_add_998_n3), .IN2(P2_add_998_n4), 
        .Q(P2_add_998_n2) );
  NOR2X0 P2_add_998_U1 ( .QN(P2_N4258), .IN1(P2_add_998_n1), 
        .IN2(P2_add_998_n2) );
  NAND2X0 P2_add_998_U122 ( .IN1(n7247), .IN2(P2_add_998_n117), 
        .QN(P2_add_998_n114) );
  OR2X1 P2_add_998_U121 ( .IN2(n7247), .IN1(P2_add_998_n117), 
        .Q(P2_add_998_n116) );
  NAND2X0 P2_add_998_U120 ( .IN1(P2_N4119), .IN2(P2_add_998_n116), 
        .QN(P2_add_998_n115) );
  NAND2X0 P2_add_998_U119 ( .IN1(P2_add_998_n114), .IN2(P2_add_998_n115), 
        .QN(P2_add_998_n107) );
  OR2X1 P2_add_998_U117 ( .IN2(P2_N4120), .IN1(n7243), .Q(P2_add_998_n111) );
  NAND2X0 P2_add_998_U116 ( .IN1(P2_N4120), .IN2(n7243), .QN(P2_add_998_n112)
         );
  NAND2X0 P2_add_998_U115 ( .IN1(P2_add_998_n111), .IN2(P2_add_998_n112), 
        .QN(P2_add_998_n110) );
  NOR2X0 P2_add_998_U114 ( .QN(P2_add_998_n108), .IN1(P2_add_998_n107), 
        .IN2(P2_add_998_n110) );
  AND2X1 P2_add_998_U113 ( .IN1(P2_add_998_n107), .IN2(P2_add_998_n110), 
        .Q(P2_add_998_n109) );
  NOR2X0 P2_add_998_U112 ( .QN(P2_N4272), .IN1(P2_add_998_n108), 
        .IN2(P2_add_998_n109) );
  NAND2X0 P2_add_998_U111 ( .IN1(n7242), .IN2(P2_add_998_n107), 
        .QN(P2_add_998_n104) );
  OR2X1 P2_add_998_U110 ( .IN2(n7242), .IN1(P2_add_998_n107), 
        .Q(P2_add_998_n106) );
  NAND2X0 P2_add_998_U109 ( .IN1(P2_N4120), .IN2(P2_add_998_n106), 
        .QN(P2_add_998_n105) );
  NAND2X0 P2_add_998_U108 ( .IN1(P2_add_998_n104), .IN2(P2_add_998_n105), 
        .QN(P2_add_998_n97) );
  OR2X1 P2_add_998_U106 ( .IN2(P2_N4121), .IN1(P2_add_998_n296), 
        .Q(P2_add_998_n101) );
  NAND2X0 P2_add_998_U105 ( .IN1(P2_N4121), .IN2(P2_add_998_n296), 
        .QN(P2_add_998_n102) );
  NAND2X0 P2_add_998_U104 ( .IN1(P2_add_998_n101), .IN2(P2_add_998_n102), 
        .QN(P2_add_998_n100) );
  NOR2X0 P2_add_998_U103 ( .QN(P2_add_998_n98), .IN1(P2_add_998_n97), 
        .IN2(P2_add_998_n100) );
  AND2X1 P2_add_998_U102 ( .IN1(P2_add_998_n97), .IN2(P2_add_998_n100), 
        .Q(P2_add_998_n99) );
  NOR2X0 P2_add_998_U101 ( .QN(P2_N4273), .IN1(P2_add_998_n98), 
        .IN2(P2_add_998_n99) );
  NAND2X0 P2_add_998_U100 ( .IN1(n7238), .IN2(P2_add_998_n97), 
        .QN(P2_add_998_n94) );
  OR2X1 P2_add_998_U99 ( .IN2(n7238), .IN1(P2_add_998_n97), .Q(P2_add_998_n96)
         );
  NAND2X0 P2_add_998_U98 ( .IN1(P2_N4121), .IN2(P2_add_998_n96), 
        .QN(P2_add_998_n95) );
  NAND2X0 P2_add_998_U97 ( .IN1(P2_add_998_n94), .IN2(P2_add_998_n95), 
        .QN(P2_add_998_n87) );
  OR2X1 P2_add_998_U95 ( .IN2(P2_N4122), .IN1(n7234), .Q(P2_add_998_n91) );
  NAND2X0 P2_add_998_U94 ( .IN1(P2_N4122), .IN2(n7234), .QN(P2_add_998_n92) );
  NAND2X0 P2_add_998_U93 ( .IN1(P2_add_998_n91), .IN2(P2_add_998_n92), 
        .QN(P2_add_998_n90) );
  NOR2X0 P2_add_998_U92 ( .QN(P2_add_998_n88), .IN1(P2_add_998_n87), 
        .IN2(P2_add_998_n90) );
  AND2X1 P2_add_998_U91 ( .IN1(P2_add_998_n87), .IN2(P2_add_998_n90), 
        .Q(P2_add_998_n89) );
  NOR2X0 P2_add_998_U90 ( .QN(P2_N4274), .IN1(P2_add_998_n88), 
        .IN2(P2_add_998_n89) );
  NAND2X0 P2_add_998_U89 ( .IN1(n7237), .IN2(P2_add_998_n87), 
        .QN(P2_add_998_n84) );
  OR2X1 P2_add_998_U88 ( .IN2(n7237), .IN1(P2_add_998_n87), .Q(P2_add_998_n86)
         );
  NAND2X0 P2_add_998_U87 ( .IN1(P2_N4122), .IN2(P2_add_998_n86), 
        .QN(P2_add_998_n85) );
  NAND2X0 P2_add_998_U86 ( .IN1(P2_add_998_n84), .IN2(P2_add_998_n85), 
        .QN(P2_add_998_n77) );
  OR2X1 P2_add_998_U84 ( .IN2(P2_N4123), .IN1(n7229), .Q(P2_add_998_n81) );
  NAND2X0 P2_add_998_U83 ( .IN1(P2_N4123), .IN2(n7229), .QN(P2_add_998_n82) );
  NAND2X0 P2_add_998_U82 ( .IN1(P2_add_998_n81), .IN2(P2_add_998_n82), 
        .QN(P2_add_998_n80) );
  NOR2X0 P2_add_998_U81 ( .QN(P2_add_998_n78), .IN1(P2_add_998_n77), 
        .IN2(P2_add_998_n80) );
  AND2X1 P2_add_998_U80 ( .IN1(P2_add_998_n77), .IN2(P2_add_998_n80), 
        .Q(P2_add_998_n79) );
  NOR2X0 P2_add_998_U79 ( .QN(P2_N4275), .IN1(P2_add_998_n78), 
        .IN2(P2_add_998_n79) );
  NAND2X0 P2_add_998_U78 ( .IN1(n7231), .IN2(P2_add_998_n77), 
        .QN(P2_add_998_n74) );
  OR2X1 P2_add_998_U77 ( .IN2(n7231), .IN1(P2_add_998_n77), .Q(P2_add_998_n76)
         );
  NAND2X0 P2_add_998_U76 ( .IN1(P2_N4123), .IN2(P2_add_998_n76), 
        .QN(P2_add_998_n75) );
  NAND2X0 P2_add_998_U75 ( .IN1(P2_add_998_n74), .IN2(P2_add_998_n75), 
        .QN(P2_add_998_n64) );
  OR2X1 P2_add_998_U73 ( .IN2(P2_N4124), .IN1(n7224), .Q(P2_add_998_n71) );
  NAND2X0 P2_add_998_U72 ( .IN1(P2_N4124), .IN2(n7224), .QN(P2_add_998_n72) );
  NAND2X0 P2_add_998_U71 ( .IN1(P2_add_998_n71), .IN2(P2_add_998_n72), 
        .QN(P2_add_998_n70) );
  NOR2X0 P2_add_998_U70 ( .QN(P2_add_998_n68), .IN1(P2_add_998_n64), 
        .IN2(P2_add_998_n70) );
  AND2X1 P2_add_998_U69 ( .IN1(P2_add_998_n64), .IN2(P2_add_998_n70), 
        .Q(P2_add_998_n69) );
  NOR2X0 P2_add_998_U68 ( .QN(P2_N4276), .IN1(P2_add_998_n68), 
        .IN2(P2_add_998_n69) );
  OR2X1 P2_add_998_U66 ( .IN2(P2_N4125), .IN1(n7222), .Q(P2_add_998_n65) );
  NAND2X0 P2_add_998_U65 ( .IN1(P2_N4125), .IN2(n7222), .QN(P2_add_998_n66) );
  NAND2X0 P2_add_998_U64 ( .IN1(P2_add_998_n65), .IN2(P2_add_998_n66), 
        .QN(P2_add_998_n60) );
  NAND2X0 P2_add_998_U63 ( .IN1(P2_N5098), .IN2(P2_add_998_n64), 
        .QN(P2_add_998_n61) );
  OR2X1 P2_add_998_U62 ( .IN2(P2_N5098), .IN1(P2_add_998_n64), 
        .Q(P2_add_998_n63) );
  NAND2X0 P2_add_998_U61 ( .IN1(P2_N4124), .IN2(P2_add_998_n63), 
        .QN(P2_add_998_n62) );
  NAND2X0 P2_add_998_U60 ( .IN1(P2_add_998_n61), .IN2(P2_add_998_n62), 
        .QN(P2_add_998_n59) );
  NOR2X0 P2_add_998_U59 ( .QN(P2_add_998_n57), .IN1(P2_add_998_n60), 
        .IN2(P2_add_998_n59) );
  AND2X1 P2_add_998_U58 ( .IN1(P2_add_998_n59), .IN2(P2_add_998_n60), 
        .Q(P2_add_998_n58) );
  NOR2X0 P2_add_998_U57 ( .QN(P2_N4277), .IN1(P2_add_998_n57), 
        .IN2(P2_add_998_n58) );
  OR2X1 P2_add_998_U55 ( .IN2(P2_N4099), .IN1(n7182), .Q(P2_add_998_n54) );
  NAND2X0 P2_add_998_U54 ( .IN1(P2_N4099), .IN2(n7182), .QN(P2_add_998_n55) );
  NAND2X0 P2_add_998_U53 ( .IN1(P2_add_998_n54), .IN2(P2_add_998_n55), 
        .QN(P2_add_998_n53) );
  NOR2X0 P2_add_998_U52 ( .QN(P2_add_998_n50), .IN1(P2_add_998_n52), 
        .IN2(P2_add_998_n53) );
  AND2X1 P2_add_998_U51 ( .IN1(P2_add_998_n52), .IN2(P2_add_998_n53), 
        .Q(P2_add_998_n51) );
  NOR2X0 P2_add_998_U50 ( .QN(P2_N4251), .IN1(P2_add_998_n50), 
        .IN2(P2_add_998_n51) );
  OR2X1 P2_add_998_U48 ( .IN2(P2_N4100), .IN1(n7178), .Q(P2_add_998_n47) );
  NAND2X0 P2_add_998_U47 ( .IN1(P2_N4100), .IN2(n7178), .QN(P2_add_998_n48) );
  NAND2X0 P2_add_998_U46 ( .IN1(P2_add_998_n47), .IN2(P2_add_998_n48), 
        .QN(P2_add_998_n46) );
  NOR2X0 P2_add_998_U45 ( .QN(P2_add_998_n43), .IN1(P2_add_998_n45), 
        .IN2(P2_add_998_n46) );
  AND2X1 P2_add_998_U44 ( .IN1(P2_add_998_n45), .IN2(P2_add_998_n46), 
        .Q(P2_add_998_n44) );
  NOR2X0 P2_add_998_U43 ( .QN(P2_N4252), .IN1(P2_add_998_n43), 
        .IN2(P2_add_998_n44) );
  OR2X1 P2_add_998_U41 ( .IN2(P2_N4101), .IN1(n7174), .Q(P2_add_998_n40) );
  NAND2X0 P2_add_998_U40 ( .IN1(P2_N4101), .IN2(n7174), .QN(P2_add_998_n41) );
  NAND2X0 P2_add_998_U39 ( .IN1(P2_add_998_n40), .IN2(P2_add_998_n41), 
        .QN(P2_add_998_n39) );
  NOR2X0 P2_add_998_U38 ( .QN(P2_add_998_n36), .IN1(P2_add_998_n38), 
        .IN2(P2_add_998_n39) );
  AND2X1 P2_add_998_U37 ( .IN1(P2_add_998_n38), .IN2(P2_add_998_n39), 
        .Q(P2_add_998_n37) );
  NOR2X0 P2_add_998_U36 ( .QN(P2_N4253), .IN1(P2_add_998_n36), 
        .IN2(P2_add_998_n37) );
  OR2X1 P2_add_998_U34 ( .IN2(P2_N4102), .IN1(n7166), .Q(P2_add_998_n33) );
  NAND2X0 P2_add_998_U33 ( .IN1(P2_N4102), .IN2(n7166), .QN(P2_add_998_n34) );
  NAND2X0 P2_add_998_U32 ( .IN1(P2_add_998_n33), .IN2(P2_add_998_n34), 
        .QN(P2_add_998_n32) );
  NOR2X0 P2_add_998_U31 ( .QN(P2_add_998_n29), .IN1(P2_add_998_n31), 
        .IN2(P2_add_998_n32) );
  AND2X1 P2_add_998_U30 ( .IN1(P2_add_998_n31), .IN2(P2_add_998_n32), 
        .Q(P2_add_998_n30) );
  OR2X1 P2_add_998_U215 ( .IN2(n7206), .IN1(P2_add_998_n204), 
        .Q(P2_add_998_n203) );
  NAND2X0 P2_add_998_U214 ( .IN1(P2_N4111), .IN2(P2_add_998_n203), 
        .QN(P2_add_998_n202) );
  NAND2X0 P2_add_998_U213 ( .IN1(P2_add_998_n201), .IN2(P2_add_998_n202), 
        .QN(P2_add_998_n194) );
  OR2X1 P2_add_998_U211 ( .IN2(P2_N4112), .IN1(n7201), .Q(P2_add_998_n198) );
  NAND2X0 P2_add_998_U210 ( .IN1(P2_N4112), .IN2(n7201), .QN(P2_add_998_n199)
         );
  NAND2X0 P2_add_998_U209 ( .IN1(P2_add_998_n198), .IN2(P2_add_998_n199), 
        .QN(P2_add_998_n197) );
  NOR2X0 P2_add_998_U208 ( .QN(P2_add_998_n195), .IN1(P2_add_998_n194), 
        .IN2(P2_add_998_n197) );
  AND2X1 P2_add_998_U207 ( .IN1(P2_add_998_n194), .IN2(P2_add_998_n197), 
        .Q(P2_add_998_n196) );
  NOR2X0 P2_add_998_U206 ( .QN(P2_N4264), .IN1(P2_add_998_n195), 
        .IN2(P2_add_998_n196) );
  NAND2X0 P2_add_998_U205 ( .IN1(n7202), .IN2(P2_add_998_n194), 
        .QN(P2_add_998_n191) );
  OR2X1 P2_add_998_U204 ( .IN2(n7202), .IN1(P2_add_998_n194), 
        .Q(P2_add_998_n193) );
  NAND2X0 P2_add_998_U203 ( .IN1(P2_N4112), .IN2(P2_add_998_n193), 
        .QN(P2_add_998_n192) );
  NAND2X0 P2_add_998_U202 ( .IN1(P2_add_998_n191), .IN2(P2_add_998_n192), 
        .QN(P2_add_998_n184) );
  OR2X1 P2_add_998_U200 ( .IN2(P2_N4113), .IN1(n7197), .Q(P2_add_998_n188) );
  NAND2X0 P2_add_998_U199 ( .IN1(P2_N4113), .IN2(n7197), .QN(P2_add_998_n189)
         );
  NAND2X0 P2_add_998_U198 ( .IN1(P2_add_998_n188), .IN2(P2_add_998_n189), 
        .QN(P2_add_998_n187) );
  NOR2X0 P2_add_998_U197 ( .QN(P2_add_998_n185), .IN1(P2_add_998_n184), 
        .IN2(P2_add_998_n187) );
  AND2X1 P2_add_998_U196 ( .IN1(P2_add_998_n184), .IN2(P2_add_998_n187), 
        .Q(P2_add_998_n186) );
  NOR2X0 P2_add_998_U195 ( .QN(P2_N4265), .IN1(P2_add_998_n185), 
        .IN2(P2_add_998_n186) );
  NAND2X0 P2_add_998_U194 ( .IN1(n7198), .IN2(P2_add_998_n184), 
        .QN(P2_add_998_n181) );
  OR2X1 P2_add_998_U193 ( .IN2(n7198), .IN1(P2_add_998_n184), 
        .Q(P2_add_998_n183) );
  NAND2X0 P2_add_998_U192 ( .IN1(P2_N4113), .IN2(P2_add_998_n183), 
        .QN(P2_add_998_n182) );
  NAND2X0 P2_add_998_U191 ( .IN1(P2_add_998_n181), .IN2(P2_add_998_n182), 
        .QN(P2_add_998_n174) );
  OR2X1 P2_add_998_U189 ( .IN2(P2_N4114), .IN1(n7195), .Q(P2_add_998_n178) );
  NAND2X0 P2_add_998_U188 ( .IN1(P2_N4114), .IN2(n7195), .QN(P2_add_998_n179)
         );
  NAND2X0 P2_add_998_U187 ( .IN1(P2_add_998_n178), .IN2(P2_add_998_n179), 
        .QN(P2_add_998_n177) );
  NOR2X0 P2_add_998_U186 ( .QN(P2_add_998_n175), .IN1(P2_add_998_n174), 
        .IN2(P2_add_998_n177) );
  AND2X1 P2_add_998_U185 ( .IN1(P2_add_998_n174), .IN2(P2_add_998_n177), 
        .Q(P2_add_998_n176) );
  NOR2X0 P2_add_998_U184 ( .QN(P2_N4266), .IN1(P2_add_998_n175), 
        .IN2(P2_add_998_n176) );
  NAND2X0 P2_add_998_U183 ( .IN1(n7194), .IN2(P2_add_998_n174), 
        .QN(P2_add_998_n171) );
  OR2X1 P2_add_998_U182 ( .IN2(n7194), .IN1(P2_add_998_n174), 
        .Q(P2_add_998_n173) );
  NAND2X0 P2_add_998_U181 ( .IN1(P2_N4114), .IN2(P2_add_998_n173), 
        .QN(P2_add_998_n172) );
  NAND2X0 P2_add_998_U180 ( .IN1(P2_add_998_n171), .IN2(P2_add_998_n172), 
        .QN(P2_add_998_n164) );
  OR2X1 P2_add_998_U178 ( .IN2(P2_N4115), .IN1(n7188), .Q(P2_add_998_n168) );
  NAND2X0 P2_add_998_U177 ( .IN1(P2_N4115), .IN2(n7188), .QN(P2_add_998_n169)
         );
  NAND2X0 P2_add_998_U176 ( .IN1(P2_add_998_n168), .IN2(P2_add_998_n169), 
        .QN(P2_add_998_n167) );
  NOR2X0 P2_add_998_U175 ( .QN(P2_add_998_n165), .IN1(P2_add_998_n164), 
        .IN2(P2_add_998_n167) );
  AND2X1 P2_add_998_U174 ( .IN1(P2_add_998_n164), .IN2(P2_add_998_n167), 
        .Q(P2_add_998_n166) );
  NOR2X0 P2_add_998_U173 ( .QN(P2_N4267), .IN1(P2_add_998_n165), 
        .IN2(P2_add_998_n166) );
  NAND2X0 P2_add_998_U172 ( .IN1(n7187), .IN2(P2_add_998_n164), 
        .QN(P2_add_998_n161) );
  OR2X1 P2_add_998_U171 ( .IN2(n7187), .IN1(P2_add_998_n164), 
        .Q(P2_add_998_n163) );
  NAND2X0 P2_add_998_U170 ( .IN1(P2_N4115), .IN2(P2_add_998_n163), 
        .QN(P2_add_998_n162) );
  NAND2X0 P2_add_998_U169 ( .IN1(P2_add_998_n161), .IN2(P2_add_998_n162), 
        .QN(P2_add_998_n147) );
  OR2X1 P2_add_998_U167 ( .IN2(P2_N4116), .IN1(n7264), .Q(P2_add_998_n158) );
  NAND2X0 P2_add_998_U166 ( .IN1(P2_N4116), .IN2(n7264), .QN(P2_add_998_n159)
         );
  NAND2X0 P2_add_998_U165 ( .IN1(P2_add_998_n158), .IN2(P2_add_998_n159), 
        .QN(P2_add_998_n157) );
  NOR2X0 P2_add_998_U164 ( .QN(P2_add_998_n155), .IN1(P2_add_998_n147), 
        .IN2(P2_add_998_n157) );
  AND2X1 P2_add_998_U163 ( .IN1(P2_add_998_n147), .IN2(P2_add_998_n157), 
        .Q(P2_add_998_n156) );
  NOR2X0 P2_add_998_U162 ( .QN(P2_N4268), .IN1(P2_add_998_n155), 
        .IN2(P2_add_998_n156) );
  OR2X1 P2_add_998_U161 ( .IN2(P2_N4098), .IN1(n7186), .Q(P2_add_998_n152) );
  NAND2X0 P2_add_998_U160 ( .IN1(P2_N4098), .IN2(n7186), .QN(P2_add_998_n153)
         );
  NAND2X0 P2_add_998_U159 ( .IN1(P2_add_998_n152), .IN2(P2_add_998_n153), 
        .QN(P2_add_998_n150) );
  NAND2X0 P2_add_998_U158 ( .IN1(P2_add_998_n150), .IN2(P2_add_998_n151), 
        .QN(P2_add_998_n148) );
  OR2X1 P2_add_998_U157 ( .IN2(P2_add_998_n151), .IN1(P2_add_998_n150), 
        .Q(P2_add_998_n149) );
  NAND2X0 P2_add_998_U156 ( .IN1(P2_add_998_n148), .IN2(P2_add_998_n149), 
        .QN(P2_N4250) );
  NAND2X0 P2_add_998_U155 ( .IN1(n7263), .IN2(P2_add_998_n147), 
        .QN(P2_add_998_n144) );
  OR2X1 P2_add_998_U154 ( .IN2(n7263), .IN1(P2_add_998_n147), 
        .Q(P2_add_998_n146) );
  NAND2X0 P2_add_998_U153 ( .IN1(P2_N4116), .IN2(P2_add_998_n146), 
        .QN(P2_add_998_n145) );
  NAND2X0 P2_add_998_U152 ( .IN1(P2_add_998_n144), .IN2(P2_add_998_n145), 
        .QN(P2_add_998_n137) );
  OR2X1 P2_add_998_U150 ( .IN2(P2_N4117), .IN1(n7260), .Q(P2_add_998_n141) );
  NAND2X0 P2_add_998_U149 ( .IN1(P2_N4117), .IN2(n7260), .QN(P2_add_998_n142)
         );
  NAND2X0 P2_add_998_U148 ( .IN1(P2_add_998_n141), .IN2(P2_add_998_n142), 
        .QN(P2_add_998_n140) );
  NOR2X0 P2_add_998_U147 ( .QN(P2_add_998_n138), .IN1(P2_add_998_n137), 
        .IN2(P2_add_998_n140) );
  AND2X1 P2_add_998_U146 ( .IN1(P2_add_998_n137), .IN2(P2_add_998_n140), 
        .Q(P2_add_998_n139) );
  NOR2X0 P2_add_998_U145 ( .QN(P2_N4269), .IN1(P2_add_998_n138), 
        .IN2(P2_add_998_n139) );
  NAND2X0 P2_add_998_U144 ( .IN1(n7259), .IN2(P2_add_998_n137), 
        .QN(P2_add_998_n134) );
  OR2X1 P2_add_998_U143 ( .IN2(n7259), .IN1(P2_add_998_n137), 
        .Q(P2_add_998_n136) );
  NAND2X0 P2_add_998_U142 ( .IN1(P2_N4117), .IN2(P2_add_998_n136), 
        .QN(P2_add_998_n135) );
  NAND2X0 P2_add_998_U141 ( .IN1(P2_add_998_n134), .IN2(P2_add_998_n135), 
        .QN(P2_add_998_n127) );
  OR2X1 P2_add_998_U139 ( .IN2(P2_N4118), .IN1(n7253), .Q(P2_add_998_n131) );
  NAND2X0 P2_add_998_U138 ( .IN1(P2_N4118), .IN2(n7253), .QN(P2_add_998_n132)
         );
  NAND2X0 P2_add_998_U137 ( .IN1(P2_add_998_n131), .IN2(P2_add_998_n132), 
        .QN(P2_add_998_n130) );
  NOR2X0 P2_add_998_U136 ( .QN(P2_add_998_n128), .IN1(P2_add_998_n127), 
        .IN2(P2_add_998_n130) );
  AND2X1 P2_add_998_U135 ( .IN1(P2_add_998_n127), .IN2(P2_add_998_n130), 
        .Q(P2_add_998_n129) );
  NOR2X0 P2_add_998_U134 ( .QN(P2_N4270), .IN1(P2_add_998_n128), 
        .IN2(P2_add_998_n129) );
  NAND2X0 P2_add_998_U133 ( .IN1(n7252), .IN2(P2_add_998_n127), 
        .QN(P2_add_998_n124) );
  OR2X1 P2_add_998_U132 ( .IN2(n7252), .IN1(P2_add_998_n127), 
        .Q(P2_add_998_n126) );
  NAND2X0 P2_add_998_U131 ( .IN1(P2_N4118), .IN2(P2_add_998_n126), 
        .QN(P2_add_998_n125) );
  NAND2X0 P2_add_998_U130 ( .IN1(P2_add_998_n124), .IN2(P2_add_998_n125), 
        .QN(P2_add_998_n117) );
  OR2X1 P2_add_998_U128 ( .IN2(P2_N4119), .IN1(n7248), .Q(P2_add_998_n121) );
  NAND2X0 P2_add_998_U127 ( .IN1(P2_N4119), .IN2(n7248), .QN(P2_add_998_n122)
         );
  NAND2X0 P2_add_998_U126 ( .IN1(P2_add_998_n121), .IN2(P2_add_998_n122), 
        .QN(P2_add_998_n120) );
  NOR2X0 P2_add_998_U125 ( .QN(P2_add_998_n118), .IN1(P2_add_998_n117), 
        .IN2(P2_add_998_n120) );
  AND2X1 P2_add_998_U124 ( .IN1(P2_add_998_n117), .IN2(P2_add_998_n120), 
        .Q(P2_add_998_n119) );
  NOR2X0 P2_add_998_U123 ( .QN(P2_N4271), .IN1(P2_add_998_n118), 
        .IN2(P2_add_998_n119) );
  OR2X1 P2_add_998_U308 ( .IN2(P2_N4097), .IN1(n2919), .Q(P2_add_998_n278) );
  NAND2X0 P2_add_998_U307 ( .IN1(P2_N4097), .IN2(n2919), .QN(P2_add_998_n279)
         );
  NAND2X0 P2_add_998_U306 ( .IN1(P2_add_998_n278), .IN2(P2_add_998_n279), 
        .QN(P2_N4249) );
  NAND2X0 P2_add_998_U304 ( .IN1(P2_N4097), .IN2(n7035), .QN(P2_add_998_n151)
         );
  OR2X1 P2_add_998_U303 ( .IN2(P2_add_998_n151), .IN1(n7186), 
        .Q(P2_add_998_n275) );
  NAND2X0 P2_add_998_U302 ( .IN1(n7186), .IN2(P2_add_998_n151), 
        .QN(P2_add_998_n277) );
  NAND2X0 P2_add_998_U301 ( .IN1(P2_N4098), .IN2(P2_add_998_n277), 
        .QN(P2_add_998_n276) );
  NAND2X0 P2_add_998_U300 ( .IN1(P2_add_998_n275), .IN2(P2_add_998_n276), 
        .QN(P2_add_998_n52) );
  NAND2X0 P2_add_998_U299 ( .IN1(n7181), .IN2(P2_add_998_n52), 
        .QN(P2_add_998_n272) );
  OR2X1 P2_add_998_U298 ( .IN2(n7181), .IN1(P2_add_998_n52), 
        .Q(P2_add_998_n274) );
  NAND2X0 P2_add_998_U297 ( .IN1(P2_N4099), .IN2(P2_add_998_n274), 
        .QN(P2_add_998_n273) );
  NAND2X0 P2_add_998_U296 ( .IN1(P2_add_998_n272), .IN2(P2_add_998_n273), 
        .QN(P2_add_998_n45) );
  NAND2X0 P2_add_998_U295 ( .IN1(n7177), .IN2(P2_add_998_n45), 
        .QN(P2_add_998_n269) );
  OR2X1 P2_add_998_U294 ( .IN2(n7177), .IN1(P2_add_998_n45), 
        .Q(P2_add_998_n271) );
  NAND2X0 P2_add_998_U293 ( .IN1(P2_N4100), .IN2(P2_add_998_n271), 
        .QN(P2_add_998_n270) );
  NAND2X0 P2_add_998_U292 ( .IN1(P2_add_998_n269), .IN2(P2_add_998_n270), 
        .QN(P2_add_998_n38) );
  NAND2X0 P2_add_998_U291 ( .IN1(n7173), .IN2(P2_add_998_n38), 
        .QN(P2_add_998_n266) );
  OR2X1 P2_add_998_U290 ( .IN2(n7173), .IN1(P2_add_998_n38), 
        .Q(P2_add_998_n268) );
  NAND2X0 P2_add_998_U289 ( .IN1(P2_N4101), .IN2(P2_add_998_n268), 
        .QN(P2_add_998_n267) );
  NAND2X0 P2_add_998_U288 ( .IN1(P2_add_998_n266), .IN2(P2_add_998_n267), 
        .QN(P2_add_998_n31) );
  NAND2X0 P2_add_998_U287 ( .IN1(n7165), .IN2(P2_add_998_n31), 
        .QN(P2_add_998_n263) );
  OR2X1 P2_add_998_U286 ( .IN2(n7165), .IN1(P2_add_998_n31), 
        .Q(P2_add_998_n265) );
  NAND2X0 P2_add_998_U285 ( .IN1(P2_N4102), .IN2(P2_add_998_n265), 
        .QN(P2_add_998_n264) );
  NAND2X0 P2_add_998_U284 ( .IN1(P2_add_998_n263), .IN2(P2_add_998_n264), 
        .QN(P2_add_998_n24) );
  NAND2X0 P2_add_998_U283 ( .IN1(P2_N5077), .IN2(P2_add_998_n24), 
        .QN(P2_add_998_n260) );
  OR2X1 P2_add_998_U282 ( .IN2(P2_N5077), .IN1(P2_add_998_n24), 
        .Q(P2_add_998_n262) );
  NAND2X0 P2_add_998_U281 ( .IN1(P2_N4103), .IN2(P2_add_998_n262), 
        .QN(P2_add_998_n261) );
  NAND2X0 P2_add_998_U280 ( .IN1(P2_add_998_n260), .IN2(P2_add_998_n261), 
        .QN(P2_add_998_n17) );
  NAND2X0 P2_add_998_U279 ( .IN1(n7158), .IN2(P2_add_998_n17), 
        .QN(P2_add_998_n257) );
  OR2X1 P2_add_998_U278 ( .IN2(n7158), .IN1(P2_add_998_n17), 
        .Q(P2_add_998_n259) );
  NAND2X0 P2_add_998_U277 ( .IN1(P2_N4104), .IN2(P2_add_998_n259), 
        .QN(P2_add_998_n258) );
  NAND2X0 P2_add_998_U276 ( .IN1(P2_add_998_n257), .IN2(P2_add_998_n258), 
        .QN(P2_add_998_n10) );
  NAND2X0 P2_add_998_U275 ( .IN1(n7154), .IN2(P2_add_998_n10), 
        .QN(P2_add_998_n254) );
  OR2X1 P2_add_998_U274 ( .IN2(n7154), .IN1(P2_add_998_n10), 
        .Q(P2_add_998_n256) );
  NAND2X0 P2_add_998_U273 ( .IN1(P2_N4105), .IN2(P2_add_998_n256), 
        .QN(P2_add_998_n255) );
  NAND2X0 P2_add_998_U272 ( .IN1(P2_add_998_n254), .IN2(P2_add_998_n255), 
        .QN(P2_add_998_n3) );
  NAND2X0 P2_add_998_U271 ( .IN1(n7151), .IN2(P2_add_998_n3), 
        .QN(P2_add_998_n251) );
  OR2X1 P2_add_998_U270 ( .IN2(n7151), .IN1(P2_add_998_n3), 
        .Q(P2_add_998_n253) );
  NAND2X0 P2_add_998_U269 ( .IN1(P2_N4106), .IN2(P2_add_998_n253), 
        .QN(P2_add_998_n252) );
  NAND2X0 P2_add_998_U268 ( .IN1(P2_add_998_n251), .IN2(P2_add_998_n252), 
        .QN(P2_add_998_n244) );
  OR2X1 P2_add_998_U266 ( .IN2(P2_N4107), .IN1(n7219), .Q(P2_add_998_n248) );
  NAND2X0 P2_add_998_U265 ( .IN1(P2_N4107), .IN2(n7219), .QN(P2_add_998_n249)
         );
  NAND2X0 P2_add_998_U264 ( .IN1(P2_add_998_n248), .IN2(P2_add_998_n249), 
        .QN(P2_add_998_n247) );
  NOR2X0 P2_add_998_U263 ( .QN(P2_add_998_n245), .IN1(P2_add_998_n244), 
        .IN2(P2_add_998_n247) );
  AND2X1 P2_add_998_U262 ( .IN1(P2_add_998_n244), .IN2(P2_add_998_n247), 
        .Q(P2_add_998_n246) );
  NOR2X0 P2_add_998_U261 ( .QN(P2_N4259), .IN1(P2_add_998_n245), 
        .IN2(P2_add_998_n246) );
  NAND2X0 P2_add_998_U260 ( .IN1(n7220), .IN2(P2_add_998_n244), 
        .QN(P2_add_998_n241) );
  OR2X1 P2_add_998_U259 ( .IN2(n7220), .IN1(P2_add_998_n244), 
        .Q(P2_add_998_n243) );
  NAND2X0 P2_add_998_U258 ( .IN1(P2_N4107), .IN2(P2_add_998_n243), 
        .QN(P2_add_998_n242) );
  NAND2X0 P2_add_998_U257 ( .IN1(P2_add_998_n241), .IN2(P2_add_998_n242), 
        .QN(P2_add_998_n234) );
  OR2X1 P2_add_998_U255 ( .IN2(P2_N4108), .IN1(n7214), .Q(P2_add_998_n238) );
  NAND2X0 P2_add_998_U254 ( .IN1(P2_N4108), .IN2(n7214), .QN(P2_add_998_n239)
         );
  NAND2X0 P2_add_998_U253 ( .IN1(P2_add_998_n238), .IN2(P2_add_998_n239), 
        .QN(P2_add_998_n237) );
  NOR2X0 P2_add_998_U252 ( .QN(P2_add_998_n235), .IN1(P2_add_998_n234), 
        .IN2(P2_add_998_n237) );
  AND2X1 P2_add_998_U251 ( .IN1(P2_add_998_n234), .IN2(P2_add_998_n237), 
        .Q(P2_add_998_n236) );
  NOR2X0 P2_add_998_U250 ( .QN(P2_N4260), .IN1(P2_add_998_n235), 
        .IN2(P2_add_998_n236) );
  NAND2X0 P2_add_998_U249 ( .IN1(n7216), .IN2(P2_add_998_n234), 
        .QN(P2_add_998_n231) );
  OR2X1 P2_add_998_U248 ( .IN2(n7216), .IN1(P2_add_998_n234), 
        .Q(P2_add_998_n233) );
  NAND2X0 P2_add_998_U247 ( .IN1(P2_N4108), .IN2(P2_add_998_n233), 
        .QN(P2_add_998_n232) );
  NAND2X0 P2_add_998_U246 ( .IN1(P2_add_998_n231), .IN2(P2_add_998_n232), 
        .QN(P2_add_998_n224) );
  OR2X1 P2_add_998_U244 ( .IN2(P2_N4109), .IN1(n7211), .Q(P2_add_998_n228) );
  NAND2X0 P2_add_998_U243 ( .IN1(P2_N4109), .IN2(n7211), .QN(P2_add_998_n229)
         );
  NAND2X0 P2_add_998_U242 ( .IN1(P2_add_998_n228), .IN2(P2_add_998_n229), 
        .QN(P2_add_998_n227) );
  NOR2X0 P2_add_998_U241 ( .QN(P2_add_998_n225), .IN1(P2_add_998_n224), 
        .IN2(P2_add_998_n227) );
  AND2X1 P2_add_998_U240 ( .IN1(P2_add_998_n224), .IN2(P2_add_998_n227), 
        .Q(P2_add_998_n226) );
  NOR2X0 P2_add_998_U239 ( .QN(P2_N4261), .IN1(P2_add_998_n225), 
        .IN2(P2_add_998_n226) );
  NAND2X0 P2_add_998_U238 ( .IN1(n7210), .IN2(P2_add_998_n224), 
        .QN(P2_add_998_n221) );
  OR2X1 P2_add_998_U237 ( .IN2(n7210), .IN1(P2_add_998_n224), 
        .Q(P2_add_998_n223) );
  NAND2X0 P2_add_998_U236 ( .IN1(P2_N4109), .IN2(P2_add_998_n223), 
        .QN(P2_add_998_n222) );
  NAND2X0 P2_add_998_U235 ( .IN1(P2_add_998_n221), .IN2(P2_add_998_n222), 
        .QN(P2_add_998_n214) );
  OR2X1 P2_add_998_U233 ( .IN2(P2_N4110), .IN1(n7208), .Q(P2_add_998_n218) );
  NAND2X0 P2_add_998_U232 ( .IN1(P2_N4110), .IN2(n7208), .QN(P2_add_998_n219)
         );
  NAND2X0 P2_add_998_U231 ( .IN1(P2_add_998_n218), .IN2(P2_add_998_n219), 
        .QN(P2_add_998_n217) );
  NOR2X0 P2_add_998_U230 ( .QN(P2_add_998_n215), .IN1(P2_add_998_n214), 
        .IN2(P2_add_998_n217) );
  AND2X1 P2_add_998_U229 ( .IN1(P2_add_998_n214), .IN2(P2_add_998_n217), 
        .Q(P2_add_998_n216) );
  NOR2X0 P2_add_998_U228 ( .QN(P2_N4262), .IN1(P2_add_998_n215), 
        .IN2(P2_add_998_n216) );
  NAND2X0 P2_add_998_U227 ( .IN1(n7209), .IN2(P2_add_998_n214), 
        .QN(P2_add_998_n211) );
  OR2X1 P2_add_998_U226 ( .IN2(n7209), .IN1(P2_add_998_n214), 
        .Q(P2_add_998_n213) );
  NAND2X0 P2_add_998_U225 ( .IN1(P2_N4110), .IN2(P2_add_998_n213), 
        .QN(P2_add_998_n212) );
  NAND2X0 P2_add_998_U224 ( .IN1(P2_add_998_n211), .IN2(P2_add_998_n212), 
        .QN(P2_add_998_n204) );
  OR2X1 P2_add_998_U222 ( .IN2(P2_N4111), .IN1(n7205), .Q(P2_add_998_n208) );
  NAND2X0 P2_add_998_U221 ( .IN1(P2_N4111), .IN2(n7205), .QN(P2_add_998_n209)
         );
  NAND2X0 P2_add_998_U220 ( .IN1(P2_add_998_n208), .IN2(P2_add_998_n209), 
        .QN(P2_add_998_n207) );
  NOR2X0 P2_add_998_U219 ( .QN(P2_add_998_n205), .IN1(P2_add_998_n204), 
        .IN2(P2_add_998_n207) );
  AND2X1 P2_add_998_U218 ( .IN1(P2_add_998_n204), .IN2(P2_add_998_n207), 
        .Q(P2_add_998_n206) );
  NOR2X0 P2_add_998_U217 ( .QN(P2_N4263), .IN1(P2_add_998_n205), 
        .IN2(P2_add_998_n206) );
  NAND2X0 P2_add_998_U216 ( .IN1(n7206), .IN2(P2_add_998_n204), 
        .QN(P2_add_998_n201) );
  INVX0 P2_add_998_U7 ( .ZN(P2_add_998_n49), .INP(n7158) );
  INVX0 P2_add_998_U14 ( .ZN(P2_add_998_n296), .INP(n7238) );
  NAND2X0 P2_sub_1030_U54 ( .IN1(n6664), .IN2(n6733), .QN(P2_sub_1030_n61) );
  NAND2X0 P2_sub_1030_U53 ( .IN1(P2_N362), .IN2(n18939), .QN(P2_sub_1030_n62)
         );
  NAND2X0 P2_sub_1030_U52 ( .IN1(P2_sub_1030_n61), .IN2(P2_sub_1030_n62), 
        .QN(P2_sub_1030_n59) );
  NAND2X0 P2_sub_1030_U51 ( .IN1(P2_sub_1030_n59), .IN2(P2_sub_1030_n60), 
        .QN(P2_sub_1030_n57) );
  OR2X1 P2_sub_1030_U50 ( .IN2(P2_sub_1030_n60), .IN1(P2_sub_1030_n59), 
        .Q(P2_sub_1030_n58) );
  NAND2X0 P2_sub_1030_U49 ( .IN1(P2_sub_1030_n57), .IN2(P2_sub_1030_n58), 
        .QN(P2_N4844) );
  NAND2X0 P2_sub_1030_U48 ( .IN1(n6665), .IN2(n6735), .QN(P2_sub_1030_n54) );
  OR2X1 P2_sub_1030_U47 ( .IN2(n6665), .IN1(n6735), .Q(P2_sub_1030_n55) );
  NAND2X0 P2_sub_1030_U46 ( .IN1(P2_sub_1030_n54), .IN2(P2_sub_1030_n55), 
        .QN(P2_sub_1030_n52) );
  NAND2X0 P2_sub_1030_U45 ( .IN1(P2_sub_1030_n52), .IN2(P2_sub_1030_n53), 
        .QN(P2_sub_1030_n50) );
  OR2X1 P2_sub_1030_U44 ( .IN2(P2_sub_1030_n53), .IN1(P2_sub_1030_n52), 
        .Q(P2_sub_1030_n51) );
  NAND2X0 P2_sub_1030_U43 ( .IN1(P2_sub_1030_n50), .IN2(P2_sub_1030_n51), 
        .QN(P2_N4845) );
  NAND2X0 P2_sub_1030_U42 ( .IN1(n6666), .IN2(n6743), .QN(P2_sub_1030_n47) );
  OR2X1 P2_sub_1030_U41 ( .IN2(n6666), .IN1(n6743), .Q(P2_sub_1030_n48) );
  NAND2X0 P2_sub_1030_U40 ( .IN1(P2_sub_1030_n47), .IN2(P2_sub_1030_n48), 
        .QN(P2_sub_1030_n45) );
  NAND2X0 P2_sub_1030_U39 ( .IN1(P2_sub_1030_n45), .IN2(P2_sub_1030_n46), 
        .QN(P2_sub_1030_n43) );
  OR2X1 P2_sub_1030_U38 ( .IN2(P2_sub_1030_n46), .IN1(P2_sub_1030_n45), 
        .Q(P2_sub_1030_n44) );
  NAND2X0 P2_sub_1030_U37 ( .IN1(P2_sub_1030_n43), .IN2(P2_sub_1030_n44), 
        .QN(P2_N4846) );
  NAND2X0 P2_sub_1030_U36 ( .IN1(n6667), .IN2(n6745), .QN(P2_sub_1030_n40) );
  OR2X1 P2_sub_1030_U35 ( .IN2(n6667), .IN1(n6745), .Q(P2_sub_1030_n41) );
  NAND2X0 P2_sub_1030_U34 ( .IN1(P2_sub_1030_n40), .IN2(P2_sub_1030_n41), 
        .QN(P2_sub_1030_n38) );
  NAND2X0 P2_sub_1030_U33 ( .IN1(P2_sub_1030_n38), .IN2(P2_sub_1030_n39), 
        .QN(P2_sub_1030_n36) );
  OR2X1 P2_sub_1030_U32 ( .IN2(P2_sub_1030_n39), .IN1(P2_sub_1030_n38), 
        .Q(P2_sub_1030_n37) );
  NAND2X0 P2_sub_1030_U31 ( .IN1(P2_sub_1030_n36), .IN2(P2_sub_1030_n37), 
        .QN(P2_N4847) );
  NAND2X0 P2_sub_1030_U30 ( .IN1(n6668), .IN2(n6749), .QN(P2_sub_1030_n33) );
  OR2X1 P2_sub_1030_U29 ( .IN2(n6668), .IN1(n6749), .Q(P2_sub_1030_n34) );
  NAND2X0 P2_sub_1030_U28 ( .IN1(P2_sub_1030_n33), .IN2(P2_sub_1030_n34), 
        .QN(P2_sub_1030_n31) );
  NAND2X0 P2_sub_1030_U27 ( .IN1(P2_sub_1030_n31), .IN2(P2_sub_1030_n32), 
        .QN(P2_sub_1030_n29) );
  OR2X1 P2_sub_1030_U26 ( .IN2(P2_sub_1030_n32), .IN1(P2_sub_1030_n31), 
        .Q(P2_sub_1030_n30) );
  NAND2X0 P2_sub_1030_U25 ( .IN1(P2_sub_1030_n29), .IN2(P2_sub_1030_n30), 
        .QN(P2_N4848) );
  NAND2X0 P2_sub_1030_U24 ( .IN1(n6669), .IN2(n6753), .QN(P2_sub_1030_n26) );
  OR2X1 P2_sub_1030_U23 ( .IN2(n6669), .IN1(n6753), .Q(P2_sub_1030_n27) );
  NAND2X0 P2_sub_1030_U22 ( .IN1(P2_sub_1030_n26), .IN2(P2_sub_1030_n27), 
        .QN(P2_sub_1030_n24) );
  NAND2X0 P2_sub_1030_U21 ( .IN1(P2_sub_1030_n24), .IN2(P2_sub_1030_n25), 
        .QN(P2_sub_1030_n22) );
  OR2X1 P2_sub_1030_U20 ( .IN2(P2_sub_1030_n25), .IN1(P2_sub_1030_n24), 
        .Q(P2_sub_1030_n23) );
  NAND2X0 P2_sub_1030_U19 ( .IN1(P2_sub_1030_n22), .IN2(P2_sub_1030_n23), 
        .QN(P2_N4849) );
  NAND2X0 P2_sub_1030_U18 ( .IN1(n6670), .IN2(n6748), .QN(P2_sub_1030_n19) );
  OR2X1 P2_sub_1030_U17 ( .IN2(n6670), .IN1(n6748), .Q(P2_sub_1030_n20) );
  NAND2X0 P2_sub_1030_U16 ( .IN1(P2_sub_1030_n19), .IN2(P2_sub_1030_n20), 
        .QN(P2_sub_1030_n17) );
  NAND2X0 P2_sub_1030_U15 ( .IN1(P2_sub_1030_n17), .IN2(P2_sub_1030_n18), 
        .QN(P2_sub_1030_n15) );
  OR2X1 P2_sub_1030_U14 ( .IN2(P2_sub_1030_n18), .IN1(P2_sub_1030_n17), 
        .Q(P2_sub_1030_n16) );
  NAND2X0 P2_sub_1030_U13 ( .IN1(P2_sub_1030_n15), .IN2(P2_sub_1030_n16), 
        .QN(P2_N4850) );
  NAND2X0 P2_sub_1030_U12 ( .IN1(n10249), .IN2(n6752), .QN(P2_sub_1030_n12) );
  OR2X1 P2_sub_1030_U11 ( .IN2(n10249), .IN1(n6752), .Q(P2_sub_1030_n13) );
  NAND2X0 P2_sub_1030_U10 ( .IN1(P2_sub_1030_n12), .IN2(P2_sub_1030_n13), 
        .QN(P2_sub_1030_n10) );
  NAND2X0 P2_sub_1030_U9 ( .IN1(P2_sub_1030_n10), .IN2(P2_sub_1030_n11), 
        .QN(P2_sub_1030_n8) );
  OR2X1 P2_sub_1030_U8 ( .IN2(P2_sub_1030_n11), .IN1(P2_sub_1030_n10), 
        .Q(P2_sub_1030_n9) );
  NAND2X0 P2_sub_1030_U7 ( .IN1(P2_sub_1030_n8), .IN2(P2_sub_1030_n9), 
        .QN(P2_N4851) );
  NAND2X0 P2_sub_1030_U6 ( .IN1(n6671), .IN2(n6757), .QN(P2_sub_1030_n5) );
  OR2X1 P2_sub_1030_U5 ( .IN2(n6671), .IN1(n6757), .Q(P2_sub_1030_n6) );
  NAND2X0 P2_sub_1030_U4 ( .IN1(P2_sub_1030_n5), .IN2(P2_sub_1030_n6), 
        .QN(P2_sub_1030_n3) );
  NAND2X0 P2_sub_1030_U3 ( .IN1(P2_sub_1030_n3), .IN2(P2_sub_1030_n4), 
        .QN(P2_sub_1030_n1) );
  OR2X1 P2_sub_1030_U2 ( .IN2(P2_sub_1030_n4), .IN1(P2_sub_1030_n3), 
        .Q(P2_sub_1030_n2) );
  NAND2X0 P2_sub_1030_U1 ( .IN1(P2_sub_1030_n1), .IN2(P2_sub_1030_n2), 
        .QN(P2_N4852) );
  NAND2X0 P2_sub_1030_U147 ( .IN1(P2_sub_1030_n152), .IN2(n6760), 
        .QN(P2_sub_1030_n151) );
  NAND2X0 P2_sub_1030_U146 ( .IN1(P2_sub_1030_n150), .IN2(P2_sub_1030_n151), 
        .QN(P2_sub_1030_n144) );
  NAND2X0 P2_sub_1030_U145 ( .IN1(P2_sub_1030_n149), .IN2(P2_sub_1030_n144), 
        .QN(P2_sub_1030_n147) );
  OR2X1 P2_sub_1030_U144 ( .IN2(P2_sub_1030_n144), .IN1(P2_sub_1030_n149), 
        .Q(P2_sub_1030_n148) );
  NAND2X0 P2_sub_1030_U143 ( .IN1(P2_sub_1030_n147), .IN2(P2_sub_1030_n148), 
        .QN(P2_N4854) );
  NAND2X0 P2_sub_1030_U141 ( .IN1(n6674), .IN2(n6761), .QN(P2_sub_1030_n145)
         );
  OR2X1 P2_sub_1030_U140 ( .IN2(n6674), .IN1(n6761), .Q(P2_sub_1030_n146) );
  NAND2X0 P2_sub_1030_U139 ( .IN1(P2_sub_1030_n145), .IN2(P2_sub_1030_n146), 
        .QN(P2_sub_1030_n139) );
  NAND2X0 P2_sub_1030_U138 ( .IN1(n6673), .IN2(P2_sub_1030_n144), 
        .QN(P2_sub_1030_n140) );
  OR2X1 P2_sub_1030_U137 ( .IN2(n6673), .IN1(P2_sub_1030_n144), 
        .Q(P2_sub_1030_n142) );
  NAND2X0 P2_sub_1030_U136 ( .IN1(P2_sub_1030_n142), .IN2(n6756), 
        .QN(P2_sub_1030_n141) );
  NAND2X0 P2_sub_1030_U135 ( .IN1(P2_sub_1030_n140), .IN2(P2_sub_1030_n141), 
        .QN(P2_sub_1030_n134) );
  NAND2X0 P2_sub_1030_U134 ( .IN1(P2_sub_1030_n139), .IN2(P2_sub_1030_n134), 
        .QN(P2_sub_1030_n137) );
  OR2X1 P2_sub_1030_U133 ( .IN2(P2_sub_1030_n134), .IN1(P2_sub_1030_n139), 
        .Q(P2_sub_1030_n138) );
  NAND2X0 P2_sub_1030_U132 ( .IN1(P2_sub_1030_n137), .IN2(P2_sub_1030_n138), 
        .QN(P2_N4855) );
  NAND2X0 P2_sub_1030_U130 ( .IN1(n6675), .IN2(n6765), .QN(P2_sub_1030_n135)
         );
  OR2X1 P2_sub_1030_U129 ( .IN2(n6675), .IN1(n6765), .Q(P2_sub_1030_n136) );
  NAND2X0 P2_sub_1030_U128 ( .IN1(P2_sub_1030_n135), .IN2(P2_sub_1030_n136), 
        .QN(P2_sub_1030_n129) );
  NAND2X0 P2_sub_1030_U127 ( .IN1(n6674), .IN2(P2_sub_1030_n134), 
        .QN(P2_sub_1030_n130) );
  OR2X1 P2_sub_1030_U126 ( .IN2(n6674), .IN1(P2_sub_1030_n134), 
        .Q(P2_sub_1030_n132) );
  NAND2X0 P2_sub_1030_U125 ( .IN1(P2_sub_1030_n132), .IN2(n6761), 
        .QN(P2_sub_1030_n131) );
  NAND2X0 P2_sub_1030_U124 ( .IN1(P2_sub_1030_n130), .IN2(P2_sub_1030_n131), 
        .QN(P2_sub_1030_n124) );
  NAND2X0 P2_sub_1030_U123 ( .IN1(P2_sub_1030_n129), .IN2(P2_sub_1030_n124), 
        .QN(P2_sub_1030_n127) );
  OR2X1 P2_sub_1030_U122 ( .IN2(P2_sub_1030_n124), .IN1(P2_sub_1030_n129), 
        .Q(P2_sub_1030_n128) );
  NAND2X0 P2_sub_1030_U121 ( .IN1(P2_sub_1030_n127), .IN2(P2_sub_1030_n128), 
        .QN(P2_N4856) );
  NAND2X0 P2_sub_1030_U119 ( .IN1(n6676), .IN2(n6769), .QN(P2_sub_1030_n125)
         );
  OR2X1 P2_sub_1030_U118 ( .IN2(n6676), .IN1(n6769), .Q(P2_sub_1030_n126) );
  NAND2X0 P2_sub_1030_U117 ( .IN1(P2_sub_1030_n125), .IN2(P2_sub_1030_n126), 
        .QN(P2_sub_1030_n119) );
  NAND2X0 P2_sub_1030_U116 ( .IN1(n6675), .IN2(P2_sub_1030_n124), 
        .QN(P2_sub_1030_n120) );
  OR2X1 P2_sub_1030_U115 ( .IN2(n6675), .IN1(P2_sub_1030_n124), 
        .Q(P2_sub_1030_n122) );
  NAND2X0 P2_sub_1030_U114 ( .IN1(P2_sub_1030_n122), .IN2(n6765), 
        .QN(P2_sub_1030_n121) );
  NAND2X0 P2_sub_1030_U113 ( .IN1(P2_sub_1030_n120), .IN2(P2_sub_1030_n121), 
        .QN(P2_sub_1030_n114) );
  NAND2X0 P2_sub_1030_U112 ( .IN1(P2_sub_1030_n119), .IN2(P2_sub_1030_n114), 
        .QN(P2_sub_1030_n117) );
  OR2X1 P2_sub_1030_U111 ( .IN2(P2_sub_1030_n114), .IN1(P2_sub_1030_n119), 
        .Q(P2_sub_1030_n118) );
  NAND2X0 P2_sub_1030_U110 ( .IN1(P2_sub_1030_n117), .IN2(P2_sub_1030_n118), 
        .QN(P2_N4857) );
  NAND2X0 P2_sub_1030_U108 ( .IN1(n6677), .IN2(n6764), .QN(P2_sub_1030_n115)
         );
  OR2X1 P2_sub_1030_U107 ( .IN2(n6677), .IN1(n6764), .Q(P2_sub_1030_n116) );
  NAND2X0 P2_sub_1030_U106 ( .IN1(P2_sub_1030_n115), .IN2(P2_sub_1030_n116), 
        .QN(P2_sub_1030_n109) );
  NAND2X0 P2_sub_1030_U105 ( .IN1(n6676), .IN2(P2_sub_1030_n114), 
        .QN(P2_sub_1030_n110) );
  OR2X1 P2_sub_1030_U104 ( .IN2(n6676), .IN1(P2_sub_1030_n114), 
        .Q(P2_sub_1030_n112) );
  NAND2X0 P2_sub_1030_U103 ( .IN1(P2_sub_1030_n112), .IN2(n6769), 
        .QN(P2_sub_1030_n111) );
  NAND2X0 P2_sub_1030_U102 ( .IN1(P2_sub_1030_n110), .IN2(P2_sub_1030_n111), 
        .QN(P2_sub_1030_n104) );
  NAND2X0 P2_sub_1030_U101 ( .IN1(P2_sub_1030_n109), .IN2(P2_sub_1030_n104), 
        .QN(P2_sub_1030_n107) );
  OR2X1 P2_sub_1030_U100 ( .IN2(P2_sub_1030_n104), .IN1(P2_sub_1030_n109), 
        .Q(P2_sub_1030_n108) );
  NAND2X0 P2_sub_1030_U99 ( .IN1(P2_sub_1030_n107), .IN2(P2_sub_1030_n108), 
        .QN(P2_N4858) );
  NAND2X0 P2_sub_1030_U97 ( .IN1(n6678), .IN2(n6768), .QN(P2_sub_1030_n105) );
  OR2X1 P2_sub_1030_U96 ( .IN2(n6678), .IN1(n6768), .Q(P2_sub_1030_n106) );
  NAND2X0 P2_sub_1030_U95 ( .IN1(P2_sub_1030_n105), .IN2(P2_sub_1030_n106), 
        .QN(P2_sub_1030_n99) );
  NAND2X0 P2_sub_1030_U94 ( .IN1(n6677), .IN2(P2_sub_1030_n104), 
        .QN(P2_sub_1030_n100) );
  OR2X1 P2_sub_1030_U93 ( .IN2(n6677), .IN1(P2_sub_1030_n104), 
        .Q(P2_sub_1030_n102) );
  NAND2X0 P2_sub_1030_U92 ( .IN1(P2_sub_1030_n102), .IN2(n6764), 
        .QN(P2_sub_1030_n101) );
  NAND2X0 P2_sub_1030_U91 ( .IN1(P2_sub_1030_n100), .IN2(P2_sub_1030_n101), 
        .QN(P2_sub_1030_n94) );
  NAND2X0 P2_sub_1030_U90 ( .IN1(P2_sub_1030_n99), .IN2(P2_sub_1030_n94), 
        .QN(P2_sub_1030_n97) );
  OR2X1 P2_sub_1030_U89 ( .IN2(P2_sub_1030_n94), .IN1(P2_sub_1030_n99), 
        .Q(P2_sub_1030_n98) );
  NAND2X0 P2_sub_1030_U88 ( .IN1(P2_sub_1030_n97), .IN2(P2_sub_1030_n98), 
        .QN(P2_N4859) );
  NAND2X0 P2_sub_1030_U86 ( .IN1(n6679), .IN2(n6772), .QN(P2_sub_1030_n95) );
  OR2X1 P2_sub_1030_U85 ( .IN2(n6679), .IN1(n6772), .Q(P2_sub_1030_n96) );
  NAND2X0 P2_sub_1030_U84 ( .IN1(P2_sub_1030_n95), .IN2(P2_sub_1030_n96), 
        .QN(P2_sub_1030_n89) );
  NAND2X0 P2_sub_1030_U83 ( .IN1(n6678), .IN2(P2_sub_1030_n94), 
        .QN(P2_sub_1030_n90) );
  OR2X1 P2_sub_1030_U82 ( .IN2(n6678), .IN1(P2_sub_1030_n94), 
        .Q(P2_sub_1030_n92) );
  NAND2X0 P2_sub_1030_U81 ( .IN1(P2_sub_1030_n92), .IN2(n6768), 
        .QN(P2_sub_1030_n91) );
  NAND2X0 P2_sub_1030_U80 ( .IN1(P2_sub_1030_n90), .IN2(P2_sub_1030_n91), 
        .QN(P2_sub_1030_n84) );
  NAND2X0 P2_sub_1030_U79 ( .IN1(P2_sub_1030_n89), .IN2(P2_sub_1030_n84), 
        .QN(P2_sub_1030_n87) );
  OR2X1 P2_sub_1030_U78 ( .IN2(P2_sub_1030_n84), .IN1(P2_sub_1030_n89), 
        .Q(P2_sub_1030_n88) );
  NAND2X0 P2_sub_1030_U77 ( .IN1(P2_sub_1030_n87), .IN2(P2_sub_1030_n88), 
        .QN(P2_N4860) );
  NAND2X0 P2_sub_1030_U75 ( .IN1(n6680), .IN2(n6774), .QN(P2_sub_1030_n85) );
  OR2X1 P2_sub_1030_U74 ( .IN2(n6680), .IN1(n6774), .Q(P2_sub_1030_n86) );
  NAND2X0 P2_sub_1030_U73 ( .IN1(P2_sub_1030_n85), .IN2(P2_sub_1030_n86), 
        .QN(P2_sub_1030_n79) );
  NAND2X0 P2_sub_1030_U72 ( .IN1(n6679), .IN2(P2_sub_1030_n84), 
        .QN(P2_sub_1030_n80) );
  OR2X1 P2_sub_1030_U71 ( .IN2(n6679), .IN1(P2_sub_1030_n84), 
        .Q(P2_sub_1030_n82) );
  NAND2X0 P2_sub_1030_U70 ( .IN1(P2_sub_1030_n82), .IN2(n6772), 
        .QN(P2_sub_1030_n81) );
  NAND2X0 P2_sub_1030_U69 ( .IN1(P2_sub_1030_n80), .IN2(P2_sub_1030_n81), 
        .QN(P2_sub_1030_n73) );
  NAND2X0 P2_sub_1030_U68 ( .IN1(P2_sub_1030_n79), .IN2(P2_sub_1030_n73), 
        .QN(P2_sub_1030_n77) );
  OR2X1 P2_sub_1030_U67 ( .IN2(P2_sub_1030_n73), .IN1(P2_sub_1030_n79), 
        .Q(P2_sub_1030_n78) );
  NAND2X0 P2_sub_1030_U66 ( .IN1(P2_sub_1030_n77), .IN2(P2_sub_1030_n78), 
        .QN(P2_N4861) );
  INVX0 P2_sub_1030_U65 ( .ZN(P2_sub_1030_n76), .INP(n10111) );
  OR2X1 P2_sub_1030_U64 ( .IN2(P2_N344), .IN1(P2_sub_1030_n76), 
        .Q(P2_sub_1030_n74) );
  NAND2X0 P2_sub_1030_U63 ( .IN1(P2_N344), .IN2(P2_sub_1030_n76), 
        .QN(P2_sub_1030_n75) );
  NAND2X0 P2_sub_1030_U62 ( .IN1(P2_sub_1030_n74), .IN2(P2_sub_1030_n75), 
        .QN(P2_sub_1030_n68) );
  NAND2X0 P2_sub_1030_U61 ( .IN1(n6680), .IN2(P2_sub_1030_n73), 
        .QN(P2_sub_1030_n69) );
  OR2X1 P2_sub_1030_U60 ( .IN2(n6680), .IN1(P2_sub_1030_n73), 
        .Q(P2_sub_1030_n71) );
  NAND2X0 P2_sub_1030_U59 ( .IN1(P2_sub_1030_n71), .IN2(n6774), 
        .QN(P2_sub_1030_n70) );
  NAND2X0 P2_sub_1030_U58 ( .IN1(P2_sub_1030_n69), .IN2(P2_sub_1030_n70), 
        .QN(P2_sub_1030_n67) );
  NAND2X0 P2_sub_1030_U57 ( .IN1(P2_sub_1030_n68), .IN2(P2_sub_1030_n67), 
        .QN(P2_sub_1030_n65) );
  OR2X1 P2_sub_1030_U56 ( .IN2(P2_sub_1030_n68), .IN1(P2_sub_1030_n67), 
        .Q(P2_sub_1030_n66) );
  NAND2X0 P2_sub_1030_U55 ( .IN1(P2_sub_1030_n65), .IN2(P2_sub_1030_n66), 
        .QN(P2_N4862) );
  NOR2X0 P2_sub_1030_U210 ( .QN(P2_sub_1030_n187), .IN1(n6731), .IN2(n9837) );
  INVX0 P2_sub_1030_U209 ( .ZN(P2_sub_1030_n60), .INP(P2_sub_1030_n187) );
  NAND2X0 P2_sub_1030_U208 ( .IN1(n9837), .IN2(n6731), .QN(P2_sub_1030_n190)
         );
  NAND2X0 P2_sub_1030_U207 ( .IN1(P2_sub_1030_n60), .IN2(P2_sub_1030_n190), 
        .QN(P2_N4843) );
  NAND2X0 P2_sub_1030_U205 ( .IN1(n6672), .IN2(n6760), .QN(P2_sub_1030_n188)
         );
  OR2X1 P2_sub_1030_U204 ( .IN2(n6672), .IN1(n6760), .Q(P2_sub_1030_n189) );
  NAND2X0 P2_sub_1030_U203 ( .IN1(P2_sub_1030_n188), .IN2(P2_sub_1030_n189), 
        .QN(P2_sub_1030_n159) );
  NAND2X0 P2_sub_1030_U202 ( .IN1(n6664), .IN2(P2_sub_1030_n60), 
        .QN(P2_sub_1030_n184) );
  NAND2X0 P2_sub_1030_U200 ( .IN1(P2_sub_1030_n187), .IN2(n18939), 
        .QN(P2_sub_1030_n186) );
  NAND2X0 P2_sub_1030_U198 ( .IN1(P2_sub_1030_n186), .IN2(n6733), 
        .QN(P2_sub_1030_n185) );
  NAND2X0 P2_sub_1030_U197 ( .IN1(P2_sub_1030_n184), .IN2(P2_sub_1030_n185), 
        .QN(P2_sub_1030_n53) );
  NAND2X0 P2_sub_1030_U196 ( .IN1(n6665), .IN2(P2_sub_1030_n53), 
        .QN(P2_sub_1030_n181) );
  OR2X1 P2_sub_1030_U195 ( .IN2(n6665), .IN1(P2_sub_1030_n53), 
        .Q(P2_sub_1030_n183) );
  NAND2X0 P2_sub_1030_U193 ( .IN1(P2_sub_1030_n183), .IN2(n6735), 
        .QN(P2_sub_1030_n182) );
  NAND2X0 P2_sub_1030_U192 ( .IN1(P2_sub_1030_n181), .IN2(P2_sub_1030_n182), 
        .QN(P2_sub_1030_n46) );
  NAND2X0 P2_sub_1030_U191 ( .IN1(n6666), .IN2(P2_sub_1030_n46), 
        .QN(P2_sub_1030_n178) );
  OR2X1 P2_sub_1030_U190 ( .IN2(n6666), .IN1(P2_sub_1030_n46), 
        .Q(P2_sub_1030_n180) );
  NAND2X0 P2_sub_1030_U188 ( .IN1(P2_sub_1030_n180), .IN2(n6743), 
        .QN(P2_sub_1030_n179) );
  NAND2X0 P2_sub_1030_U187 ( .IN1(P2_sub_1030_n178), .IN2(P2_sub_1030_n179), 
        .QN(P2_sub_1030_n39) );
  NAND2X0 P2_sub_1030_U186 ( .IN1(n6667), .IN2(P2_sub_1030_n39), 
        .QN(P2_sub_1030_n175) );
  OR2X1 P2_sub_1030_U185 ( .IN2(n6667), .IN1(P2_sub_1030_n39), 
        .Q(P2_sub_1030_n177) );
  NAND2X0 P2_sub_1030_U183 ( .IN1(P2_sub_1030_n177), .IN2(n6745), 
        .QN(P2_sub_1030_n176) );
  NAND2X0 P2_sub_1030_U182 ( .IN1(P2_sub_1030_n175), .IN2(P2_sub_1030_n176), 
        .QN(P2_sub_1030_n32) );
  NAND2X0 P2_sub_1030_U181 ( .IN1(n6668), .IN2(P2_sub_1030_n32), 
        .QN(P2_sub_1030_n172) );
  OR2X1 P2_sub_1030_U180 ( .IN2(n6668), .IN1(P2_sub_1030_n32), 
        .Q(P2_sub_1030_n174) );
  NAND2X0 P2_sub_1030_U178 ( .IN1(P2_sub_1030_n174), .IN2(n6749), 
        .QN(P2_sub_1030_n173) );
  NAND2X0 P2_sub_1030_U177 ( .IN1(P2_sub_1030_n172), .IN2(P2_sub_1030_n173), 
        .QN(P2_sub_1030_n25) );
  NAND2X0 P2_sub_1030_U176 ( .IN1(n6669), .IN2(P2_sub_1030_n25), 
        .QN(P2_sub_1030_n169) );
  OR2X1 P2_sub_1030_U175 ( .IN2(n6669), .IN1(P2_sub_1030_n25), 
        .Q(P2_sub_1030_n171) );
  NAND2X0 P2_sub_1030_U173 ( .IN1(P2_sub_1030_n171), .IN2(n6753), 
        .QN(P2_sub_1030_n170) );
  NAND2X0 P2_sub_1030_U172 ( .IN1(P2_sub_1030_n169), .IN2(P2_sub_1030_n170), 
        .QN(P2_sub_1030_n18) );
  NAND2X0 P2_sub_1030_U171 ( .IN1(n6670), .IN2(P2_sub_1030_n18), 
        .QN(P2_sub_1030_n166) );
  OR2X1 P2_sub_1030_U170 ( .IN2(n6670), .IN1(P2_sub_1030_n18), 
        .Q(P2_sub_1030_n168) );
  NAND2X0 P2_sub_1030_U168 ( .IN1(P2_sub_1030_n168), .IN2(n6748), 
        .QN(P2_sub_1030_n167) );
  NAND2X0 P2_sub_1030_U167 ( .IN1(P2_sub_1030_n166), .IN2(P2_sub_1030_n167), 
        .QN(P2_sub_1030_n11) );
  NAND2X0 P2_sub_1030_U166 ( .IN1(n10249), .IN2(P2_sub_1030_n11), 
        .QN(P2_sub_1030_n163) );
  OR2X1 P2_sub_1030_U165 ( .IN2(n10249), .IN1(P2_sub_1030_n11), 
        .Q(P2_sub_1030_n165) );
  NAND2X0 P2_sub_1030_U163 ( .IN1(P2_sub_1030_n165), .IN2(n6752), 
        .QN(P2_sub_1030_n164) );
  NAND2X0 P2_sub_1030_U162 ( .IN1(P2_sub_1030_n163), .IN2(P2_sub_1030_n164), 
        .QN(P2_sub_1030_n4) );
  NAND2X0 P2_sub_1030_U161 ( .IN1(n6671), .IN2(P2_sub_1030_n4), 
        .QN(P2_sub_1030_n160) );
  OR2X1 P2_sub_1030_U160 ( .IN2(n6671), .IN1(P2_sub_1030_n4), 
        .Q(P2_sub_1030_n162) );
  NAND2X0 P2_sub_1030_U158 ( .IN1(P2_sub_1030_n162), .IN2(n6757), 
        .QN(P2_sub_1030_n161) );
  NAND2X0 P2_sub_1030_U157 ( .IN1(P2_sub_1030_n160), .IN2(P2_sub_1030_n161), 
        .QN(P2_sub_1030_n154) );
  NAND2X0 P2_sub_1030_U156 ( .IN1(P2_sub_1030_n159), .IN2(P2_sub_1030_n154), 
        .QN(P2_sub_1030_n157) );
  OR2X1 P2_sub_1030_U155 ( .IN2(P2_sub_1030_n154), .IN1(P2_sub_1030_n159), 
        .Q(P2_sub_1030_n158) );
  NAND2X0 P2_sub_1030_U154 ( .IN1(P2_sub_1030_n157), .IN2(P2_sub_1030_n158), 
        .QN(P2_N4853) );
  NAND2X0 P2_sub_1030_U152 ( .IN1(n6673), .IN2(n6756), .QN(P2_sub_1030_n155)
         );
  OR2X1 P2_sub_1030_U151 ( .IN2(n6673), .IN1(n6756), .Q(P2_sub_1030_n156) );
  NAND2X0 P2_sub_1030_U150 ( .IN1(P2_sub_1030_n155), .IN2(P2_sub_1030_n156), 
        .QN(P2_sub_1030_n149) );
  NAND2X0 P2_sub_1030_U149 ( .IN1(n6672), .IN2(P2_sub_1030_n154), 
        .QN(P2_sub_1030_n150) );
  OR2X1 P2_sub_1030_U148 ( .IN2(n6672), .IN1(P2_sub_1030_n154), 
        .Q(P2_sub_1030_n152) );
  NAND2X0 P2_sub_1031_U79 ( .IN1(P2_sub_1031_n89), .IN2(P2_sub_1031_n84), 
        .QN(P2_sub_1031_n87) );
  OR2X1 P2_sub_1031_U78 ( .IN2(P2_sub_1031_n84), .IN1(P2_sub_1031_n89), 
        .Q(P2_sub_1031_n88) );
  NAND2X0 P2_sub_1031_U77 ( .IN1(P2_sub_1031_n87), .IN2(P2_sub_1031_n88), 
        .QN(P2_N4880) );
  NAND2X0 P2_sub_1031_U75 ( .IN1(n6663), .IN2(n6774), .QN(P2_sub_1031_n85) );
  OR2X1 P2_sub_1031_U74 ( .IN2(n6663), .IN1(n6774), .Q(P2_sub_1031_n86) );
  NAND2X0 P2_sub_1031_U73 ( .IN1(P2_sub_1031_n85), .IN2(P2_sub_1031_n86), 
        .QN(P2_sub_1031_n79) );
  NAND2X0 P2_sub_1031_U72 ( .IN1(n6662), .IN2(P2_sub_1031_n84), 
        .QN(P2_sub_1031_n80) );
  OR2X1 P2_sub_1031_U71 ( .IN2(n6662), .IN1(P2_sub_1031_n84), 
        .Q(P2_sub_1031_n82) );
  NAND2X0 P2_sub_1031_U70 ( .IN1(P2_sub_1031_n82), .IN2(n6772), 
        .QN(P2_sub_1031_n81) );
  NAND2X0 P2_sub_1031_U69 ( .IN1(P2_sub_1031_n80), .IN2(P2_sub_1031_n81), 
        .QN(P2_sub_1031_n73) );
  NAND2X0 P2_sub_1031_U68 ( .IN1(P2_sub_1031_n79), .IN2(P2_sub_1031_n73), 
        .QN(P2_sub_1031_n77) );
  OR2X1 P2_sub_1031_U67 ( .IN2(P2_sub_1031_n73), .IN1(P2_sub_1031_n79), 
        .Q(P2_sub_1031_n78) );
  NAND2X0 P2_sub_1031_U66 ( .IN1(P2_sub_1031_n77), .IN2(P2_sub_1031_n78), 
        .QN(P2_N4881) );
  INVX0 P2_sub_1031_U65 ( .ZN(P2_sub_1031_n76), .INP(n10116) );
  OR2X1 P2_sub_1031_U64 ( .IN2(P2_N344), .IN1(P2_sub_1031_n76), 
        .Q(P2_sub_1031_n74) );
  NAND2X0 P2_sub_1031_U63 ( .IN1(P2_N344), .IN2(P2_sub_1031_n76), 
        .QN(P2_sub_1031_n75) );
  NAND2X0 P2_sub_1031_U62 ( .IN1(P2_sub_1031_n74), .IN2(P2_sub_1031_n75), 
        .QN(P2_sub_1031_n68) );
  NAND2X0 P2_sub_1031_U61 ( .IN1(n6663), .IN2(P2_sub_1031_n73), 
        .QN(P2_sub_1031_n69) );
  OR2X1 P2_sub_1031_U60 ( .IN2(n6663), .IN1(P2_sub_1031_n73), 
        .Q(P2_sub_1031_n71) );
  NAND2X0 P2_sub_1031_U59 ( .IN1(P2_sub_1031_n71), .IN2(n6774), 
        .QN(P2_sub_1031_n70) );
  NAND2X0 P2_sub_1031_U58 ( .IN1(P2_sub_1031_n69), .IN2(P2_sub_1031_n70), 
        .QN(P2_sub_1031_n67) );
  NAND2X0 P2_sub_1031_U57 ( .IN1(P2_sub_1031_n68), .IN2(P2_sub_1031_n67), 
        .QN(P2_sub_1031_n65) );
  OR2X1 P2_sub_1031_U56 ( .IN2(P2_sub_1031_n68), .IN1(P2_sub_1031_n67), 
        .Q(P2_sub_1031_n66) );
  NAND2X0 P2_sub_1031_U55 ( .IN1(P2_sub_1031_n65), .IN2(P2_sub_1031_n66), 
        .QN(P2_N4882) );
  NAND2X0 P2_sub_1031_U54 ( .IN1(n6720), .IN2(n6733), .QN(P2_sub_1031_n61) );
  NAND2X0 P2_sub_1031_U53 ( .IN1(P2_N362), .IN2(n18997), .QN(P2_sub_1031_n62)
         );
  NAND2X0 P2_sub_1031_U52 ( .IN1(P2_sub_1031_n61), .IN2(P2_sub_1031_n62), 
        .QN(P2_sub_1031_n59) );
  NAND2X0 P2_sub_1031_U51 ( .IN1(P2_sub_1031_n59), .IN2(P2_sub_1031_n60), 
        .QN(P2_sub_1031_n57) );
  OR2X1 P2_sub_1031_U50 ( .IN2(P2_sub_1031_n60), .IN1(P2_sub_1031_n59), 
        .Q(P2_sub_1031_n58) );
  NAND2X0 P2_sub_1031_U49 ( .IN1(P2_sub_1031_n57), .IN2(P2_sub_1031_n58), 
        .QN(P2_N4864) );
  NAND2X0 P2_sub_1031_U48 ( .IN1(n6721), .IN2(n6735), .QN(P2_sub_1031_n54) );
  OR2X1 P2_sub_1031_U47 ( .IN2(n6721), .IN1(n6735), .Q(P2_sub_1031_n55) );
  NAND2X0 P2_sub_1031_U46 ( .IN1(P2_sub_1031_n54), .IN2(P2_sub_1031_n55), 
        .QN(P2_sub_1031_n52) );
  NAND2X0 P2_sub_1031_U45 ( .IN1(P2_sub_1031_n52), .IN2(P2_sub_1031_n53), 
        .QN(P2_sub_1031_n50) );
  OR2X1 P2_sub_1031_U44 ( .IN2(P2_sub_1031_n53), .IN1(P2_sub_1031_n52), 
        .Q(P2_sub_1031_n51) );
  NAND2X0 P2_sub_1031_U43 ( .IN1(P2_sub_1031_n50), .IN2(P2_sub_1031_n51), 
        .QN(P2_N4865) );
  NAND2X0 P2_sub_1031_U42 ( .IN1(n6648), .IN2(n6743), .QN(P2_sub_1031_n47) );
  OR2X1 P2_sub_1031_U41 ( .IN2(n6648), .IN1(n6743), .Q(P2_sub_1031_n48) );
  NAND2X0 P2_sub_1031_U40 ( .IN1(P2_sub_1031_n47), .IN2(P2_sub_1031_n48), 
        .QN(P2_sub_1031_n45) );
  NAND2X0 P2_sub_1031_U39 ( .IN1(P2_sub_1031_n45), .IN2(P2_sub_1031_n46), 
        .QN(P2_sub_1031_n43) );
  OR2X1 P2_sub_1031_U38 ( .IN2(P2_sub_1031_n46), .IN1(P2_sub_1031_n45), 
        .Q(P2_sub_1031_n44) );
  NAND2X0 P2_sub_1031_U37 ( .IN1(P2_sub_1031_n43), .IN2(P2_sub_1031_n44), 
        .QN(P2_N4866) );
  NAND2X0 P2_sub_1031_U36 ( .IN1(n6649), .IN2(n6745), .QN(P2_sub_1031_n40) );
  OR2X1 P2_sub_1031_U35 ( .IN2(n6649), .IN1(n6745), .Q(P2_sub_1031_n41) );
  NAND2X0 P2_sub_1031_U34 ( .IN1(P2_sub_1031_n40), .IN2(P2_sub_1031_n41), 
        .QN(P2_sub_1031_n38) );
  NAND2X0 P2_sub_1031_U33 ( .IN1(P2_sub_1031_n38), .IN2(P2_sub_1031_n39), 
        .QN(P2_sub_1031_n36) );
  OR2X1 P2_sub_1031_U32 ( .IN2(P2_sub_1031_n39), .IN1(P2_sub_1031_n38), 
        .Q(P2_sub_1031_n37) );
  NAND2X0 P2_sub_1031_U31 ( .IN1(P2_sub_1031_n36), .IN2(P2_sub_1031_n37), 
        .QN(P2_N4867) );
  NAND2X0 P2_sub_1031_U30 ( .IN1(n6650), .IN2(n6749), .QN(P2_sub_1031_n33) );
  OR2X1 P2_sub_1031_U29 ( .IN2(n6650), .IN1(n6749), .Q(P2_sub_1031_n34) );
  NAND2X0 P2_sub_1031_U28 ( .IN1(P2_sub_1031_n33), .IN2(P2_sub_1031_n34), 
        .QN(P2_sub_1031_n31) );
  NAND2X0 P2_sub_1031_U27 ( .IN1(P2_sub_1031_n31), .IN2(P2_sub_1031_n32), 
        .QN(P2_sub_1031_n29) );
  OR2X1 P2_sub_1031_U26 ( .IN2(P2_sub_1031_n32), .IN1(P2_sub_1031_n31), 
        .Q(P2_sub_1031_n30) );
  NAND2X0 P2_sub_1031_U25 ( .IN1(P2_sub_1031_n29), .IN2(P2_sub_1031_n30), 
        .QN(P2_N4868) );
  NAND2X0 P2_sub_1031_U24 ( .IN1(n6651), .IN2(n6753), .QN(P2_sub_1031_n26) );
  OR2X1 P2_sub_1031_U23 ( .IN2(n6651), .IN1(n6753), .Q(P2_sub_1031_n27) );
  NAND2X0 P2_sub_1031_U22 ( .IN1(P2_sub_1031_n26), .IN2(P2_sub_1031_n27), 
        .QN(P2_sub_1031_n24) );
  NAND2X0 P2_sub_1031_U21 ( .IN1(P2_sub_1031_n24), .IN2(P2_sub_1031_n25), 
        .QN(P2_sub_1031_n22) );
  OR2X1 P2_sub_1031_U20 ( .IN2(P2_sub_1031_n25), .IN1(P2_sub_1031_n24), 
        .Q(P2_sub_1031_n23) );
  NAND2X0 P2_sub_1031_U19 ( .IN1(P2_sub_1031_n22), .IN2(P2_sub_1031_n23), 
        .QN(P2_N4869) );
  NAND2X0 P2_sub_1031_U18 ( .IN1(n6652), .IN2(n6748), .QN(P2_sub_1031_n19) );
  OR2X1 P2_sub_1031_U17 ( .IN2(n6652), .IN1(n6748), .Q(P2_sub_1031_n20) );
  NAND2X0 P2_sub_1031_U16 ( .IN1(P2_sub_1031_n19), .IN2(P2_sub_1031_n20), 
        .QN(P2_sub_1031_n17) );
  NAND2X0 P2_sub_1031_U15 ( .IN1(P2_sub_1031_n17), .IN2(P2_sub_1031_n18), 
        .QN(P2_sub_1031_n15) );
  OR2X1 P2_sub_1031_U14 ( .IN2(P2_sub_1031_n18), .IN1(P2_sub_1031_n17), 
        .Q(P2_sub_1031_n16) );
  NAND2X0 P2_sub_1031_U13 ( .IN1(P2_sub_1031_n15), .IN2(P2_sub_1031_n16), 
        .QN(P2_N4870) );
  NAND2X0 P2_sub_1031_U12 ( .IN1(n6653), .IN2(n6752), .QN(P2_sub_1031_n12) );
  OR2X1 P2_sub_1031_U11 ( .IN2(n6653), .IN1(n6752), .Q(P2_sub_1031_n13) );
  NAND2X0 P2_sub_1031_U10 ( .IN1(P2_sub_1031_n12), .IN2(P2_sub_1031_n13), 
        .QN(P2_sub_1031_n10) );
  NAND2X0 P2_sub_1031_U9 ( .IN1(P2_sub_1031_n10), .IN2(P2_sub_1031_n11), 
        .QN(P2_sub_1031_n8) );
  OR2X1 P2_sub_1031_U8 ( .IN2(P2_sub_1031_n11), .IN1(P2_sub_1031_n10), 
        .Q(P2_sub_1031_n9) );
  NAND2X0 P2_sub_1031_U7 ( .IN1(P2_sub_1031_n8), .IN2(P2_sub_1031_n9), 
        .QN(P2_N4871) );
  NAND2X0 P2_sub_1031_U6 ( .IN1(n6654), .IN2(n6757), .QN(P2_sub_1031_n5) );
  OR2X1 P2_sub_1031_U5 ( .IN2(n6654), .IN1(n6757), .Q(P2_sub_1031_n6) );
  NAND2X0 P2_sub_1031_U4 ( .IN1(P2_sub_1031_n5), .IN2(P2_sub_1031_n6), 
        .QN(P2_sub_1031_n3) );
  NAND2X0 P2_sub_1031_U3 ( .IN1(P2_sub_1031_n3), .IN2(P2_sub_1031_n4), 
        .QN(P2_sub_1031_n1) );
  OR2X1 P2_sub_1031_U2 ( .IN2(P2_sub_1031_n4), .IN1(P2_sub_1031_n3), 
        .Q(P2_sub_1031_n2) );
  NAND2X0 P2_sub_1031_U1 ( .IN1(P2_sub_1031_n1), .IN2(P2_sub_1031_n2), 
        .QN(P2_N4872) );
  NAND2X0 P2_sub_1031_U172 ( .IN1(P2_sub_1031_n169), .IN2(P2_sub_1031_n170), 
        .QN(P2_sub_1031_n18) );
  NAND2X0 P2_sub_1031_U171 ( .IN1(n6652), .IN2(P2_sub_1031_n18), 
        .QN(P2_sub_1031_n166) );
  OR2X1 P2_sub_1031_U170 ( .IN2(n6652), .IN1(P2_sub_1031_n18), 
        .Q(P2_sub_1031_n168) );
  NAND2X0 P2_sub_1031_U168 ( .IN1(P2_sub_1031_n168), .IN2(n6748), 
        .QN(P2_sub_1031_n167) );
  NAND2X0 P2_sub_1031_U167 ( .IN1(P2_sub_1031_n166), .IN2(P2_sub_1031_n167), 
        .QN(P2_sub_1031_n11) );
  NAND2X0 P2_sub_1031_U166 ( .IN1(n6653), .IN2(P2_sub_1031_n11), 
        .QN(P2_sub_1031_n163) );
  OR2X1 P2_sub_1031_U165 ( .IN2(n6653), .IN1(P2_sub_1031_n11), 
        .Q(P2_sub_1031_n165) );
  NAND2X0 P2_sub_1031_U163 ( .IN1(P2_sub_1031_n165), .IN2(n6752), 
        .QN(P2_sub_1031_n164) );
  NAND2X0 P2_sub_1031_U162 ( .IN1(P2_sub_1031_n163), .IN2(P2_sub_1031_n164), 
        .QN(P2_sub_1031_n4) );
  NAND2X0 P2_sub_1031_U161 ( .IN1(n6654), .IN2(P2_sub_1031_n4), 
        .QN(P2_sub_1031_n160) );
  OR2X1 P2_sub_1031_U160 ( .IN2(n6654), .IN1(P2_sub_1031_n4), 
        .Q(P2_sub_1031_n162) );
  NAND2X0 P2_sub_1031_U158 ( .IN1(P2_sub_1031_n162), .IN2(n6757), 
        .QN(P2_sub_1031_n161) );
  NAND2X0 P2_sub_1031_U157 ( .IN1(P2_sub_1031_n160), .IN2(P2_sub_1031_n161), 
        .QN(P2_sub_1031_n154) );
  NAND2X0 P2_sub_1031_U156 ( .IN1(P2_sub_1031_n159), .IN2(P2_sub_1031_n154), 
        .QN(P2_sub_1031_n157) );
  OR2X1 P2_sub_1031_U155 ( .IN2(P2_sub_1031_n154), .IN1(P2_sub_1031_n159), 
        .Q(P2_sub_1031_n158) );
  NAND2X0 P2_sub_1031_U154 ( .IN1(P2_sub_1031_n157), .IN2(P2_sub_1031_n158), 
        .QN(P2_N4873) );
  NAND2X0 P2_sub_1031_U152 ( .IN1(n6656), .IN2(n6756), .QN(P2_sub_1031_n155)
         );
  OR2X1 P2_sub_1031_U151 ( .IN2(n6656), .IN1(n6756), .Q(P2_sub_1031_n156) );
  NAND2X0 P2_sub_1031_U150 ( .IN1(P2_sub_1031_n155), .IN2(P2_sub_1031_n156), 
        .QN(P2_sub_1031_n149) );
  NAND2X0 P2_sub_1031_U149 ( .IN1(n6655), .IN2(P2_sub_1031_n154), 
        .QN(P2_sub_1031_n150) );
  OR2X1 P2_sub_1031_U148 ( .IN2(n6655), .IN1(P2_sub_1031_n154), 
        .Q(P2_sub_1031_n152) );
  NAND2X0 P2_sub_1031_U147 ( .IN1(P2_sub_1031_n152), .IN2(n6760), 
        .QN(P2_sub_1031_n151) );
  NAND2X0 P2_sub_1031_U146 ( .IN1(P2_sub_1031_n150), .IN2(P2_sub_1031_n151), 
        .QN(P2_sub_1031_n144) );
  NAND2X0 P2_sub_1031_U145 ( .IN1(P2_sub_1031_n149), .IN2(P2_sub_1031_n144), 
        .QN(P2_sub_1031_n147) );
  OR2X1 P2_sub_1031_U144 ( .IN2(P2_sub_1031_n144), .IN1(P2_sub_1031_n149), 
        .Q(P2_sub_1031_n148) );
  NAND2X0 P2_sub_1031_U143 ( .IN1(P2_sub_1031_n147), .IN2(P2_sub_1031_n148), 
        .QN(P2_N4874) );
  NAND2X0 P2_sub_1031_U141 ( .IN1(n6657), .IN2(n6761), .QN(P2_sub_1031_n145)
         );
  OR2X1 P2_sub_1031_U140 ( .IN2(n6657), .IN1(n6761), .Q(P2_sub_1031_n146) );
  NAND2X0 P2_sub_1031_U139 ( .IN1(P2_sub_1031_n145), .IN2(P2_sub_1031_n146), 
        .QN(P2_sub_1031_n139) );
  NAND2X0 P2_sub_1031_U138 ( .IN1(n6656), .IN2(P2_sub_1031_n144), 
        .QN(P2_sub_1031_n140) );
  OR2X1 P2_sub_1031_U137 ( .IN2(n6656), .IN1(P2_sub_1031_n144), 
        .Q(P2_sub_1031_n142) );
  NAND2X0 P2_sub_1031_U136 ( .IN1(P2_sub_1031_n142), .IN2(n6756), 
        .QN(P2_sub_1031_n141) );
  NAND2X0 P2_sub_1031_U135 ( .IN1(P2_sub_1031_n140), .IN2(P2_sub_1031_n141), 
        .QN(P2_sub_1031_n134) );
  NAND2X0 P2_sub_1031_U134 ( .IN1(P2_sub_1031_n139), .IN2(P2_sub_1031_n134), 
        .QN(P2_sub_1031_n137) );
  OR2X1 P2_sub_1031_U133 ( .IN2(P2_sub_1031_n134), .IN1(P2_sub_1031_n139), 
        .Q(P2_sub_1031_n138) );
  NAND2X0 P2_sub_1031_U132 ( .IN1(P2_sub_1031_n137), .IN2(P2_sub_1031_n138), 
        .QN(P2_N4875) );
  NAND2X0 P2_sub_1031_U130 ( .IN1(n6658), .IN2(n6765), .QN(P2_sub_1031_n135)
         );
  OR2X1 P2_sub_1031_U129 ( .IN2(n6658), .IN1(n6765), .Q(P2_sub_1031_n136) );
  NAND2X0 P2_sub_1031_U128 ( .IN1(P2_sub_1031_n135), .IN2(P2_sub_1031_n136), 
        .QN(P2_sub_1031_n129) );
  NAND2X0 P2_sub_1031_U127 ( .IN1(n6657), .IN2(P2_sub_1031_n134), 
        .QN(P2_sub_1031_n130) );
  OR2X1 P2_sub_1031_U126 ( .IN2(n6657), .IN1(P2_sub_1031_n134), 
        .Q(P2_sub_1031_n132) );
  NAND2X0 P2_sub_1031_U125 ( .IN1(P2_sub_1031_n132), .IN2(n6761), 
        .QN(P2_sub_1031_n131) );
  NAND2X0 P2_sub_1031_U124 ( .IN1(P2_sub_1031_n130), .IN2(P2_sub_1031_n131), 
        .QN(P2_sub_1031_n124) );
  NAND2X0 P2_sub_1031_U123 ( .IN1(P2_sub_1031_n129), .IN2(P2_sub_1031_n124), 
        .QN(P2_sub_1031_n127) );
  OR2X1 P2_sub_1031_U122 ( .IN2(P2_sub_1031_n124), .IN1(P2_sub_1031_n129), 
        .Q(P2_sub_1031_n128) );
  NAND2X0 P2_sub_1031_U121 ( .IN1(P2_sub_1031_n127), .IN2(P2_sub_1031_n128), 
        .QN(P2_N4876) );
  NAND2X0 P2_sub_1031_U119 ( .IN1(n6659), .IN2(n6769), .QN(P2_sub_1031_n125)
         );
  OR2X1 P2_sub_1031_U118 ( .IN2(n6659), .IN1(n6769), .Q(P2_sub_1031_n126) );
  NAND2X0 P2_sub_1031_U117 ( .IN1(P2_sub_1031_n125), .IN2(P2_sub_1031_n126), 
        .QN(P2_sub_1031_n119) );
  NAND2X0 P2_sub_1031_U116 ( .IN1(n6658), .IN2(P2_sub_1031_n124), 
        .QN(P2_sub_1031_n120) );
  OR2X1 P2_sub_1031_U115 ( .IN2(n6658), .IN1(P2_sub_1031_n124), 
        .Q(P2_sub_1031_n122) );
  NAND2X0 P2_sub_1031_U114 ( .IN1(P2_sub_1031_n122), .IN2(n6765), 
        .QN(P2_sub_1031_n121) );
  NAND2X0 P2_sub_1031_U113 ( .IN1(P2_sub_1031_n120), .IN2(P2_sub_1031_n121), 
        .QN(P2_sub_1031_n114) );
  NAND2X0 P2_sub_1031_U112 ( .IN1(P2_sub_1031_n119), .IN2(P2_sub_1031_n114), 
        .QN(P2_sub_1031_n117) );
  OR2X1 P2_sub_1031_U111 ( .IN2(P2_sub_1031_n114), .IN1(P2_sub_1031_n119), 
        .Q(P2_sub_1031_n118) );
  NAND2X0 P2_sub_1031_U110 ( .IN1(P2_sub_1031_n117), .IN2(P2_sub_1031_n118), 
        .QN(P2_N4877) );
  NAND2X0 P2_sub_1031_U108 ( .IN1(n6660), .IN2(n6764), .QN(P2_sub_1031_n115)
         );
  OR2X1 P2_sub_1031_U107 ( .IN2(n6660), .IN1(n6764), .Q(P2_sub_1031_n116) );
  NAND2X0 P2_sub_1031_U106 ( .IN1(P2_sub_1031_n115), .IN2(P2_sub_1031_n116), 
        .QN(P2_sub_1031_n109) );
  NAND2X0 P2_sub_1031_U105 ( .IN1(n6659), .IN2(P2_sub_1031_n114), 
        .QN(P2_sub_1031_n110) );
  OR2X1 P2_sub_1031_U104 ( .IN2(n6659), .IN1(P2_sub_1031_n114), 
        .Q(P2_sub_1031_n112) );
  NAND2X0 P2_sub_1031_U103 ( .IN1(P2_sub_1031_n112), .IN2(n6769), 
        .QN(P2_sub_1031_n111) );
  NAND2X0 P2_sub_1031_U102 ( .IN1(P2_sub_1031_n110), .IN2(P2_sub_1031_n111), 
        .QN(P2_sub_1031_n104) );
  NAND2X0 P2_sub_1031_U101 ( .IN1(P2_sub_1031_n109), .IN2(P2_sub_1031_n104), 
        .QN(P2_sub_1031_n107) );
  OR2X1 P2_sub_1031_U100 ( .IN2(P2_sub_1031_n104), .IN1(P2_sub_1031_n109), 
        .Q(P2_sub_1031_n108) );
  NAND2X0 P2_sub_1031_U99 ( .IN1(P2_sub_1031_n107), .IN2(P2_sub_1031_n108), 
        .QN(P2_N4878) );
  NAND2X0 P2_sub_1031_U97 ( .IN1(n6661), .IN2(n6768), .QN(P2_sub_1031_n105) );
  OR2X1 P2_sub_1031_U96 ( .IN2(n6661), .IN1(n6768), .Q(P2_sub_1031_n106) );
  NAND2X0 P2_sub_1031_U95 ( .IN1(P2_sub_1031_n105), .IN2(P2_sub_1031_n106), 
        .QN(P2_sub_1031_n99) );
  NAND2X0 P2_sub_1031_U94 ( .IN1(n6660), .IN2(P2_sub_1031_n104), 
        .QN(P2_sub_1031_n100) );
  OR2X1 P2_sub_1031_U93 ( .IN2(n6660), .IN1(P2_sub_1031_n104), 
        .Q(P2_sub_1031_n102) );
  NAND2X0 P2_sub_1031_U92 ( .IN1(P2_sub_1031_n102), .IN2(n6764), 
        .QN(P2_sub_1031_n101) );
  NAND2X0 P2_sub_1031_U91 ( .IN1(P2_sub_1031_n100), .IN2(P2_sub_1031_n101), 
        .QN(P2_sub_1031_n94) );
  NAND2X0 P2_sub_1031_U90 ( .IN1(P2_sub_1031_n99), .IN2(P2_sub_1031_n94), 
        .QN(P2_sub_1031_n97) );
  OR2X1 P2_sub_1031_U89 ( .IN2(P2_sub_1031_n94), .IN1(P2_sub_1031_n99), 
        .Q(P2_sub_1031_n98) );
  NAND2X0 P2_sub_1031_U88 ( .IN1(P2_sub_1031_n97), .IN2(P2_sub_1031_n98), 
        .QN(P2_N4879) );
  NAND2X0 P2_sub_1031_U86 ( .IN1(n6662), .IN2(n6772), .QN(P2_sub_1031_n95) );
  OR2X1 P2_sub_1031_U85 ( .IN2(n6662), .IN1(n6772), .Q(P2_sub_1031_n96) );
  NAND2X0 P2_sub_1031_U84 ( .IN1(P2_sub_1031_n95), .IN2(P2_sub_1031_n96), 
        .QN(P2_sub_1031_n89) );
  NAND2X0 P2_sub_1031_U83 ( .IN1(n6661), .IN2(P2_sub_1031_n94), 
        .QN(P2_sub_1031_n90) );
  OR2X1 P2_sub_1031_U82 ( .IN2(n6661), .IN1(P2_sub_1031_n94), 
        .Q(P2_sub_1031_n92) );
  NAND2X0 P2_sub_1031_U81 ( .IN1(P2_sub_1031_n92), .IN2(n6768), 
        .QN(P2_sub_1031_n91) );
  NAND2X0 P2_sub_1031_U80 ( .IN1(P2_sub_1031_n90), .IN2(P2_sub_1031_n91), 
        .QN(P2_sub_1031_n84) );
  NOR2X0 P2_sub_1031_U210 ( .QN(P2_sub_1031_n187), .IN1(n6731), .IN2(n9842) );
  INVX0 P2_sub_1031_U209 ( .ZN(P2_sub_1031_n60), .INP(P2_sub_1031_n187) );
  NAND2X0 P2_sub_1031_U208 ( .IN1(n9842), .IN2(n6731), .QN(P2_sub_1031_n190)
         );
  NAND2X0 P2_sub_1031_U207 ( .IN1(P2_sub_1031_n60), .IN2(P2_sub_1031_n190), 
        .QN(P2_N4863) );
  NAND2X0 P2_sub_1031_U205 ( .IN1(n6655), .IN2(n6760), .QN(P2_sub_1031_n188)
         );
  OR2X1 P2_sub_1031_U204 ( .IN2(n6655), .IN1(n6760), .Q(P2_sub_1031_n189) );
  NAND2X0 P2_sub_1031_U203 ( .IN1(P2_sub_1031_n188), .IN2(P2_sub_1031_n189), 
        .QN(P2_sub_1031_n159) );
  NAND2X0 P2_sub_1031_U202 ( .IN1(n6720), .IN2(P2_sub_1031_n60), 
        .QN(P2_sub_1031_n184) );
  NAND2X0 P2_sub_1031_U200 ( .IN1(P2_sub_1031_n187), .IN2(n18997), 
        .QN(P2_sub_1031_n186) );
  NAND2X0 P2_sub_1031_U198 ( .IN1(P2_sub_1031_n186), .IN2(n6733), 
        .QN(P2_sub_1031_n185) );
  NAND2X0 P2_sub_1031_U197 ( .IN1(P2_sub_1031_n184), .IN2(P2_sub_1031_n185), 
        .QN(P2_sub_1031_n53) );
  NAND2X0 P2_sub_1031_U196 ( .IN1(n6721), .IN2(P2_sub_1031_n53), 
        .QN(P2_sub_1031_n181) );
  OR2X1 P2_sub_1031_U195 ( .IN2(n6721), .IN1(P2_sub_1031_n53), 
        .Q(P2_sub_1031_n183) );
  NAND2X0 P2_sub_1031_U193 ( .IN1(P2_sub_1031_n183), .IN2(n6735), 
        .QN(P2_sub_1031_n182) );
  NAND2X0 P2_sub_1031_U192 ( .IN1(P2_sub_1031_n181), .IN2(P2_sub_1031_n182), 
        .QN(P2_sub_1031_n46) );
  NAND2X0 P2_sub_1031_U191 ( .IN1(n6648), .IN2(P2_sub_1031_n46), 
        .QN(P2_sub_1031_n178) );
  OR2X1 P2_sub_1031_U190 ( .IN2(n6648), .IN1(P2_sub_1031_n46), 
        .Q(P2_sub_1031_n180) );
  NAND2X0 P2_sub_1031_U188 ( .IN1(P2_sub_1031_n180), .IN2(n6743), 
        .QN(P2_sub_1031_n179) );
  NAND2X0 P2_sub_1031_U187 ( .IN1(P2_sub_1031_n178), .IN2(P2_sub_1031_n179), 
        .QN(P2_sub_1031_n39) );
  NAND2X0 P2_sub_1031_U186 ( .IN1(n6649), .IN2(P2_sub_1031_n39), 
        .QN(P2_sub_1031_n175) );
  OR2X1 P2_sub_1031_U185 ( .IN2(n6649), .IN1(P2_sub_1031_n39), 
        .Q(P2_sub_1031_n177) );
  NAND2X0 P2_sub_1031_U183 ( .IN1(P2_sub_1031_n177), .IN2(n6745), 
        .QN(P2_sub_1031_n176) );
  NAND2X0 P2_sub_1031_U182 ( .IN1(P2_sub_1031_n175), .IN2(P2_sub_1031_n176), 
        .QN(P2_sub_1031_n32) );
  NAND2X0 P2_sub_1031_U181 ( .IN1(n6650), .IN2(P2_sub_1031_n32), 
        .QN(P2_sub_1031_n172) );
  OR2X1 P2_sub_1031_U180 ( .IN2(n6650), .IN1(P2_sub_1031_n32), 
        .Q(P2_sub_1031_n174) );
  NAND2X0 P2_sub_1031_U178 ( .IN1(P2_sub_1031_n174), .IN2(n6749), 
        .QN(P2_sub_1031_n173) );
  NAND2X0 P2_sub_1031_U177 ( .IN1(P2_sub_1031_n172), .IN2(P2_sub_1031_n173), 
        .QN(P2_sub_1031_n25) );
  NAND2X0 P2_sub_1031_U176 ( .IN1(n6651), .IN2(P2_sub_1031_n25), 
        .QN(P2_sub_1031_n169) );
  OR2X1 P2_sub_1031_U175 ( .IN2(n6651), .IN1(P2_sub_1031_n25), 
        .Q(P2_sub_1031_n171) );
  NAND2X0 P2_sub_1031_U173 ( .IN1(P2_sub_1031_n171), .IN2(n6753), 
        .QN(P2_sub_1031_n170) );
  NOR2X0 P2_lt_688_U50 ( .QN(P2_lt_688_n62), .IN1(P2_N5025), 
        .IN2(P2_lt_688_n63) );
  NOR2X0 P2_lt_688_U49 ( .QN(P2_lt_688_n59), .IN1(P2_lt_688_n61), 
        .IN2(P2_lt_688_n62) );
  INVX0 P2_lt_688_U48 ( .ZN(P2_lt_688_n58), .INP(P2_N5341) );
  OR2X1 P2_lt_688_U47 ( .IN2(P2_N5026), .IN1(P2_lt_688_n58), .Q(P2_lt_688_n60)
         );
  NAND2X0 P2_lt_688_U46 ( .IN1(P2_lt_688_n59), .IN2(P2_lt_688_n60), 
        .QN(P2_lt_688_n56) );
  NAND2X0 P2_lt_688_U45 ( .IN1(P2_N5026), .IN2(P2_lt_688_n58), 
        .QN(P2_lt_688_n57) );
  NAND2X0 P2_lt_688_U44 ( .IN1(P2_lt_688_n56), .IN2(P2_lt_688_n57), 
        .QN(P2_lt_688_n55) );
  NOR2X0 P2_lt_688_U43 ( .QN(P2_lt_688_n51), .IN1(P2_lt_688_n54), 
        .IN2(P2_lt_688_n55) );
  NOR2X0 P2_lt_688_U42 ( .QN(P2_lt_688_n52), .IN1(P2_N5027), 
        .IN2(P2_lt_688_n53) );
  NOR2X0 P2_lt_688_U41 ( .QN(P2_lt_688_n49), .IN1(P2_lt_688_n51), 
        .IN2(P2_lt_688_n52) );
  INVX0 P2_lt_688_U40 ( .ZN(P2_lt_688_n48), .INP(P2_N5343) );
  OR2X1 P2_lt_688_U39 ( .IN2(P2_N5028), .IN1(P2_lt_688_n48), .Q(P2_lt_688_n50)
         );
  NAND2X0 P2_lt_688_U38 ( .IN1(P2_lt_688_n49), .IN2(P2_lt_688_n50), 
        .QN(P2_lt_688_n46) );
  NAND2X0 P2_lt_688_U37 ( .IN1(P2_N5028), .IN2(P2_lt_688_n48), 
        .QN(P2_lt_688_n47) );
  NAND2X0 P2_lt_688_U36 ( .IN1(P2_lt_688_n46), .IN2(P2_lt_688_n47), 
        .QN(P2_lt_688_n45) );
  NOR2X0 P2_lt_688_U35 ( .QN(P2_lt_688_n41), .IN1(P2_lt_688_n44), 
        .IN2(P2_lt_688_n45) );
  NOR2X0 P2_lt_688_U34 ( .QN(P2_lt_688_n42), .IN1(P2_N5029), 
        .IN2(P2_lt_688_n43) );
  NOR2X0 P2_lt_688_U33 ( .QN(P2_lt_688_n39), .IN1(P2_lt_688_n41), 
        .IN2(P2_lt_688_n42) );
  INVX0 P2_lt_688_U32 ( .ZN(P2_lt_688_n38), .INP(P2_N5345) );
  OR2X1 P2_lt_688_U31 ( .IN2(P2_N5030), .IN1(P2_lt_688_n38), .Q(P2_lt_688_n40)
         );
  NAND2X0 P2_lt_688_U30 ( .IN1(P2_lt_688_n39), .IN2(P2_lt_688_n40), 
        .QN(P2_lt_688_n36) );
  NAND2X0 P2_lt_688_U29 ( .IN1(P2_N5030), .IN2(P2_lt_688_n38), 
        .QN(P2_lt_688_n37) );
  NAND2X0 P2_lt_688_U28 ( .IN1(P2_lt_688_n36), .IN2(P2_lt_688_n37), 
        .QN(P2_lt_688_n35) );
  NOR2X0 P2_lt_688_U27 ( .QN(P2_lt_688_n31), .IN1(P2_lt_688_n34), 
        .IN2(P2_lt_688_n35) );
  NOR2X0 P2_lt_688_U26 ( .QN(P2_lt_688_n32), .IN1(P2_N5031), 
        .IN2(P2_lt_688_n33) );
  NOR2X0 P2_lt_688_U25 ( .QN(P2_lt_688_n29), .IN1(P2_lt_688_n31), 
        .IN2(P2_lt_688_n32) );
  INVX0 P2_lt_688_U24 ( .ZN(P2_lt_688_n28), .INP(P2_N5347) );
  OR2X1 P2_lt_688_U23 ( .IN2(P2_N5032), .IN1(P2_lt_688_n28), .Q(P2_lt_688_n30)
         );
  NAND2X0 P2_lt_688_U22 ( .IN1(P2_lt_688_n29), .IN2(P2_lt_688_n30), 
        .QN(P2_lt_688_n26) );
  NAND2X0 P2_lt_688_U21 ( .IN1(P2_N5032), .IN2(P2_lt_688_n28), 
        .QN(P2_lt_688_n27) );
  NAND2X0 P2_lt_688_U20 ( .IN1(P2_lt_688_n26), .IN2(P2_lt_688_n27), 
        .QN(P2_lt_688_n25) );
  NOR2X0 P2_lt_688_U19 ( .QN(P2_lt_688_n21), .IN1(P2_lt_688_n24), 
        .IN2(P2_lt_688_n25) );
  NOR2X0 P2_lt_688_U18 ( .QN(P2_lt_688_n22), .IN1(P2_N5033), 
        .IN2(P2_lt_688_n23) );
  NOR2X0 P2_lt_688_U17 ( .QN(P2_lt_688_n19), .IN1(P2_lt_688_n21), 
        .IN2(P2_lt_688_n22) );
  INVX0 P2_lt_688_U16 ( .ZN(P2_lt_688_n18), .INP(P2_N5349) );
  OR2X1 P2_lt_688_U15 ( .IN2(P2_N5034), .IN1(P2_lt_688_n18), .Q(P2_lt_688_n20)
         );
  NAND2X0 P2_lt_688_U14 ( .IN1(P2_lt_688_n19), .IN2(P2_lt_688_n20), 
        .QN(P2_lt_688_n16) );
  NAND2X0 P2_lt_688_U13 ( .IN1(P2_N5034), .IN2(P2_lt_688_n18), 
        .QN(P2_lt_688_n17) );
  NAND2X0 P2_lt_688_U12 ( .IN1(P2_lt_688_n16), .IN2(P2_lt_688_n17), 
        .QN(P2_lt_688_n15) );
  NOR2X0 P2_lt_688_U11 ( .QN(P2_lt_688_n11), .IN1(P2_lt_688_n14), 
        .IN2(P2_lt_688_n15) );
  NOR2X0 P2_lt_688_U10 ( .QN(P2_lt_688_n12), .IN1(P2_N5035), 
        .IN2(P2_lt_688_n13) );
  NOR2X0 P2_lt_688_U9 ( .QN(P2_lt_688_n9), .IN1(P2_lt_688_n11), 
        .IN2(P2_lt_688_n12) );
  INVX0 P2_lt_688_U8 ( .ZN(P2_lt_688_n8), .INP(P2_N5351) );
  OR2X1 P2_lt_688_U7 ( .IN2(P2_N5036), .IN1(P2_lt_688_n8), .Q(P2_lt_688_n10)
         );
  NAND2X0 P2_lt_688_U6 ( .IN1(P2_lt_688_n9), .IN2(P2_lt_688_n10), 
        .QN(P2_lt_688_n6) );
  NAND2X0 P2_lt_688_U5 ( .IN1(P2_N5036), .IN2(P2_lt_688_n8), .QN(P2_lt_688_n7)
         );
  NAND2X0 P2_lt_688_U4 ( .IN1(P2_lt_688_n6), .IN2(P2_lt_688_n7), 
        .QN(P2_lt_688_n3) );
  NAND2X0 P2_lt_688_U3 ( .IN1(P2_N5037), .IN2(P2_lt_688_n5), .QN(P2_lt_688_n4)
         );
  NAND2X0 P2_lt_688_U2 ( .IN1(P2_lt_688_n3), .IN2(P2_lt_688_n4), 
        .QN(P2_lt_688_n2) );
  NAND2X0 P2_lt_688_U1 ( .IN1(P2_lt_688_n1), .IN2(P2_lt_688_n2), .QN(P2_N5135)
         );
  INVX0 P2_lt_688_U143 ( .ZN(P2_lt_688_n73), .INP(P2_N5338) );
  AND2X1 P2_lt_688_U142 ( .IN1(P2_lt_688_n73), .IN2(P2_N5023), 
        .Q(P2_lt_688_n74) );
  INVX0 P2_lt_688_U141 ( .ZN(P2_lt_688_n83), .INP(P2_N5336) );
  AND2X1 P2_lt_688_U140 ( .IN1(P2_lt_688_n83), .IN2(P2_N5021), 
        .Q(P2_lt_688_n84) );
  INVX0 P2_lt_688_U139 ( .ZN(P2_lt_688_n93), .INP(P2_N5334) );
  AND2X1 P2_lt_688_U138 ( .IN1(P2_lt_688_n93), .IN2(P2_N5019), 
        .Q(P2_lt_688_n94) );
  INVX0 P2_lt_688_U137 ( .ZN(P2_lt_688_n103), .INP(P2_N5332) );
  AND2X1 P2_lt_688_U136 ( .IN1(P2_lt_688_n103), .IN2(P2_N5017), 
        .Q(P2_lt_688_n104) );
  NOR2X0 P2_lt_688_U134 ( .QN(P2_lt_688_n114), .IN1(P2_N5330), .IN2(n7275) );
  INVX0 P2_lt_688_U133 ( .ZN(P2_lt_688_n123), .INP(P2_N5328) );
  AND2X1 P2_lt_688_U132 ( .IN1(P2_lt_688_n123), .IN2(P2_N5013), 
        .Q(P2_lt_688_n124) );
  INVX0 P2_lt_688_U131 ( .ZN(P2_lt_688_n133), .INP(P2_N5326) );
  AND2X1 P2_lt_688_U130 ( .IN1(P2_lt_688_n133), .IN2(P2_N5011), 
        .Q(P2_lt_688_n134) );
  INVX0 P2_lt_688_U129 ( .ZN(P2_lt_688_n143), .INP(P2_N5324) );
  AND2X1 P2_lt_688_U128 ( .IN1(P2_lt_688_n143), .IN2(P2_N5009), 
        .Q(P2_lt_688_n144) );
  INVX0 P2_lt_688_U127 ( .ZN(P2_lt_688_n154), .INP(P2_N5322) );
  INVX0 P2_lt_688_U126 ( .ZN(P2_lt_688_n156), .INP(P2_N5006) );
  NOR2X0 P2_lt_688_U125 ( .QN(P2_lt_688_n153), .IN1(P2_lt_688_n156), 
        .IN2(P2_N5321) );
  AND2X1 P2_lt_688_U124 ( .IN1(P2_lt_688_n154), .IN2(P2_lt_688_n153), 
        .Q(P2_lt_688_n155) );
  NOR2X0 P2_lt_688_U123 ( .QN(P2_lt_688_n151), .IN1(P2_N5007), 
        .IN2(P2_lt_688_n155) );
  NOR2X0 P2_lt_688_U122 ( .QN(P2_lt_688_n152), .IN1(P2_lt_688_n153), 
        .IN2(P2_lt_688_n154) );
  NOR2X0 P2_lt_688_U121 ( .QN(P2_lt_688_n149), .IN1(P2_lt_688_n151), 
        .IN2(P2_lt_688_n152) );
  INVX0 P2_lt_688_U120 ( .ZN(P2_lt_688_n148), .INP(P2_N5323) );
  OR2X1 P2_lt_688_U119 ( .IN2(P2_N5008), .IN1(P2_lt_688_n148), 
        .Q(P2_lt_688_n150) );
  NAND2X0 P2_lt_688_U118 ( .IN1(P2_lt_688_n149), .IN2(P2_lt_688_n150), 
        .QN(P2_lt_688_n146) );
  NAND2X0 P2_lt_688_U117 ( .IN1(P2_N5008), .IN2(P2_lt_688_n148), 
        .QN(P2_lt_688_n147) );
  NAND2X0 P2_lt_688_U116 ( .IN1(P2_lt_688_n146), .IN2(P2_lt_688_n147), 
        .QN(P2_lt_688_n145) );
  NOR2X0 P2_lt_688_U115 ( .QN(P2_lt_688_n141), .IN1(P2_lt_688_n144), 
        .IN2(P2_lt_688_n145) );
  NOR2X0 P2_lt_688_U114 ( .QN(P2_lt_688_n142), .IN1(P2_N5009), 
        .IN2(P2_lt_688_n143) );
  NOR2X0 P2_lt_688_U113 ( .QN(P2_lt_688_n139), .IN1(P2_lt_688_n141), 
        .IN2(P2_lt_688_n142) );
  INVX0 P2_lt_688_U112 ( .ZN(P2_lt_688_n138), .INP(P2_N5325) );
  OR2X1 P2_lt_688_U111 ( .IN2(P2_N5010), .IN1(P2_lt_688_n138), 
        .Q(P2_lt_688_n140) );
  NAND2X0 P2_lt_688_U110 ( .IN1(P2_lt_688_n139), .IN2(P2_lt_688_n140), 
        .QN(P2_lt_688_n136) );
  NAND2X0 P2_lt_688_U109 ( .IN1(P2_N5010), .IN2(P2_lt_688_n138), 
        .QN(P2_lt_688_n137) );
  NAND2X0 P2_lt_688_U108 ( .IN1(P2_lt_688_n136), .IN2(P2_lt_688_n137), 
        .QN(P2_lt_688_n135) );
  NOR2X0 P2_lt_688_U107 ( .QN(P2_lt_688_n131), .IN1(P2_lt_688_n134), 
        .IN2(P2_lt_688_n135) );
  NOR2X0 P2_lt_688_U106 ( .QN(P2_lt_688_n132), .IN1(P2_N5011), 
        .IN2(P2_lt_688_n133) );
  NOR2X0 P2_lt_688_U105 ( .QN(P2_lt_688_n129), .IN1(P2_lt_688_n131), 
        .IN2(P2_lt_688_n132) );
  INVX0 P2_lt_688_U104 ( .ZN(P2_lt_688_n128), .INP(P2_N5327) );
  OR2X1 P2_lt_688_U103 ( .IN2(P2_N5012), .IN1(P2_lt_688_n128), 
        .Q(P2_lt_688_n130) );
  NAND2X0 P2_lt_688_U102 ( .IN1(P2_lt_688_n129), .IN2(P2_lt_688_n130), 
        .QN(P2_lt_688_n126) );
  NAND2X0 P2_lt_688_U101 ( .IN1(P2_N5012), .IN2(P2_lt_688_n128), 
        .QN(P2_lt_688_n127) );
  NAND2X0 P2_lt_688_U100 ( .IN1(P2_lt_688_n126), .IN2(P2_lt_688_n127), 
        .QN(P2_lt_688_n125) );
  NOR2X0 P2_lt_688_U99 ( .QN(P2_lt_688_n121), .IN1(P2_lt_688_n124), 
        .IN2(P2_lt_688_n125) );
  NOR2X0 P2_lt_688_U98 ( .QN(P2_lt_688_n122), .IN1(P2_N5013), 
        .IN2(P2_lt_688_n123) );
  NOR2X0 P2_lt_688_U97 ( .QN(P2_lt_688_n119), .IN1(P2_lt_688_n121), 
        .IN2(P2_lt_688_n122) );
  INVX0 P2_lt_688_U96 ( .ZN(P2_lt_688_n118), .INP(P2_N5329) );
  OR2X1 P2_lt_688_U95 ( .IN2(P2_N5014), .IN1(P2_lt_688_n118), 
        .Q(P2_lt_688_n120) );
  NAND2X0 P2_lt_688_U94 ( .IN1(P2_lt_688_n119), .IN2(P2_lt_688_n120), 
        .QN(P2_lt_688_n116) );
  NAND2X0 P2_lt_688_U93 ( .IN1(P2_N5014), .IN2(P2_lt_688_n118), 
        .QN(P2_lt_688_n117) );
  NAND2X0 P2_lt_688_U92 ( .IN1(P2_lt_688_n116), .IN2(P2_lt_688_n117), 
        .QN(P2_lt_688_n115) );
  NOR2X0 P2_lt_688_U91 ( .QN(P2_lt_688_n112), .IN1(P2_lt_688_n114), 
        .IN2(P2_lt_688_n115) );
  INVX0 P2_lt_688_U90 ( .ZN(P2_lt_688_n108), .INP(P2_N5331) );
  NOR2X0 P2_lt_688_U89 ( .QN(P2_lt_688_n113), .IN1(P2_N5016), 
        .IN2(P2_lt_688_n108) );
  NOR2X0 P2_lt_688_U88 ( .QN(P2_lt_688_n109), .IN1(P2_lt_688_n112), 
        .IN2(P2_lt_688_n113) );
  NAND2X0 P2_lt_688_U87 ( .IN1(P2_N5330), .IN2(n7275), .QN(P2_lt_688_n110) );
  NAND2X0 P2_lt_688_U86 ( .IN1(P2_lt_688_n109), .IN2(P2_lt_688_n110), 
        .QN(P2_lt_688_n106) );
  NAND2X0 P2_lt_688_U85 ( .IN1(P2_N5016), .IN2(P2_lt_688_n108), 
        .QN(P2_lt_688_n107) );
  NAND2X0 P2_lt_688_U84 ( .IN1(P2_lt_688_n106), .IN2(P2_lt_688_n107), 
        .QN(P2_lt_688_n105) );
  NOR2X0 P2_lt_688_U83 ( .QN(P2_lt_688_n101), .IN1(P2_lt_688_n104), 
        .IN2(P2_lt_688_n105) );
  NOR2X0 P2_lt_688_U82 ( .QN(P2_lt_688_n102), .IN1(P2_N5017), 
        .IN2(P2_lt_688_n103) );
  NOR2X0 P2_lt_688_U81 ( .QN(P2_lt_688_n99), .IN1(P2_lt_688_n101), 
        .IN2(P2_lt_688_n102) );
  INVX0 P2_lt_688_U80 ( .ZN(P2_lt_688_n98), .INP(P2_N5333) );
  OR2X1 P2_lt_688_U79 ( .IN2(P2_N5018), .IN1(P2_lt_688_n98), 
        .Q(P2_lt_688_n100) );
  NAND2X0 P2_lt_688_U78 ( .IN1(P2_lt_688_n99), .IN2(P2_lt_688_n100), 
        .QN(P2_lt_688_n96) );
  NAND2X0 P2_lt_688_U77 ( .IN1(P2_N5018), .IN2(P2_lt_688_n98), 
        .QN(P2_lt_688_n97) );
  NAND2X0 P2_lt_688_U76 ( .IN1(P2_lt_688_n96), .IN2(P2_lt_688_n97), 
        .QN(P2_lt_688_n95) );
  NOR2X0 P2_lt_688_U75 ( .QN(P2_lt_688_n91), .IN1(P2_lt_688_n94), 
        .IN2(P2_lt_688_n95) );
  NOR2X0 P2_lt_688_U74 ( .QN(P2_lt_688_n92), .IN1(P2_N5019), 
        .IN2(P2_lt_688_n93) );
  NOR2X0 P2_lt_688_U73 ( .QN(P2_lt_688_n89), .IN1(P2_lt_688_n91), 
        .IN2(P2_lt_688_n92) );
  INVX0 P2_lt_688_U72 ( .ZN(P2_lt_688_n88), .INP(P2_N5335) );
  OR2X1 P2_lt_688_U71 ( .IN2(P2_N5020), .IN1(P2_lt_688_n88), .Q(P2_lt_688_n90)
         );
  NAND2X0 P2_lt_688_U70 ( .IN1(P2_lt_688_n89), .IN2(P2_lt_688_n90), 
        .QN(P2_lt_688_n86) );
  NAND2X0 P2_lt_688_U69 ( .IN1(P2_N5020), .IN2(P2_lt_688_n88), 
        .QN(P2_lt_688_n87) );
  NAND2X0 P2_lt_688_U68 ( .IN1(P2_lt_688_n86), .IN2(P2_lt_688_n87), 
        .QN(P2_lt_688_n85) );
  NOR2X0 P2_lt_688_U67 ( .QN(P2_lt_688_n81), .IN1(P2_lt_688_n84), 
        .IN2(P2_lt_688_n85) );
  NOR2X0 P2_lt_688_U66 ( .QN(P2_lt_688_n82), .IN1(P2_N5021), 
        .IN2(P2_lt_688_n83) );
  NOR2X0 P2_lt_688_U65 ( .QN(P2_lt_688_n79), .IN1(P2_lt_688_n81), 
        .IN2(P2_lt_688_n82) );
  INVX0 P2_lt_688_U64 ( .ZN(P2_lt_688_n78), .INP(P2_N5337) );
  OR2X1 P2_lt_688_U63 ( .IN2(P2_N5022), .IN1(P2_lt_688_n78), .Q(P2_lt_688_n80)
         );
  NAND2X0 P2_lt_688_U62 ( .IN1(P2_lt_688_n79), .IN2(P2_lt_688_n80), 
        .QN(P2_lt_688_n76) );
  NAND2X0 P2_lt_688_U61 ( .IN1(P2_N5022), .IN2(P2_lt_688_n78), 
        .QN(P2_lt_688_n77) );
  NAND2X0 P2_lt_688_U60 ( .IN1(P2_lt_688_n76), .IN2(P2_lt_688_n77), 
        .QN(P2_lt_688_n75) );
  NOR2X0 P2_lt_688_U59 ( .QN(P2_lt_688_n71), .IN1(P2_lt_688_n74), 
        .IN2(P2_lt_688_n75) );
  NOR2X0 P2_lt_688_U58 ( .QN(P2_lt_688_n72), .IN1(P2_N5023), 
        .IN2(P2_lt_688_n73) );
  NOR2X0 P2_lt_688_U57 ( .QN(P2_lt_688_n69), .IN1(P2_lt_688_n71), 
        .IN2(P2_lt_688_n72) );
  INVX0 P2_lt_688_U56 ( .ZN(P2_lt_688_n68), .INP(P2_N5339) );
  OR2X1 P2_lt_688_U55 ( .IN2(P2_N5024), .IN1(P2_lt_688_n68), .Q(P2_lt_688_n70)
         );
  NAND2X0 P2_lt_688_U54 ( .IN1(P2_lt_688_n69), .IN2(P2_lt_688_n70), 
        .QN(P2_lt_688_n66) );
  NAND2X0 P2_lt_688_U53 ( .IN1(P2_N5024), .IN2(P2_lt_688_n68), 
        .QN(P2_lt_688_n67) );
  NAND2X0 P2_lt_688_U52 ( .IN1(P2_lt_688_n66), .IN2(P2_lt_688_n67), 
        .QN(P2_lt_688_n65) );
  NOR2X0 P2_lt_688_U51 ( .QN(P2_lt_688_n61), .IN1(P2_lt_688_n64), 
        .IN2(P2_lt_688_n65) );
  INVX0 P2_lt_688_U157 ( .ZN(P2_lt_688_n5), .INP(P2_N5352) );
  OR2X1 P2_lt_688_U156 ( .IN2(P2_N5037), .IN1(P2_lt_688_n5), .Q(P2_lt_688_n1)
         );
  INVX0 P2_lt_688_U155 ( .ZN(P2_lt_688_n13), .INP(P2_N5350) );
  AND2X1 P2_lt_688_U154 ( .IN1(P2_lt_688_n13), .IN2(P2_N5035), 
        .Q(P2_lt_688_n14) );
  INVX0 P2_lt_688_U153 ( .ZN(P2_lt_688_n23), .INP(P2_N5348) );
  AND2X1 P2_lt_688_U152 ( .IN1(P2_lt_688_n23), .IN2(P2_N5033), 
        .Q(P2_lt_688_n24) );
  INVX0 P2_lt_688_U151 ( .ZN(P2_lt_688_n33), .INP(P2_N5346) );
  AND2X1 P2_lt_688_U150 ( .IN1(P2_lt_688_n33), .IN2(P2_N5031), 
        .Q(P2_lt_688_n34) );
  INVX0 P2_lt_688_U149 ( .ZN(P2_lt_688_n43), .INP(P2_N5344) );
  AND2X1 P2_lt_688_U148 ( .IN1(P2_lt_688_n43), .IN2(P2_N5029), 
        .Q(P2_lt_688_n44) );
  INVX0 P2_lt_688_U147 ( .ZN(P2_lt_688_n53), .INP(P2_N5342) );
  AND2X1 P2_lt_688_U146 ( .IN1(P2_lt_688_n53), .IN2(P2_N5027), 
        .Q(P2_lt_688_n54) );
  INVX0 P2_lt_688_U145 ( .ZN(P2_lt_688_n63), .INP(P2_N5340) );
  AND2X1 P2_lt_688_U144 ( .IN1(P2_lt_688_n63), .IN2(P2_N5025), 
        .Q(P2_lt_688_n64) );
  OR2X1 P1_sub_488_U87 ( .IN2(P1_N5173), .IN1(P1_sub_488_n96), 
        .Q(P1_sub_488_n94) );
  NAND2X0 P1_sub_488_U86 ( .IN1(P1_sub_488_n94), .IN2(P1_sub_488_n95), 
        .QN(P1_sub_488_n93) );
  NAND2X0 P1_sub_488_U85 ( .IN1(P1_sub_488_n92), .IN2(P1_sub_488_n93), 
        .QN(P1_sub_488_n86) );
  NAND2X0 P1_sub_488_U84 ( .IN1(P1_sub_488_n91), .IN2(P1_sub_488_n86), 
        .QN(P1_sub_488_n89) );
  OR2X1 P1_sub_488_U83 ( .IN2(P1_sub_488_n86), .IN1(P1_sub_488_n91), 
        .Q(P1_sub_488_n90) );
  NAND2X0 P1_sub_488_U82 ( .IN1(P1_sub_488_n89), .IN2(P1_sub_488_n90), 
        .QN(P1_N4490) );
  INVX0 P1_sub_488_U81 ( .ZN(P1_sub_488_n75), .INP(P1_N4249) );
  NAND2X0 P1_sub_488_U80 ( .IN1(P1_N5175), .IN2(P1_sub_488_n75), 
        .QN(P1_sub_488_n87) );
  OR2X1 P1_sub_488_U79 ( .IN2(P1_N5175), .IN1(P1_sub_488_n75), 
        .Q(P1_sub_488_n88) );
  NAND2X0 P1_sub_488_U78 ( .IN1(P1_sub_488_n87), .IN2(P1_sub_488_n88), 
        .QN(P1_sub_488_n81) );
  NAND2X0 P1_sub_488_U77 ( .IN1(n7129), .IN2(P1_sub_488_n86), 
        .QN(P1_sub_488_n82) );
  OR2X1 P1_sub_488_U76 ( .IN2(n7129), .IN1(P1_sub_488_n86), .Q(P1_sub_488_n84)
         );
  NAND2X0 P1_sub_488_U75 ( .IN1(P1_sub_488_n84), .IN2(P1_sub_488_n85), 
        .QN(P1_sub_488_n83) );
  NAND2X0 P1_sub_488_U74 ( .IN1(P1_sub_488_n82), .IN2(P1_sub_488_n83), 
        .QN(P1_sub_488_n76) );
  NAND2X0 P1_sub_488_U73 ( .IN1(P1_sub_488_n81), .IN2(P1_sub_488_n76), 
        .QN(P1_sub_488_n79) );
  OR2X1 P1_sub_488_U72 ( .IN2(P1_sub_488_n76), .IN1(P1_sub_488_n81), 
        .Q(P1_sub_488_n80) );
  NAND2X0 P1_sub_488_U71 ( .IN1(P1_sub_488_n79), .IN2(P1_sub_488_n80), 
        .QN(P1_N4491) );
  INVX0 P1_sub_488_U70 ( .ZN(P1_sub_488_n64), .INP(P1_N4250) );
  NAND2X0 P1_sub_488_U69 ( .IN1(P1_N5176), .IN2(P1_sub_488_n64), 
        .QN(P1_sub_488_n77) );
  OR2X1 P1_sub_488_U68 ( .IN2(P1_N5176), .IN1(P1_sub_488_n64), 
        .Q(P1_sub_488_n78) );
  NAND2X0 P1_sub_488_U67 ( .IN1(P1_sub_488_n77), .IN2(P1_sub_488_n78), 
        .QN(P1_sub_488_n71) );
  NAND2X0 P1_sub_488_U66 ( .IN1(P1_N5175), .IN2(P1_sub_488_n76), 
        .QN(P1_sub_488_n72) );
  OR2X1 P1_sub_488_U65 ( .IN2(P1_N5175), .IN1(P1_sub_488_n76), 
        .Q(P1_sub_488_n74) );
  NAND2X0 P1_sub_488_U64 ( .IN1(P1_sub_488_n74), .IN2(P1_sub_488_n75), 
        .QN(P1_sub_488_n73) );
  NAND2X0 P1_sub_488_U63 ( .IN1(P1_sub_488_n72), .IN2(P1_sub_488_n73), 
        .QN(P1_sub_488_n65) );
  NAND2X0 P1_sub_488_U62 ( .IN1(P1_sub_488_n71), .IN2(P1_sub_488_n65), 
        .QN(P1_sub_488_n69) );
  OR2X1 P1_sub_488_U61 ( .IN2(P1_sub_488_n65), .IN1(P1_sub_488_n71), 
        .Q(P1_sub_488_n70) );
  NAND2X0 P1_sub_488_U60 ( .IN1(P1_sub_488_n69), .IN2(P1_sub_488_n70), 
        .QN(P1_N4492) );
  OR2X1 P1_sub_488_U58 ( .IN2(P1_N4251), .IN1(n7117), .Q(P1_sub_488_n66) );
  NAND2X0 P1_sub_488_U57 ( .IN1(P1_N4251), .IN2(n7117), .QN(P1_sub_488_n67) );
  NAND2X0 P1_sub_488_U56 ( .IN1(P1_sub_488_n66), .IN2(P1_sub_488_n67), 
        .QN(P1_sub_488_n60) );
  NAND2X0 P1_sub_488_U55 ( .IN1(P1_N5176), .IN2(P1_sub_488_n65), 
        .QN(P1_sub_488_n61) );
  OR2X1 P1_sub_488_U54 ( .IN2(P1_N5176), .IN1(P1_sub_488_n65), 
        .Q(P1_sub_488_n63) );
  NAND2X0 P1_sub_488_U53 ( .IN1(P1_sub_488_n63), .IN2(P1_sub_488_n64), 
        .QN(P1_sub_488_n62) );
  NAND2X0 P1_sub_488_U52 ( .IN1(P1_sub_488_n61), .IN2(P1_sub_488_n62), 
        .QN(P1_sub_488_n59) );
  NAND2X0 P1_sub_488_U51 ( .IN1(P1_sub_488_n60), .IN2(P1_sub_488_n59), 
        .QN(P1_sub_488_n57) );
  OR2X1 P1_sub_488_U50 ( .IN2(P1_sub_488_n60), .IN1(P1_sub_488_n59), 
        .Q(P1_sub_488_n58) );
  NAND2X0 P1_sub_488_U49 ( .IN1(P1_sub_488_n57), .IN2(P1_sub_488_n58), 
        .QN(P1_N4493) );
  NAND2X0 P1_sub_488_U48 ( .IN1(n7046), .IN2(P1_sub_488_n56), 
        .QN(P1_sub_488_n54) );
  OR2X1 P1_sub_488_U47 ( .IN2(n7046), .IN1(P1_sub_488_n56), .Q(P1_sub_488_n55)
         );
  NAND2X0 P1_sub_488_U46 ( .IN1(P1_sub_488_n54), .IN2(P1_sub_488_n55), 
        .QN(P1_sub_488_n52) );
  NAND2X0 P1_sub_488_U45 ( .IN1(P1_sub_488_n52), .IN2(P1_sub_488_n53), 
        .QN(P1_sub_488_n50) );
  OR2X1 P1_sub_488_U44 ( .IN2(P1_sub_488_n53), .IN1(P1_sub_488_n52), 
        .Q(P1_sub_488_n51) );
  NAND2X0 P1_sub_488_U43 ( .IN1(P1_sub_488_n50), .IN2(P1_sub_488_n51), 
        .QN(P1_N4467) );
  NAND2X0 P1_sub_488_U42 ( .IN1(n7041), .IN2(P1_sub_488_n49), 
        .QN(P1_sub_488_n47) );
  OR2X1 P1_sub_488_U41 ( .IN2(n7041), .IN1(P1_sub_488_n49), .Q(P1_sub_488_n48)
         );
  NAND2X0 P1_sub_488_U40 ( .IN1(P1_sub_488_n47), .IN2(P1_sub_488_n48), 
        .QN(P1_sub_488_n45) );
  NAND2X0 P1_sub_488_U39 ( .IN1(P1_sub_488_n45), .IN2(P1_sub_488_n46), 
        .QN(P1_sub_488_n43) );
  OR2X1 P1_sub_488_U38 ( .IN2(P1_sub_488_n46), .IN1(P1_sub_488_n45), 
        .Q(P1_sub_488_n44) );
  NAND2X0 P1_sub_488_U37 ( .IN1(P1_sub_488_n43), .IN2(P1_sub_488_n44), 
        .QN(P1_N4468) );
  NAND2X0 P1_sub_488_U36 ( .IN1(n7036), .IN2(P1_sub_488_n42), 
        .QN(P1_sub_488_n40) );
  OR2X1 P1_sub_488_U35 ( .IN2(n7036), .IN1(P1_sub_488_n42), .Q(P1_sub_488_n41)
         );
  NAND2X0 P1_sub_488_U34 ( .IN1(P1_sub_488_n40), .IN2(P1_sub_488_n41), 
        .QN(P1_sub_488_n38) );
  NAND2X0 P1_sub_488_U33 ( .IN1(P1_sub_488_n38), .IN2(P1_sub_488_n39), 
        .QN(P1_sub_488_n36) );
  OR2X1 P1_sub_488_U32 ( .IN2(P1_sub_488_n39), .IN1(P1_sub_488_n38), 
        .Q(P1_sub_488_n37) );
  NAND2X0 P1_sub_488_U31 ( .IN1(P1_sub_488_n36), .IN2(P1_sub_488_n37), 
        .QN(P1_N4469) );
  NAND2X0 P1_sub_488_U30 ( .IN1(n7081), .IN2(P1_sub_488_n35), 
        .QN(P1_sub_488_n33) );
  OR2X1 P1_sub_488_U29 ( .IN2(n7081), .IN1(P1_sub_488_n35), .Q(P1_sub_488_n34)
         );
  NAND2X0 P1_sub_488_U28 ( .IN1(P1_sub_488_n33), .IN2(P1_sub_488_n34), 
        .QN(P1_sub_488_n31) );
  NAND2X0 P1_sub_488_U27 ( .IN1(P1_sub_488_n31), .IN2(P1_sub_488_n32), 
        .QN(P1_sub_488_n29) );
  OR2X1 P1_sub_488_U26 ( .IN2(P1_sub_488_n32), .IN1(P1_sub_488_n31), 
        .Q(P1_sub_488_n30) );
  NAND2X0 P1_sub_488_U25 ( .IN1(P1_sub_488_n29), .IN2(P1_sub_488_n30), 
        .QN(P1_N4470) );
  NAND2X0 P1_sub_488_U24 ( .IN1(n7080), .IN2(P1_sub_488_n28), 
        .QN(P1_sub_488_n26) );
  OR2X1 P1_sub_488_U23 ( .IN2(n7080), .IN1(P1_sub_488_n28), .Q(P1_sub_488_n27)
         );
  NAND2X0 P1_sub_488_U22 ( .IN1(P1_sub_488_n26), .IN2(P1_sub_488_n27), 
        .QN(P1_sub_488_n24) );
  NAND2X0 P1_sub_488_U21 ( .IN1(P1_sub_488_n24), .IN2(P1_sub_488_n25), 
        .QN(P1_sub_488_n22) );
  OR2X1 P1_sub_488_U20 ( .IN2(P1_sub_488_n25), .IN1(P1_sub_488_n24), 
        .Q(P1_sub_488_n23) );
  NAND2X0 P1_sub_488_U19 ( .IN1(P1_sub_488_n22), .IN2(P1_sub_488_n23), 
        .QN(P1_N4471) );
  NAND2X0 P1_sub_488_U18 ( .IN1(P1_N5156), .IN2(P1_sub_488_n21), 
        .QN(P1_sub_488_n19) );
  OR2X1 P1_sub_488_U17 ( .IN2(P1_N5156), .IN1(P1_sub_488_n21), 
        .Q(P1_sub_488_n20) );
  NAND2X0 P1_sub_488_U16 ( .IN1(P1_sub_488_n19), .IN2(P1_sub_488_n20), 
        .QN(P1_sub_488_n17) );
  NAND2X0 P1_sub_488_U15 ( .IN1(P1_sub_488_n17), .IN2(P1_sub_488_n18), 
        .QN(P1_sub_488_n15) );
  OR2X1 P1_sub_488_U14 ( .IN2(P1_sub_488_n18), .IN1(P1_sub_488_n17), 
        .Q(P1_sub_488_n16) );
  NAND2X0 P1_sub_488_U13 ( .IN1(P1_sub_488_n15), .IN2(P1_sub_488_n16), 
        .QN(P1_N4472) );
  NAND2X0 P1_sub_488_U12 ( .IN1(P1_N5157), .IN2(P1_sub_488_n14), 
        .QN(P1_sub_488_n12) );
  OR2X1 P1_sub_488_U11 ( .IN2(P1_N5157), .IN1(P1_sub_488_n14), 
        .Q(P1_sub_488_n13) );
  NAND2X0 P1_sub_488_U10 ( .IN1(P1_sub_488_n12), .IN2(P1_sub_488_n13), 
        .QN(P1_sub_488_n10) );
  NAND2X0 P1_sub_488_U9 ( .IN1(P1_sub_488_n10), .IN2(P1_sub_488_n11), 
        .QN(P1_sub_488_n8) );
  OR2X1 P1_sub_488_U8 ( .IN2(P1_sub_488_n11), .IN1(P1_sub_488_n10), 
        .Q(P1_sub_488_n9) );
  NAND2X0 P1_sub_488_U7 ( .IN1(P1_sub_488_n8), .IN2(P1_sub_488_n9), 
        .QN(P1_N4473) );
  NAND2X0 P1_sub_488_U6 ( .IN1(n7070), .IN2(P1_sub_488_n7), .QN(P1_sub_488_n5)
         );
  OR2X1 P1_sub_488_U5 ( .IN2(n7070), .IN1(P1_sub_488_n7), .Q(P1_sub_488_n6) );
  NAND2X0 P1_sub_488_U4 ( .IN1(P1_sub_488_n5), .IN2(P1_sub_488_n6), 
        .QN(P1_sub_488_n3) );
  NAND2X0 P1_sub_488_U3 ( .IN1(P1_sub_488_n3), .IN2(P1_sub_488_n4), 
        .QN(P1_sub_488_n1) );
  OR2X1 P1_sub_488_U2 ( .IN2(P1_sub_488_n4), .IN1(P1_sub_488_n3), 
        .Q(P1_sub_488_n2) );
  NAND2X0 P1_sub_488_U1 ( .IN1(P1_sub_488_n1), .IN2(P1_sub_488_n2), 
        .QN(P1_N4474) );
  NAND2X0 P1_sub_488_U180 ( .IN1(P1_sub_488_n182), .IN2(P1_sub_488_n183), 
        .QN(P1_sub_488_n181) );
  NAND2X0 P1_sub_488_U179 ( .IN1(P1_sub_488_n180), .IN2(P1_sub_488_n181), 
        .QN(P1_sub_488_n174) );
  NAND2X0 P1_sub_488_U178 ( .IN1(P1_sub_488_n179), .IN2(P1_sub_488_n174), 
        .QN(P1_sub_488_n177) );
  OR2X1 P1_sub_488_U177 ( .IN2(P1_sub_488_n174), .IN1(P1_sub_488_n179), 
        .Q(P1_sub_488_n178) );
  NAND2X0 P1_sub_488_U176 ( .IN1(P1_sub_488_n177), .IN2(P1_sub_488_n178), 
        .QN(P1_N4482) );
  INVX0 P1_sub_488_U175 ( .ZN(P1_sub_488_n163), .INP(P1_N4241) );
  NAND2X0 P1_sub_488_U174 ( .IN1(n7103), .IN2(P1_sub_488_n163), 
        .QN(P1_sub_488_n175) );
  OR2X1 P1_sub_488_U173 ( .IN2(n7103), .IN1(P1_sub_488_n163), 
        .Q(P1_sub_488_n176) );
  NAND2X0 P1_sub_488_U172 ( .IN1(P1_sub_488_n175), .IN2(P1_sub_488_n176), 
        .QN(P1_sub_488_n169) );
  NAND2X0 P1_sub_488_U171 ( .IN1(P1_N5166), .IN2(P1_sub_488_n174), 
        .QN(P1_sub_488_n170) );
  OR2X1 P1_sub_488_U170 ( .IN2(P1_N5166), .IN1(P1_sub_488_n174), 
        .Q(P1_sub_488_n172) );
  NAND2X0 P1_sub_488_U169 ( .IN1(P1_sub_488_n172), .IN2(P1_sub_488_n173), 
        .QN(P1_sub_488_n171) );
  NAND2X0 P1_sub_488_U168 ( .IN1(P1_sub_488_n170), .IN2(P1_sub_488_n171), 
        .QN(P1_sub_488_n164) );
  NAND2X0 P1_sub_488_U167 ( .IN1(P1_sub_488_n169), .IN2(P1_sub_488_n164), 
        .QN(P1_sub_488_n167) );
  OR2X1 P1_sub_488_U166 ( .IN2(P1_sub_488_n164), .IN1(P1_sub_488_n169), 
        .Q(P1_sub_488_n168) );
  NAND2X0 P1_sub_488_U165 ( .IN1(P1_sub_488_n167), .IN2(P1_sub_488_n168), 
        .QN(P1_N4483) );
  INVX0 P1_sub_488_U164 ( .ZN(P1_sub_488_n145), .INP(P1_N4242) );
  NAND2X0 P1_sub_488_U163 ( .IN1(P1_N5168), .IN2(P1_sub_488_n145), 
        .QN(P1_sub_488_n165) );
  OR2X1 P1_sub_488_U162 ( .IN2(P1_N5168), .IN1(P1_sub_488_n145), 
        .Q(P1_sub_488_n166) );
  NAND2X0 P1_sub_488_U161 ( .IN1(P1_sub_488_n165), .IN2(P1_sub_488_n166), 
        .QN(P1_sub_488_n159) );
  NAND2X0 P1_sub_488_U160 ( .IN1(n7103), .IN2(P1_sub_488_n164), 
        .QN(P1_sub_488_n160) );
  OR2X1 P1_sub_488_U159 ( .IN2(n7103), .IN1(P1_sub_488_n164), 
        .Q(P1_sub_488_n162) );
  NAND2X0 P1_sub_488_U158 ( .IN1(P1_sub_488_n162), .IN2(P1_sub_488_n163), 
        .QN(P1_sub_488_n161) );
  NAND2X0 P1_sub_488_U157 ( .IN1(P1_sub_488_n160), .IN2(P1_sub_488_n161), 
        .QN(P1_sub_488_n146) );
  NAND2X0 P1_sub_488_U156 ( .IN1(P1_sub_488_n159), .IN2(P1_sub_488_n146), 
        .QN(P1_sub_488_n157) );
  OR2X1 P1_sub_488_U155 ( .IN2(P1_sub_488_n146), .IN1(P1_sub_488_n159), 
        .Q(P1_sub_488_n158) );
  NAND2X0 P1_sub_488_U154 ( .IN1(P1_sub_488_n157), .IN2(P1_sub_488_n158), 
        .QN(P1_N4484) );
  NAND2X0 P1_sub_488_U153 ( .IN1(P1_N5150), .IN2(P1_sub_488_n156), 
        .QN(P1_sub_488_n153) );
  NAND2X0 P1_sub_488_U152 ( .IN1(P1_N4224), .IN2(n7048), .QN(P1_sub_488_n154)
         );
  NAND2X0 P1_sub_488_U151 ( .IN1(P1_sub_488_n153), .IN2(P1_sub_488_n154), 
        .QN(P1_sub_488_n151) );
  NAND2X0 P1_sub_488_U150 ( .IN1(P1_sub_488_n151), .IN2(P1_sub_488_n152), 
        .QN(P1_sub_488_n149) );
  OR2X1 P1_sub_488_U149 ( .IN2(P1_sub_488_n152), .IN1(P1_sub_488_n151), 
        .Q(P1_sub_488_n150) );
  NAND2X0 P1_sub_488_U148 ( .IN1(P1_sub_488_n149), .IN2(P1_sub_488_n150), 
        .QN(P1_N4466) );
  INVX0 P1_sub_488_U147 ( .ZN(P1_sub_488_n135), .INP(P1_N4243) );
  NAND2X0 P1_sub_488_U146 ( .IN1(n7096), .IN2(P1_sub_488_n135), 
        .QN(P1_sub_488_n147) );
  OR2X1 P1_sub_488_U145 ( .IN2(n7096), .IN1(P1_sub_488_n135), 
        .Q(P1_sub_488_n148) );
  NAND2X0 P1_sub_488_U144 ( .IN1(P1_sub_488_n147), .IN2(P1_sub_488_n148), 
        .QN(P1_sub_488_n141) );
  NAND2X0 P1_sub_488_U143 ( .IN1(P1_N5168), .IN2(P1_sub_488_n146), 
        .QN(P1_sub_488_n142) );
  OR2X1 P1_sub_488_U142 ( .IN2(P1_N5168), .IN1(P1_sub_488_n146), 
        .Q(P1_sub_488_n144) );
  NAND2X0 P1_sub_488_U141 ( .IN1(P1_sub_488_n144), .IN2(P1_sub_488_n145), 
        .QN(P1_sub_488_n143) );
  NAND2X0 P1_sub_488_U140 ( .IN1(P1_sub_488_n142), .IN2(P1_sub_488_n143), 
        .QN(P1_sub_488_n136) );
  NAND2X0 P1_sub_488_U139 ( .IN1(P1_sub_488_n141), .IN2(P1_sub_488_n136), 
        .QN(P1_sub_488_n139) );
  OR2X1 P1_sub_488_U138 ( .IN2(P1_sub_488_n136), .IN1(P1_sub_488_n141), 
        .Q(P1_sub_488_n140) );
  NAND2X0 P1_sub_488_U137 ( .IN1(P1_sub_488_n139), .IN2(P1_sub_488_n140), 
        .QN(P1_N4485) );
  INVX0 P1_sub_488_U136 ( .ZN(P1_sub_488_n125), .INP(P1_N4244) );
  NAND2X0 P1_sub_488_U135 ( .IN1(n7093), .IN2(P1_sub_488_n125), 
        .QN(P1_sub_488_n137) );
  OR2X1 P1_sub_488_U134 ( .IN2(n7093), .IN1(P1_sub_488_n125), 
        .Q(P1_sub_488_n138) );
  NAND2X0 P1_sub_488_U133 ( .IN1(P1_sub_488_n137), .IN2(P1_sub_488_n138), 
        .QN(P1_sub_488_n131) );
  NAND2X0 P1_sub_488_U132 ( .IN1(n7096), .IN2(P1_sub_488_n136), 
        .QN(P1_sub_488_n132) );
  OR2X1 P1_sub_488_U131 ( .IN2(n7096), .IN1(P1_sub_488_n136), 
        .Q(P1_sub_488_n134) );
  NAND2X0 P1_sub_488_U130 ( .IN1(P1_sub_488_n134), .IN2(P1_sub_488_n135), 
        .QN(P1_sub_488_n133) );
  NAND2X0 P1_sub_488_U129 ( .IN1(P1_sub_488_n132), .IN2(P1_sub_488_n133), 
        .QN(P1_sub_488_n126) );
  NAND2X0 P1_sub_488_U128 ( .IN1(P1_sub_488_n131), .IN2(P1_sub_488_n126), 
        .QN(P1_sub_488_n129) );
  OR2X1 P1_sub_488_U127 ( .IN2(P1_sub_488_n126), .IN1(P1_sub_488_n131), 
        .Q(P1_sub_488_n130) );
  NAND2X0 P1_sub_488_U126 ( .IN1(P1_sub_488_n129), .IN2(P1_sub_488_n130), 
        .QN(P1_N4486) );
  INVX0 P1_sub_488_U125 ( .ZN(P1_sub_488_n115), .INP(P1_N4245) );
  NAND2X0 P1_sub_488_U124 ( .IN1(n7089), .IN2(P1_sub_488_n115), 
        .QN(P1_sub_488_n127) );
  OR2X1 P1_sub_488_U123 ( .IN2(n7089), .IN1(P1_sub_488_n115), 
        .Q(P1_sub_488_n128) );
  NAND2X0 P1_sub_488_U122 ( .IN1(P1_sub_488_n127), .IN2(P1_sub_488_n128), 
        .QN(P1_sub_488_n121) );
  NAND2X0 P1_sub_488_U121 ( .IN1(n7093), .IN2(P1_sub_488_n126), 
        .QN(P1_sub_488_n122) );
  OR2X1 P1_sub_488_U120 ( .IN2(n7093), .IN1(P1_sub_488_n126), 
        .Q(P1_sub_488_n124) );
  NAND2X0 P1_sub_488_U119 ( .IN1(P1_sub_488_n124), .IN2(P1_sub_488_n125), 
        .QN(P1_sub_488_n123) );
  NAND2X0 P1_sub_488_U118 ( .IN1(P1_sub_488_n122), .IN2(P1_sub_488_n123), 
        .QN(P1_sub_488_n116) );
  NAND2X0 P1_sub_488_U117 ( .IN1(P1_sub_488_n121), .IN2(P1_sub_488_n116), 
        .QN(P1_sub_488_n119) );
  OR2X1 P1_sub_488_U116 ( .IN2(P1_sub_488_n116), .IN1(P1_sub_488_n121), 
        .Q(P1_sub_488_n120) );
  NAND2X0 P1_sub_488_U115 ( .IN1(P1_sub_488_n119), .IN2(P1_sub_488_n120), 
        .QN(P1_N4487) );
  INVX0 P1_sub_488_U114 ( .ZN(P1_sub_488_n105), .INP(P1_N4246) );
  NAND2X0 P1_sub_488_U113 ( .IN1(P1_N5172), .IN2(P1_sub_488_n105), 
        .QN(P1_sub_488_n117) );
  OR2X1 P1_sub_488_U112 ( .IN2(P1_N5172), .IN1(P1_sub_488_n105), 
        .Q(P1_sub_488_n118) );
  NAND2X0 P1_sub_488_U111 ( .IN1(P1_sub_488_n117), .IN2(P1_sub_488_n118), 
        .QN(P1_sub_488_n111) );
  NAND2X0 P1_sub_488_U110 ( .IN1(n7089), .IN2(P1_sub_488_n116), 
        .QN(P1_sub_488_n112) );
  OR2X1 P1_sub_488_U109 ( .IN2(n7089), .IN1(P1_sub_488_n116), 
        .Q(P1_sub_488_n114) );
  NAND2X0 P1_sub_488_U108 ( .IN1(P1_sub_488_n114), .IN2(P1_sub_488_n115), 
        .QN(P1_sub_488_n113) );
  NAND2X0 P1_sub_488_U107 ( .IN1(P1_sub_488_n112), .IN2(P1_sub_488_n113), 
        .QN(P1_sub_488_n106) );
  NAND2X0 P1_sub_488_U106 ( .IN1(P1_sub_488_n111), .IN2(P1_sub_488_n106), 
        .QN(P1_sub_488_n109) );
  OR2X1 P1_sub_488_U105 ( .IN2(P1_sub_488_n106), .IN1(P1_sub_488_n111), 
        .Q(P1_sub_488_n110) );
  NAND2X0 P1_sub_488_U104 ( .IN1(P1_sub_488_n109), .IN2(P1_sub_488_n110), 
        .QN(P1_N4488) );
  INVX0 P1_sub_488_U103 ( .ZN(P1_sub_488_n95), .INP(P1_N4247) );
  NAND2X0 P1_sub_488_U102 ( .IN1(P1_N5173), .IN2(P1_sub_488_n95), 
        .QN(P1_sub_488_n107) );
  OR2X1 P1_sub_488_U101 ( .IN2(P1_N5173), .IN1(P1_sub_488_n95), 
        .Q(P1_sub_488_n108) );
  NAND2X0 P1_sub_488_U100 ( .IN1(P1_sub_488_n107), .IN2(P1_sub_488_n108), 
        .QN(P1_sub_488_n101) );
  NAND2X0 P1_sub_488_U99 ( .IN1(P1_N5172), .IN2(P1_sub_488_n106), 
        .QN(P1_sub_488_n102) );
  OR2X1 P1_sub_488_U98 ( .IN2(P1_N5172), .IN1(P1_sub_488_n106), 
        .Q(P1_sub_488_n104) );
  NAND2X0 P1_sub_488_U97 ( .IN1(P1_sub_488_n104), .IN2(P1_sub_488_n105), 
        .QN(P1_sub_488_n103) );
  NAND2X0 P1_sub_488_U96 ( .IN1(P1_sub_488_n102), .IN2(P1_sub_488_n103), 
        .QN(P1_sub_488_n96) );
  NAND2X0 P1_sub_488_U95 ( .IN1(P1_sub_488_n101), .IN2(P1_sub_488_n96), 
        .QN(P1_sub_488_n99) );
  OR2X1 P1_sub_488_U94 ( .IN2(P1_sub_488_n96), .IN1(P1_sub_488_n101), 
        .Q(P1_sub_488_n100) );
  NAND2X0 P1_sub_488_U93 ( .IN1(P1_sub_488_n99), .IN2(P1_sub_488_n100), 
        .QN(P1_N4489) );
  INVX0 P1_sub_488_U92 ( .ZN(P1_sub_488_n85), .INP(P1_N4248) );
  NAND2X0 P1_sub_488_U91 ( .IN1(n7129), .IN2(P1_sub_488_n85), 
        .QN(P1_sub_488_n97) );
  OR2X1 P1_sub_488_U90 ( .IN2(n7129), .IN1(P1_sub_488_n85), .Q(P1_sub_488_n98)
         );
  NAND2X0 P1_sub_488_U89 ( .IN1(P1_sub_488_n97), .IN2(P1_sub_488_n98), 
        .QN(P1_sub_488_n91) );
  NAND2X0 P1_sub_488_U88 ( .IN1(P1_N5173), .IN2(P1_sub_488_n96), 
        .QN(P1_sub_488_n92) );
  INVX0 P1_sub_488_U273 ( .ZN(P1_sub_488_n28), .INP(P1_N4229) );
  NAND2X0 P1_sub_488_U272 ( .IN1(P1_sub_488_n261), .IN2(P1_sub_488_n28), 
        .QN(P1_sub_488_n260) );
  NAND2X0 P1_sub_488_U271 ( .IN1(P1_sub_488_n259), .IN2(P1_sub_488_n260), 
        .QN(P1_sub_488_n18) );
  NAND2X0 P1_sub_488_U270 ( .IN1(P1_N5156), .IN2(P1_sub_488_n18), 
        .QN(P1_sub_488_n256) );
  OR2X1 P1_sub_488_U269 ( .IN2(P1_N5156), .IN1(P1_sub_488_n18), 
        .Q(P1_sub_488_n258) );
  INVX0 P1_sub_488_U268 ( .ZN(P1_sub_488_n21), .INP(P1_N4230) );
  NAND2X0 P1_sub_488_U267 ( .IN1(P1_sub_488_n258), .IN2(P1_sub_488_n21), 
        .QN(P1_sub_488_n257) );
  NAND2X0 P1_sub_488_U266 ( .IN1(P1_sub_488_n256), .IN2(P1_sub_488_n257), 
        .QN(P1_sub_488_n11) );
  NAND2X0 P1_sub_488_U265 ( .IN1(P1_N5157), .IN2(P1_sub_488_n11), 
        .QN(P1_sub_488_n253) );
  OR2X1 P1_sub_488_U264 ( .IN2(P1_N5157), .IN1(P1_sub_488_n11), 
        .Q(P1_sub_488_n255) );
  INVX0 P1_sub_488_U263 ( .ZN(P1_sub_488_n14), .INP(P1_N4231) );
  NAND2X0 P1_sub_488_U262 ( .IN1(P1_sub_488_n255), .IN2(P1_sub_488_n14), 
        .QN(P1_sub_488_n254) );
  NAND2X0 P1_sub_488_U261 ( .IN1(P1_sub_488_n253), .IN2(P1_sub_488_n254), 
        .QN(P1_sub_488_n4) );
  NAND2X0 P1_sub_488_U260 ( .IN1(n7070), .IN2(P1_sub_488_n4), 
        .QN(P1_sub_488_n250) );
  OR2X1 P1_sub_488_U259 ( .IN2(n7070), .IN1(P1_sub_488_n4), 
        .Q(P1_sub_488_n252) );
  INVX0 P1_sub_488_U258 ( .ZN(P1_sub_488_n7), .INP(P1_N4232) );
  NAND2X0 P1_sub_488_U257 ( .IN1(P1_sub_488_n252), .IN2(P1_sub_488_n7), 
        .QN(P1_sub_488_n251) );
  NAND2X0 P1_sub_488_U256 ( .IN1(P1_sub_488_n250), .IN2(P1_sub_488_n251), 
        .QN(P1_sub_488_n244) );
  NAND2X0 P1_sub_488_U255 ( .IN1(P1_sub_488_n249), .IN2(P1_sub_488_n244), 
        .QN(P1_sub_488_n247) );
  OR2X1 P1_sub_488_U254 ( .IN2(P1_sub_488_n244), .IN1(P1_sub_488_n249), 
        .Q(P1_sub_488_n248) );
  NAND2X0 P1_sub_488_U253 ( .IN1(P1_sub_488_n247), .IN2(P1_sub_488_n248), 
        .QN(P1_N4475) );
  INVX0 P1_sub_488_U252 ( .ZN(P1_sub_488_n233), .INP(P1_N4234) );
  NAND2X0 P1_sub_488_U251 ( .IN1(n7062), .IN2(P1_sub_488_n233), 
        .QN(P1_sub_488_n245) );
  OR2X1 P1_sub_488_U250 ( .IN2(n7062), .IN1(P1_sub_488_n233), 
        .Q(P1_sub_488_n246) );
  NAND2X0 P1_sub_488_U249 ( .IN1(P1_sub_488_n245), .IN2(P1_sub_488_n246), 
        .QN(P1_sub_488_n239) );
  NAND2X0 P1_sub_488_U248 ( .IN1(n7066), .IN2(P1_sub_488_n244), 
        .QN(P1_sub_488_n240) );
  OR2X1 P1_sub_488_U247 ( .IN2(n7066), .IN1(P1_sub_488_n244), 
        .Q(P1_sub_488_n242) );
  NAND2X0 P1_sub_488_U246 ( .IN1(P1_sub_488_n242), .IN2(P1_sub_488_n243), 
        .QN(P1_sub_488_n241) );
  NAND2X0 P1_sub_488_U245 ( .IN1(P1_sub_488_n240), .IN2(P1_sub_488_n241), 
        .QN(P1_sub_488_n234) );
  NAND2X0 P1_sub_488_U244 ( .IN1(P1_sub_488_n239), .IN2(P1_sub_488_n234), 
        .QN(P1_sub_488_n237) );
  OR2X1 P1_sub_488_U243 ( .IN2(P1_sub_488_n234), .IN1(P1_sub_488_n239), 
        .Q(P1_sub_488_n238) );
  NAND2X0 P1_sub_488_U242 ( .IN1(P1_sub_488_n237), .IN2(P1_sub_488_n238), 
        .QN(P1_N4476) );
  INVX0 P1_sub_488_U241 ( .ZN(P1_sub_488_n223), .INP(P1_N4235) );
  NAND2X0 P1_sub_488_U240 ( .IN1(n7059), .IN2(P1_sub_488_n223), 
        .QN(P1_sub_488_n235) );
  OR2X1 P1_sub_488_U239 ( .IN2(n7059), .IN1(P1_sub_488_n223), 
        .Q(P1_sub_488_n236) );
  NAND2X0 P1_sub_488_U238 ( .IN1(P1_sub_488_n235), .IN2(P1_sub_488_n236), 
        .QN(P1_sub_488_n229) );
  NAND2X0 P1_sub_488_U237 ( .IN1(n7062), .IN2(P1_sub_488_n234), 
        .QN(P1_sub_488_n230) );
  OR2X1 P1_sub_488_U236 ( .IN2(n7062), .IN1(P1_sub_488_n234), 
        .Q(P1_sub_488_n232) );
  NAND2X0 P1_sub_488_U235 ( .IN1(P1_sub_488_n232), .IN2(P1_sub_488_n233), 
        .QN(P1_sub_488_n231) );
  NAND2X0 P1_sub_488_U234 ( .IN1(P1_sub_488_n230), .IN2(P1_sub_488_n231), 
        .QN(P1_sub_488_n224) );
  NAND2X0 P1_sub_488_U233 ( .IN1(P1_sub_488_n229), .IN2(P1_sub_488_n224), 
        .QN(P1_sub_488_n227) );
  OR2X1 P1_sub_488_U232 ( .IN2(P1_sub_488_n224), .IN1(P1_sub_488_n229), 
        .Q(P1_sub_488_n228) );
  NAND2X0 P1_sub_488_U231 ( .IN1(P1_sub_488_n227), .IN2(P1_sub_488_n228), 
        .QN(P1_N4477) );
  INVX0 P1_sub_488_U230 ( .ZN(P1_sub_488_n213), .INP(P1_N4236) );
  NAND2X0 P1_sub_488_U229 ( .IN1(n7055), .IN2(P1_sub_488_n213), 
        .QN(P1_sub_488_n225) );
  OR2X1 P1_sub_488_U228 ( .IN2(n7055), .IN1(P1_sub_488_n213), 
        .Q(P1_sub_488_n226) );
  NAND2X0 P1_sub_488_U227 ( .IN1(P1_sub_488_n225), .IN2(P1_sub_488_n226), 
        .QN(P1_sub_488_n219) );
  NAND2X0 P1_sub_488_U226 ( .IN1(n7059), .IN2(P1_sub_488_n224), 
        .QN(P1_sub_488_n220) );
  OR2X1 P1_sub_488_U225 ( .IN2(n7059), .IN1(P1_sub_488_n224), 
        .Q(P1_sub_488_n222) );
  NAND2X0 P1_sub_488_U224 ( .IN1(P1_sub_488_n222), .IN2(P1_sub_488_n223), 
        .QN(P1_sub_488_n221) );
  NAND2X0 P1_sub_488_U223 ( .IN1(P1_sub_488_n220), .IN2(P1_sub_488_n221), 
        .QN(P1_sub_488_n214) );
  NAND2X0 P1_sub_488_U222 ( .IN1(P1_sub_488_n219), .IN2(P1_sub_488_n214), 
        .QN(P1_sub_488_n217) );
  OR2X1 P1_sub_488_U221 ( .IN2(P1_sub_488_n214), .IN1(P1_sub_488_n219), 
        .Q(P1_sub_488_n218) );
  NAND2X0 P1_sub_488_U220 ( .IN1(P1_sub_488_n217), .IN2(P1_sub_488_n218), 
        .QN(P1_N4478) );
  INVX0 P1_sub_488_U219 ( .ZN(P1_sub_488_n203), .INP(P1_N4237) );
  NAND2X0 P1_sub_488_U218 ( .IN1(n7116), .IN2(P1_sub_488_n203), 
        .QN(P1_sub_488_n215) );
  OR2X1 P1_sub_488_U217 ( .IN2(n7116), .IN1(P1_sub_488_n203), 
        .Q(P1_sub_488_n216) );
  NAND2X0 P1_sub_488_U216 ( .IN1(P1_sub_488_n215), .IN2(P1_sub_488_n216), 
        .QN(P1_sub_488_n209) );
  NAND2X0 P1_sub_488_U215 ( .IN1(n7055), .IN2(P1_sub_488_n214), 
        .QN(P1_sub_488_n210) );
  OR2X1 P1_sub_488_U214 ( .IN2(n7055), .IN1(P1_sub_488_n214), 
        .Q(P1_sub_488_n212) );
  NAND2X0 P1_sub_488_U213 ( .IN1(P1_sub_488_n212), .IN2(P1_sub_488_n213), 
        .QN(P1_sub_488_n211) );
  NAND2X0 P1_sub_488_U212 ( .IN1(P1_sub_488_n210), .IN2(P1_sub_488_n211), 
        .QN(P1_sub_488_n204) );
  NAND2X0 P1_sub_488_U211 ( .IN1(P1_sub_488_n209), .IN2(P1_sub_488_n204), 
        .QN(P1_sub_488_n207) );
  OR2X1 P1_sub_488_U210 ( .IN2(P1_sub_488_n204), .IN1(P1_sub_488_n209), 
        .Q(P1_sub_488_n208) );
  NAND2X0 P1_sub_488_U209 ( .IN1(P1_sub_488_n207), .IN2(P1_sub_488_n208), 
        .QN(P1_N4479) );
  INVX0 P1_sub_488_U208 ( .ZN(P1_sub_488_n193), .INP(P1_N4238) );
  NAND2X0 P1_sub_488_U207 ( .IN1(P1_N5164), .IN2(P1_sub_488_n193), 
        .QN(P1_sub_488_n205) );
  OR2X1 P1_sub_488_U206 ( .IN2(P1_N5164), .IN1(P1_sub_488_n193), 
        .Q(P1_sub_488_n206) );
  NAND2X0 P1_sub_488_U205 ( .IN1(P1_sub_488_n205), .IN2(P1_sub_488_n206), 
        .QN(P1_sub_488_n199) );
  NAND2X0 P1_sub_488_U204 ( .IN1(n7116), .IN2(P1_sub_488_n204), 
        .QN(P1_sub_488_n200) );
  OR2X1 P1_sub_488_U203 ( .IN2(n7116), .IN1(P1_sub_488_n204), 
        .Q(P1_sub_488_n202) );
  NAND2X0 P1_sub_488_U202 ( .IN1(P1_sub_488_n202), .IN2(P1_sub_488_n203), 
        .QN(P1_sub_488_n201) );
  NAND2X0 P1_sub_488_U201 ( .IN1(P1_sub_488_n200), .IN2(P1_sub_488_n201), 
        .QN(P1_sub_488_n194) );
  NAND2X0 P1_sub_488_U200 ( .IN1(P1_sub_488_n199), .IN2(P1_sub_488_n194), 
        .QN(P1_sub_488_n197) );
  OR2X1 P1_sub_488_U199 ( .IN2(P1_sub_488_n194), .IN1(P1_sub_488_n199), 
        .Q(P1_sub_488_n198) );
  NAND2X0 P1_sub_488_U198 ( .IN1(P1_sub_488_n197), .IN2(P1_sub_488_n198), 
        .QN(P1_N4480) );
  INVX0 P1_sub_488_U197 ( .ZN(P1_sub_488_n183), .INP(P1_N4239) );
  NAND2X0 P1_sub_488_U196 ( .IN1(P1_N5165), .IN2(P1_sub_488_n183), 
        .QN(P1_sub_488_n195) );
  OR2X1 P1_sub_488_U195 ( .IN2(P1_N5165), .IN1(P1_sub_488_n183), 
        .Q(P1_sub_488_n196) );
  NAND2X0 P1_sub_488_U194 ( .IN1(P1_sub_488_n195), .IN2(P1_sub_488_n196), 
        .QN(P1_sub_488_n189) );
  NAND2X0 P1_sub_488_U193 ( .IN1(n7113), .IN2(P1_sub_488_n194), 
        .QN(P1_sub_488_n190) );
  OR2X1 P1_sub_488_U192 ( .IN2(n7113), .IN1(P1_sub_488_n194), 
        .Q(P1_sub_488_n192) );
  NAND2X0 P1_sub_488_U191 ( .IN1(P1_sub_488_n192), .IN2(P1_sub_488_n193), 
        .QN(P1_sub_488_n191) );
  NAND2X0 P1_sub_488_U190 ( .IN1(P1_sub_488_n190), .IN2(P1_sub_488_n191), 
        .QN(P1_sub_488_n184) );
  NAND2X0 P1_sub_488_U189 ( .IN1(P1_sub_488_n189), .IN2(P1_sub_488_n184), 
        .QN(P1_sub_488_n187) );
  OR2X1 P1_sub_488_U188 ( .IN2(P1_sub_488_n184), .IN1(P1_sub_488_n189), 
        .Q(P1_sub_488_n188) );
  NAND2X0 P1_sub_488_U187 ( .IN1(P1_sub_488_n187), .IN2(P1_sub_488_n188), 
        .QN(P1_N4481) );
  INVX0 P1_sub_488_U186 ( .ZN(P1_sub_488_n173), .INP(P1_N4240) );
  NAND2X0 P1_sub_488_U185 ( .IN1(P1_N5166), .IN2(P1_sub_488_n173), 
        .QN(P1_sub_488_n185) );
  OR2X1 P1_sub_488_U184 ( .IN2(P1_N5166), .IN1(P1_sub_488_n173), 
        .Q(P1_sub_488_n186) );
  NAND2X0 P1_sub_488_U183 ( .IN1(P1_sub_488_n185), .IN2(P1_sub_488_n186), 
        .QN(P1_sub_488_n179) );
  NAND2X0 P1_sub_488_U182 ( .IN1(n7110), .IN2(P1_sub_488_n184), 
        .QN(P1_sub_488_n180) );
  OR2X1 P1_sub_488_U181 ( .IN2(P1_N5165), .IN1(P1_sub_488_n184), 
        .Q(P1_sub_488_n182) );
  INVX0 P1_sub_488_U310 ( .ZN(P1_sub_488_n281), .INP(P1_N4223) );
  NOR2X0 P1_sub_488_U309 ( .QN(P1_sub_488_n277), .IN1(P1_sub_488_n281), 
        .IN2(n7034) );
  INVX0 P1_sub_488_U308 ( .ZN(P1_sub_488_n152), .INP(P1_sub_488_n277) );
  NAND2X0 P1_sub_488_U307 ( .IN1(n7034), .IN2(P1_sub_488_n281), 
        .QN(P1_sub_488_n280) );
  NAND2X0 P1_sub_488_U306 ( .IN1(P1_sub_488_n152), .IN2(P1_sub_488_n280), 
        .QN(P1_N4465) );
  INVX0 P1_sub_488_U305 ( .ZN(P1_sub_488_n243), .INP(P1_N4233) );
  NAND2X0 P1_sub_488_U304 ( .IN1(n7066), .IN2(P1_sub_488_n243), 
        .QN(P1_sub_488_n278) );
  OR2X1 P1_sub_488_U303 ( .IN2(n7066), .IN1(P1_sub_488_n243), 
        .Q(P1_sub_488_n279) );
  NAND2X0 P1_sub_488_U302 ( .IN1(P1_sub_488_n278), .IN2(P1_sub_488_n279), 
        .QN(P1_sub_488_n249) );
  NAND2X0 P1_sub_488_U301 ( .IN1(P1_N5150), .IN2(P1_sub_488_n152), 
        .QN(P1_sub_488_n274) );
  NAND2X0 P1_sub_488_U299 ( .IN1(P1_sub_488_n277), .IN2(n7048), 
        .QN(P1_sub_488_n276) );
  INVX0 P1_sub_488_U298 ( .ZN(P1_sub_488_n156), .INP(P1_N4224) );
  NAND2X0 P1_sub_488_U297 ( .IN1(P1_sub_488_n276), .IN2(P1_sub_488_n156), 
        .QN(P1_sub_488_n275) );
  NAND2X0 P1_sub_488_U296 ( .IN1(P1_sub_488_n274), .IN2(P1_sub_488_n275), 
        .QN(P1_sub_488_n53) );
  NAND2X0 P1_sub_488_U295 ( .IN1(n7046), .IN2(P1_sub_488_n53), 
        .QN(P1_sub_488_n271) );
  OR2X1 P1_sub_488_U294 ( .IN2(n7046), .IN1(P1_sub_488_n53), 
        .Q(P1_sub_488_n273) );
  INVX0 P1_sub_488_U293 ( .ZN(P1_sub_488_n56), .INP(P1_N4225) );
  NAND2X0 P1_sub_488_U292 ( .IN1(P1_sub_488_n273), .IN2(P1_sub_488_n56), 
        .QN(P1_sub_488_n272) );
  NAND2X0 P1_sub_488_U291 ( .IN1(P1_sub_488_n271), .IN2(P1_sub_488_n272), 
        .QN(P1_sub_488_n46) );
  NAND2X0 P1_sub_488_U290 ( .IN1(n7041), .IN2(P1_sub_488_n46), 
        .QN(P1_sub_488_n268) );
  OR2X1 P1_sub_488_U289 ( .IN2(n7041), .IN1(P1_sub_488_n46), 
        .Q(P1_sub_488_n270) );
  INVX0 P1_sub_488_U288 ( .ZN(P1_sub_488_n49), .INP(P1_N4226) );
  NAND2X0 P1_sub_488_U287 ( .IN1(P1_sub_488_n270), .IN2(P1_sub_488_n49), 
        .QN(P1_sub_488_n269) );
  NAND2X0 P1_sub_488_U286 ( .IN1(P1_sub_488_n268), .IN2(P1_sub_488_n269), 
        .QN(P1_sub_488_n39) );
  NAND2X0 P1_sub_488_U285 ( .IN1(n7036), .IN2(P1_sub_488_n39), 
        .QN(P1_sub_488_n265) );
  OR2X1 P1_sub_488_U284 ( .IN2(n7036), .IN1(P1_sub_488_n39), 
        .Q(P1_sub_488_n267) );
  INVX0 P1_sub_488_U283 ( .ZN(P1_sub_488_n42), .INP(P1_N4227) );
  NAND2X0 P1_sub_488_U282 ( .IN1(P1_sub_488_n267), .IN2(P1_sub_488_n42), 
        .QN(P1_sub_488_n266) );
  NAND2X0 P1_sub_488_U281 ( .IN1(P1_sub_488_n265), .IN2(P1_sub_488_n266), 
        .QN(P1_sub_488_n32) );
  NAND2X0 P1_sub_488_U280 ( .IN1(n7081), .IN2(P1_sub_488_n32), 
        .QN(P1_sub_488_n262) );
  OR2X1 P1_sub_488_U279 ( .IN2(n7081), .IN1(P1_sub_488_n32), 
        .Q(P1_sub_488_n264) );
  INVX0 P1_sub_488_U278 ( .ZN(P1_sub_488_n35), .INP(P1_N4228) );
  NAND2X0 P1_sub_488_U277 ( .IN1(P1_sub_488_n264), .IN2(P1_sub_488_n35), 
        .QN(P1_sub_488_n263) );
  NAND2X0 P1_sub_488_U276 ( .IN1(P1_sub_488_n262), .IN2(P1_sub_488_n263), 
        .QN(P1_sub_488_n25) );
  NAND2X0 P1_sub_488_U275 ( .IN1(n7080), .IN2(P1_sub_488_n25), 
        .QN(P1_sub_488_n259) );
  OR2X1 P1_sub_488_U274 ( .IN2(n7080), .IN1(P1_sub_488_n25), 
        .Q(P1_sub_488_n261) );
  NOR2X0 P1_lt_178_U58 ( .QN(P1_lt_178_n72), .IN1(P1_N5101), 
        .IN2(P1_lt_178_n73) );
  NOR2X0 P1_lt_178_U57 ( .QN(P1_lt_178_n69), .IN1(P1_lt_178_n71), 
        .IN2(P1_lt_178_n72) );
  INVX0 P1_lt_178_U56 ( .ZN(P1_lt_178_n68), .INP(P1_N5417) );
  OR2X1 P1_lt_178_U55 ( .IN2(P1_N5102), .IN1(P1_lt_178_n68), .Q(P1_lt_178_n70)
         );
  NAND2X0 P1_lt_178_U54 ( .IN1(P1_lt_178_n69), .IN2(P1_lt_178_n70), 
        .QN(P1_lt_178_n66) );
  NAND2X0 P1_lt_178_U53 ( .IN1(P1_N5102), .IN2(P1_lt_178_n68), 
        .QN(P1_lt_178_n67) );
  NAND2X0 P1_lt_178_U52 ( .IN1(P1_lt_178_n66), .IN2(P1_lt_178_n67), 
        .QN(P1_lt_178_n65) );
  NOR2X0 P1_lt_178_U51 ( .QN(P1_lt_178_n61), .IN1(P1_lt_178_n64), 
        .IN2(P1_lt_178_n65) );
  NOR2X0 P1_lt_178_U50 ( .QN(P1_lt_178_n62), .IN1(P1_N5103), 
        .IN2(P1_lt_178_n63) );
  NOR2X0 P1_lt_178_U49 ( .QN(P1_lt_178_n59), .IN1(P1_lt_178_n61), 
        .IN2(P1_lt_178_n62) );
  INVX0 P1_lt_178_U48 ( .ZN(P1_lt_178_n58), .INP(P1_N5419) );
  OR2X1 P1_lt_178_U47 ( .IN2(P1_N5104), .IN1(P1_lt_178_n58), .Q(P1_lt_178_n60)
         );
  NAND2X0 P1_lt_178_U46 ( .IN1(P1_lt_178_n59), .IN2(P1_lt_178_n60), 
        .QN(P1_lt_178_n56) );
  NAND2X0 P1_lt_178_U45 ( .IN1(P1_N5104), .IN2(P1_lt_178_n58), 
        .QN(P1_lt_178_n57) );
  NAND2X0 P1_lt_178_U44 ( .IN1(P1_lt_178_n56), .IN2(P1_lt_178_n57), 
        .QN(P1_lt_178_n55) );
  NOR2X0 P1_lt_178_U43 ( .QN(P1_lt_178_n51), .IN1(P1_lt_178_n54), 
        .IN2(P1_lt_178_n55) );
  NOR2X0 P1_lt_178_U42 ( .QN(P1_lt_178_n52), .IN1(P1_N5105), 
        .IN2(P1_lt_178_n53) );
  NOR2X0 P1_lt_178_U41 ( .QN(P1_lt_178_n49), .IN1(P1_lt_178_n51), 
        .IN2(P1_lt_178_n52) );
  INVX0 P1_lt_178_U40 ( .ZN(P1_lt_178_n48), .INP(P1_N5421) );
  OR2X1 P1_lt_178_U39 ( .IN2(P1_N5106), .IN1(P1_lt_178_n48), .Q(P1_lt_178_n50)
         );
  NAND2X0 P1_lt_178_U38 ( .IN1(P1_lt_178_n49), .IN2(P1_lt_178_n50), 
        .QN(P1_lt_178_n46) );
  NAND2X0 P1_lt_178_U37 ( .IN1(P1_N5106), .IN2(P1_lt_178_n48), 
        .QN(P1_lt_178_n47) );
  NAND2X0 P1_lt_178_U36 ( .IN1(P1_lt_178_n46), .IN2(P1_lt_178_n47), 
        .QN(P1_lt_178_n45) );
  NOR2X0 P1_lt_178_U35 ( .QN(P1_lt_178_n41), .IN1(P1_lt_178_n44), 
        .IN2(P1_lt_178_n45) );
  NOR2X0 P1_lt_178_U34 ( .QN(P1_lt_178_n42), .IN1(P1_N5107), 
        .IN2(P1_lt_178_n43) );
  NOR2X0 P1_lt_178_U33 ( .QN(P1_lt_178_n39), .IN1(P1_lt_178_n41), 
        .IN2(P1_lt_178_n42) );
  INVX0 P1_lt_178_U32 ( .ZN(P1_lt_178_n38), .INP(P1_N5423) );
  OR2X1 P1_lt_178_U31 ( .IN2(P1_N5108), .IN1(P1_lt_178_n38), .Q(P1_lt_178_n40)
         );
  NAND2X0 P1_lt_178_U30 ( .IN1(P1_lt_178_n39), .IN2(P1_lt_178_n40), 
        .QN(P1_lt_178_n36) );
  NAND2X0 P1_lt_178_U29 ( .IN1(P1_N5108), .IN2(P1_lt_178_n38), 
        .QN(P1_lt_178_n37) );
  NAND2X0 P1_lt_178_U28 ( .IN1(P1_lt_178_n36), .IN2(P1_lt_178_n37), 
        .QN(P1_lt_178_n35) );
  NOR2X0 P1_lt_178_U27 ( .QN(P1_lt_178_n31), .IN1(P1_lt_178_n34), 
        .IN2(P1_lt_178_n35) );
  NOR2X0 P1_lt_178_U26 ( .QN(P1_lt_178_n32), .IN1(P1_N5109), 
        .IN2(P1_lt_178_n33) );
  NOR2X0 P1_lt_178_U25 ( .QN(P1_lt_178_n29), .IN1(P1_lt_178_n31), 
        .IN2(P1_lt_178_n32) );
  INVX0 P1_lt_178_U24 ( .ZN(P1_lt_178_n28), .INP(P1_N5425) );
  OR2X1 P1_lt_178_U23 ( .IN2(P1_N5110), .IN1(P1_lt_178_n28), .Q(P1_lt_178_n30)
         );
  NAND2X0 P1_lt_178_U22 ( .IN1(P1_lt_178_n29), .IN2(P1_lt_178_n30), 
        .QN(P1_lt_178_n26) );
  NAND2X0 P1_lt_178_U21 ( .IN1(P1_N5110), .IN2(P1_lt_178_n28), 
        .QN(P1_lt_178_n27) );
  NAND2X0 P1_lt_178_U20 ( .IN1(P1_lt_178_n26), .IN2(P1_lt_178_n27), 
        .QN(P1_lt_178_n25) );
  NOR2X0 P1_lt_178_U19 ( .QN(P1_lt_178_n21), .IN1(P1_lt_178_n24), 
        .IN2(P1_lt_178_n25) );
  NOR2X0 P1_lt_178_U18 ( .QN(P1_lt_178_n22), .IN1(P1_N5111), 
        .IN2(P1_lt_178_n23) );
  NOR2X0 P1_lt_178_U17 ( .QN(P1_lt_178_n19), .IN1(P1_lt_178_n21), 
        .IN2(P1_lt_178_n22) );
  INVX0 P1_lt_178_U16 ( .ZN(P1_lt_178_n18), .INP(P1_N5427) );
  OR2X1 P1_lt_178_U15 ( .IN2(P1_N5112), .IN1(P1_lt_178_n18), .Q(P1_lt_178_n20)
         );
  NAND2X0 P1_lt_178_U14 ( .IN1(P1_lt_178_n19), .IN2(P1_lt_178_n20), 
        .QN(P1_lt_178_n16) );
  NAND2X0 P1_lt_178_U13 ( .IN1(P1_N5112), .IN2(P1_lt_178_n18), 
        .QN(P1_lt_178_n17) );
  NAND2X0 P1_lt_178_U12 ( .IN1(P1_lt_178_n16), .IN2(P1_lt_178_n17), 
        .QN(P1_lt_178_n15) );
  NOR2X0 P1_lt_178_U11 ( .QN(P1_lt_178_n11), .IN1(P1_lt_178_n14), 
        .IN2(P1_lt_178_n15) );
  NOR2X0 P1_lt_178_U10 ( .QN(P1_lt_178_n12), .IN1(P1_N5113), 
        .IN2(P1_lt_178_n13) );
  NOR2X0 P1_lt_178_U9 ( .QN(P1_lt_178_n9), .IN1(P1_lt_178_n11), 
        .IN2(P1_lt_178_n12) );
  INVX0 P1_lt_178_U8 ( .ZN(P1_lt_178_n8), .INP(P1_N5429) );
  OR2X1 P1_lt_178_U7 ( .IN2(P1_N5114), .IN1(P1_lt_178_n8), .Q(P1_lt_178_n10)
         );
  NAND2X0 P1_lt_178_U6 ( .IN1(P1_lt_178_n9), .IN2(P1_lt_178_n10), 
        .QN(P1_lt_178_n6) );
  NAND2X0 P1_lt_178_U5 ( .IN1(P1_N5114), .IN2(P1_lt_178_n8), .QN(P1_lt_178_n7)
         );
  NAND2X0 P1_lt_178_U4 ( .IN1(P1_lt_178_n6), .IN2(P1_lt_178_n7), 
        .QN(P1_lt_178_n3) );
  NAND2X0 P1_lt_178_U3 ( .IN1(P1_N5115), .IN2(P1_lt_178_n5), .QN(P1_lt_178_n4)
         );
  NAND2X0 P1_lt_178_U2 ( .IN1(P1_lt_178_n3), .IN2(P1_lt_178_n4), 
        .QN(P1_lt_178_n2) );
  NAND2X0 P1_lt_178_U1 ( .IN1(P1_lt_178_n1), .IN2(P1_lt_178_n2), .QN(P1_N5213)
         );
  INVX0 P1_lt_178_U151 ( .ZN(P1_lt_178_n33), .INP(P1_N5424) );
  AND2X1 P1_lt_178_U150 ( .IN1(P1_lt_178_n33), .IN2(P1_N5109), 
        .Q(P1_lt_178_n34) );
  INVX0 P1_lt_178_U149 ( .ZN(P1_lt_178_n43), .INP(P1_N5422) );
  AND2X1 P1_lt_178_U148 ( .IN1(P1_lt_178_n43), .IN2(P1_N5107), 
        .Q(P1_lt_178_n44) );
  INVX0 P1_lt_178_U147 ( .ZN(P1_lt_178_n53), .INP(P1_N5420) );
  AND2X1 P1_lt_178_U146 ( .IN1(P1_lt_178_n53), .IN2(P1_N5105), 
        .Q(P1_lt_178_n54) );
  INVX0 P1_lt_178_U145 ( .ZN(P1_lt_178_n63), .INP(P1_N5418) );
  AND2X1 P1_lt_178_U144 ( .IN1(P1_lt_178_n63), .IN2(P1_N5103), 
        .Q(P1_lt_178_n64) );
  INVX0 P1_lt_178_U143 ( .ZN(P1_lt_178_n73), .INP(P1_N5416) );
  AND2X1 P1_lt_178_U142 ( .IN1(P1_lt_178_n73), .IN2(P1_N5101), 
        .Q(P1_lt_178_n74) );
  INVX0 P1_lt_178_U141 ( .ZN(P1_lt_178_n83), .INP(P1_N5414) );
  AND2X1 P1_lt_178_U140 ( .IN1(P1_lt_178_n83), .IN2(P1_N5099), 
        .Q(P1_lt_178_n84) );
  INVX0 P1_lt_178_U139 ( .ZN(P1_lt_178_n93), .INP(P1_N5412) );
  AND2X1 P1_lt_178_U138 ( .IN1(P1_lt_178_n93), .IN2(P1_N5097), 
        .Q(P1_lt_178_n94) );
  INVX0 P1_lt_178_U137 ( .ZN(P1_lt_178_n103), .INP(P1_N5410) );
  AND2X1 P1_lt_178_U136 ( .IN1(P1_lt_178_n103), .IN2(P1_N5095), 
        .Q(P1_lt_178_n104) );
  NOR2X0 P1_lt_178_U134 ( .QN(P1_lt_178_n114), .IN1(P1_N5408), .IN2(n7273) );
  INVX0 P1_lt_178_U133 ( .ZN(P1_lt_178_n123), .INP(P1_N5406) );
  AND2X1 P1_lt_178_U132 ( .IN1(P1_lt_178_n123), .IN2(P1_N5091), 
        .Q(P1_lt_178_n124) );
  INVX0 P1_lt_178_U131 ( .ZN(P1_lt_178_n133), .INP(P1_N5404) );
  AND2X1 P1_lt_178_U130 ( .IN1(P1_lt_178_n133), .IN2(P1_N5089), 
        .Q(P1_lt_178_n134) );
  INVX0 P1_lt_178_U129 ( .ZN(P1_lt_178_n143), .INP(P1_N5402) );
  AND2X1 P1_lt_178_U128 ( .IN1(P1_lt_178_n143), .IN2(P1_N5087), 
        .Q(P1_lt_178_n144) );
  INVX0 P1_lt_178_U127 ( .ZN(P1_lt_178_n154), .INP(P1_N5400) );
  INVX0 P1_lt_178_U126 ( .ZN(P1_lt_178_n156), .INP(P1_N5084) );
  NOR2X0 P1_lt_178_U125 ( .QN(P1_lt_178_n153), .IN1(P1_lt_178_n156), 
        .IN2(P1_N5399) );
  AND2X1 P1_lt_178_U124 ( .IN1(P1_lt_178_n154), .IN2(P1_lt_178_n153), 
        .Q(P1_lt_178_n155) );
  NOR2X0 P1_lt_178_U123 ( .QN(P1_lt_178_n151), .IN1(P1_N5085), 
        .IN2(P1_lt_178_n155) );
  NOR2X0 P1_lt_178_U122 ( .QN(P1_lt_178_n152), .IN1(P1_lt_178_n153), 
        .IN2(P1_lt_178_n154) );
  NOR2X0 P1_lt_178_U121 ( .QN(P1_lt_178_n149), .IN1(P1_lt_178_n151), 
        .IN2(P1_lt_178_n152) );
  INVX0 P1_lt_178_U120 ( .ZN(P1_lt_178_n148), .INP(P1_N5401) );
  OR2X1 P1_lt_178_U119 ( .IN2(P1_N5086), .IN1(P1_lt_178_n148), 
        .Q(P1_lt_178_n150) );
  NAND2X0 P1_lt_178_U118 ( .IN1(P1_lt_178_n149), .IN2(P1_lt_178_n150), 
        .QN(P1_lt_178_n146) );
  NAND2X0 P1_lt_178_U117 ( .IN1(P1_N5086), .IN2(P1_lt_178_n148), 
        .QN(P1_lt_178_n147) );
  NAND2X0 P1_lt_178_U116 ( .IN1(P1_lt_178_n146), .IN2(P1_lt_178_n147), 
        .QN(P1_lt_178_n145) );
  NOR2X0 P1_lt_178_U115 ( .QN(P1_lt_178_n141), .IN1(P1_lt_178_n144), 
        .IN2(P1_lt_178_n145) );
  NOR2X0 P1_lt_178_U114 ( .QN(P1_lt_178_n142), .IN1(P1_N5087), 
        .IN2(P1_lt_178_n143) );
  NOR2X0 P1_lt_178_U113 ( .QN(P1_lt_178_n139), .IN1(P1_lt_178_n141), 
        .IN2(P1_lt_178_n142) );
  INVX0 P1_lt_178_U112 ( .ZN(P1_lt_178_n138), .INP(P1_N5403) );
  OR2X1 P1_lt_178_U111 ( .IN2(P1_N5088), .IN1(P1_lt_178_n138), 
        .Q(P1_lt_178_n140) );
  NAND2X0 P1_lt_178_U110 ( .IN1(P1_lt_178_n139), .IN2(P1_lt_178_n140), 
        .QN(P1_lt_178_n136) );
  NAND2X0 P1_lt_178_U109 ( .IN1(P1_N5088), .IN2(P1_lt_178_n138), 
        .QN(P1_lt_178_n137) );
  NAND2X0 P1_lt_178_U108 ( .IN1(P1_lt_178_n136), .IN2(P1_lt_178_n137), 
        .QN(P1_lt_178_n135) );
  NOR2X0 P1_lt_178_U107 ( .QN(P1_lt_178_n131), .IN1(P1_lt_178_n134), 
        .IN2(P1_lt_178_n135) );
  NOR2X0 P1_lt_178_U106 ( .QN(P1_lt_178_n132), .IN1(P1_N5089), 
        .IN2(P1_lt_178_n133) );
  NOR2X0 P1_lt_178_U105 ( .QN(P1_lt_178_n129), .IN1(P1_lt_178_n131), 
        .IN2(P1_lt_178_n132) );
  INVX0 P1_lt_178_U104 ( .ZN(P1_lt_178_n128), .INP(P1_N5405) );
  OR2X1 P1_lt_178_U103 ( .IN2(P1_N5090), .IN1(P1_lt_178_n128), 
        .Q(P1_lt_178_n130) );
  NAND2X0 P1_lt_178_U102 ( .IN1(P1_lt_178_n129), .IN2(P1_lt_178_n130), 
        .QN(P1_lt_178_n126) );
  NAND2X0 P1_lt_178_U101 ( .IN1(P1_N5090), .IN2(P1_lt_178_n128), 
        .QN(P1_lt_178_n127) );
  NAND2X0 P1_lt_178_U100 ( .IN1(P1_lt_178_n126), .IN2(P1_lt_178_n127), 
        .QN(P1_lt_178_n125) );
  NOR2X0 P1_lt_178_U99 ( .QN(P1_lt_178_n121), .IN1(P1_lt_178_n124), 
        .IN2(P1_lt_178_n125) );
  NOR2X0 P1_lt_178_U98 ( .QN(P1_lt_178_n122), .IN1(P1_N5091), 
        .IN2(P1_lt_178_n123) );
  NOR2X0 P1_lt_178_U97 ( .QN(P1_lt_178_n119), .IN1(P1_lt_178_n121), 
        .IN2(P1_lt_178_n122) );
  INVX0 P1_lt_178_U96 ( .ZN(P1_lt_178_n118), .INP(P1_N5407) );
  OR2X1 P1_lt_178_U95 ( .IN2(P1_N5092), .IN1(P1_lt_178_n118), 
        .Q(P1_lt_178_n120) );
  NAND2X0 P1_lt_178_U94 ( .IN1(P1_lt_178_n119), .IN2(P1_lt_178_n120), 
        .QN(P1_lt_178_n116) );
  NAND2X0 P1_lt_178_U93 ( .IN1(P1_N5092), .IN2(P1_lt_178_n118), 
        .QN(P1_lt_178_n117) );
  NAND2X0 P1_lt_178_U92 ( .IN1(P1_lt_178_n116), .IN2(P1_lt_178_n117), 
        .QN(P1_lt_178_n115) );
  NOR2X0 P1_lt_178_U91 ( .QN(P1_lt_178_n112), .IN1(P1_lt_178_n114), 
        .IN2(P1_lt_178_n115) );
  INVX0 P1_lt_178_U90 ( .ZN(P1_lt_178_n108), .INP(P1_N5409) );
  NOR2X0 P1_lt_178_U89 ( .QN(P1_lt_178_n113), .IN1(P1_N5094), 
        .IN2(P1_lt_178_n108) );
  NOR2X0 P1_lt_178_U88 ( .QN(P1_lt_178_n109), .IN1(P1_lt_178_n112), 
        .IN2(P1_lt_178_n113) );
  NAND2X0 P1_lt_178_U87 ( .IN1(P1_N5408), .IN2(n7273), .QN(P1_lt_178_n110) );
  NAND2X0 P1_lt_178_U86 ( .IN1(P1_lt_178_n109), .IN2(P1_lt_178_n110), 
        .QN(P1_lt_178_n106) );
  NAND2X0 P1_lt_178_U85 ( .IN1(P1_N5094), .IN2(P1_lt_178_n108), 
        .QN(P1_lt_178_n107) );
  NAND2X0 P1_lt_178_U84 ( .IN1(P1_lt_178_n106), .IN2(P1_lt_178_n107), 
        .QN(P1_lt_178_n105) );
  NOR2X0 P1_lt_178_U83 ( .QN(P1_lt_178_n101), .IN1(P1_lt_178_n104), 
        .IN2(P1_lt_178_n105) );
  NOR2X0 P1_lt_178_U82 ( .QN(P1_lt_178_n102), .IN1(P1_N5095), 
        .IN2(P1_lt_178_n103) );
  NOR2X0 P1_lt_178_U81 ( .QN(P1_lt_178_n99), .IN1(P1_lt_178_n101), 
        .IN2(P1_lt_178_n102) );
  INVX0 P1_lt_178_U80 ( .ZN(P1_lt_178_n98), .INP(P1_N5411) );
  OR2X1 P1_lt_178_U79 ( .IN2(P1_N5096), .IN1(P1_lt_178_n98), 
        .Q(P1_lt_178_n100) );
  NAND2X0 P1_lt_178_U78 ( .IN1(P1_lt_178_n99), .IN2(P1_lt_178_n100), 
        .QN(P1_lt_178_n96) );
  NAND2X0 P1_lt_178_U77 ( .IN1(P1_N5096), .IN2(P1_lt_178_n98), 
        .QN(P1_lt_178_n97) );
  NAND2X0 P1_lt_178_U76 ( .IN1(P1_lt_178_n96), .IN2(P1_lt_178_n97), 
        .QN(P1_lt_178_n95) );
  NOR2X0 P1_lt_178_U75 ( .QN(P1_lt_178_n91), .IN1(P1_lt_178_n94), 
        .IN2(P1_lt_178_n95) );
  NOR2X0 P1_lt_178_U74 ( .QN(P1_lt_178_n92), .IN1(P1_N5097), 
        .IN2(P1_lt_178_n93) );
  NOR2X0 P1_lt_178_U73 ( .QN(P1_lt_178_n89), .IN1(P1_lt_178_n91), 
        .IN2(P1_lt_178_n92) );
  INVX0 P1_lt_178_U72 ( .ZN(P1_lt_178_n88), .INP(P1_N5413) );
  OR2X1 P1_lt_178_U71 ( .IN2(P1_N5098), .IN1(P1_lt_178_n88), .Q(P1_lt_178_n90)
         );
  NAND2X0 P1_lt_178_U70 ( .IN1(P1_lt_178_n89), .IN2(P1_lt_178_n90), 
        .QN(P1_lt_178_n86) );
  NAND2X0 P1_lt_178_U69 ( .IN1(P1_N5098), .IN2(P1_lt_178_n88), 
        .QN(P1_lt_178_n87) );
  NAND2X0 P1_lt_178_U68 ( .IN1(P1_lt_178_n86), .IN2(P1_lt_178_n87), 
        .QN(P1_lt_178_n85) );
  NOR2X0 P1_lt_178_U67 ( .QN(P1_lt_178_n81), .IN1(P1_lt_178_n84), 
        .IN2(P1_lt_178_n85) );
  NOR2X0 P1_lt_178_U66 ( .QN(P1_lt_178_n82), .IN1(P1_N5099), 
        .IN2(P1_lt_178_n83) );
  NOR2X0 P1_lt_178_U65 ( .QN(P1_lt_178_n79), .IN1(P1_lt_178_n81), 
        .IN2(P1_lt_178_n82) );
  INVX0 P1_lt_178_U64 ( .ZN(P1_lt_178_n78), .INP(P1_N5415) );
  OR2X1 P1_lt_178_U63 ( .IN2(P1_N5100), .IN1(P1_lt_178_n78), .Q(P1_lt_178_n80)
         );
  NAND2X0 P1_lt_178_U62 ( .IN1(P1_lt_178_n79), .IN2(P1_lt_178_n80), 
        .QN(P1_lt_178_n76) );
  NAND2X0 P1_lt_178_U61 ( .IN1(P1_N5100), .IN2(P1_lt_178_n78), 
        .QN(P1_lt_178_n77) );
  NAND2X0 P1_lt_178_U60 ( .IN1(P1_lt_178_n76), .IN2(P1_lt_178_n77), 
        .QN(P1_lt_178_n75) );
  NOR2X0 P1_lt_178_U59 ( .QN(P1_lt_178_n71), .IN1(P1_lt_178_n74), 
        .IN2(P1_lt_178_n75) );
  INVX0 P1_lt_178_U157 ( .ZN(P1_lt_178_n5), .INP(P1_N5430) );
  OR2X1 P1_lt_178_U156 ( .IN2(P1_N5115), .IN1(P1_lt_178_n5), .Q(P1_lt_178_n1)
         );
  INVX0 P1_lt_178_U155 ( .ZN(P1_lt_178_n13), .INP(P1_N5428) );
  AND2X1 P1_lt_178_U154 ( .IN1(P1_lt_178_n13), .IN2(P1_N5113), 
        .Q(P1_lt_178_n14) );
  INVX0 P1_lt_178_U153 ( .ZN(P1_lt_178_n23), .INP(P1_N5426) );
  AND2X1 P1_lt_178_U152 ( .IN1(P1_lt_178_n23), .IN2(P1_N5111), 
        .Q(P1_lt_178_n24) );
  NAND2X0 P1_lt_186_U29 ( .IN1(P1_N5108), .IN2(P1_lt_186_n38), 
        .QN(P1_lt_186_n37) );
  NAND2X0 P1_lt_186_U28 ( .IN1(P1_lt_186_n36), .IN2(P1_lt_186_n37), 
        .QN(P1_lt_186_n35) );
  NOR2X0 P1_lt_186_U27 ( .QN(P1_lt_186_n31), .IN1(P1_lt_186_n34), 
        .IN2(P1_lt_186_n35) );
  NOR2X0 P1_lt_186_U26 ( .QN(P1_lt_186_n32), .IN1(P1_N5109), 
        .IN2(P1_lt_186_n33) );
  NOR2X0 P1_lt_186_U25 ( .QN(P1_lt_186_n29), .IN1(P1_lt_186_n31), 
        .IN2(P1_lt_186_n32) );
  INVX0 P1_lt_186_U24 ( .ZN(P1_lt_186_n28), .INP(P1_N5425) );
  OR2X1 P1_lt_186_U23 ( .IN2(P1_N5110), .IN1(P1_lt_186_n28), .Q(P1_lt_186_n30)
         );
  NAND2X0 P1_lt_186_U22 ( .IN1(P1_lt_186_n29), .IN2(P1_lt_186_n30), 
        .QN(P1_lt_186_n26) );
  NAND2X0 P1_lt_186_U21 ( .IN1(P1_N5110), .IN2(P1_lt_186_n28), 
        .QN(P1_lt_186_n27) );
  NAND2X0 P1_lt_186_U20 ( .IN1(P1_lt_186_n26), .IN2(P1_lt_186_n27), 
        .QN(P1_lt_186_n25) );
  NOR2X0 P1_lt_186_U19 ( .QN(P1_lt_186_n21), .IN1(P1_lt_186_n24), 
        .IN2(P1_lt_186_n25) );
  NOR2X0 P1_lt_186_U18 ( .QN(P1_lt_186_n22), .IN1(P1_N5111), 
        .IN2(P1_lt_186_n23) );
  NOR2X0 P1_lt_186_U17 ( .QN(P1_lt_186_n19), .IN1(P1_lt_186_n21), 
        .IN2(P1_lt_186_n22) );
  INVX0 P1_lt_186_U16 ( .ZN(P1_lt_186_n18), .INP(P1_N5427) );
  OR2X1 P1_lt_186_U15 ( .IN2(P1_N5112), .IN1(P1_lt_186_n18), .Q(P1_lt_186_n20)
         );
  NAND2X0 P1_lt_186_U14 ( .IN1(P1_lt_186_n19), .IN2(P1_lt_186_n20), 
        .QN(P1_lt_186_n16) );
  NAND2X0 P1_lt_186_U13 ( .IN1(P1_N5112), .IN2(P1_lt_186_n18), 
        .QN(P1_lt_186_n17) );
  NAND2X0 P1_lt_186_U12 ( .IN1(P1_lt_186_n16), .IN2(P1_lt_186_n17), 
        .QN(P1_lt_186_n15) );
  NOR2X0 P1_lt_186_U11 ( .QN(P1_lt_186_n11), .IN1(P1_lt_186_n14), 
        .IN2(P1_lt_186_n15) );
  NOR2X0 P1_lt_186_U10 ( .QN(P1_lt_186_n12), .IN1(P1_N5113), 
        .IN2(P1_lt_186_n13) );
  NOR2X0 P1_lt_186_U9 ( .QN(P1_lt_186_n9), .IN1(P1_lt_186_n11), 
        .IN2(P1_lt_186_n12) );
  INVX0 P1_lt_186_U8 ( .ZN(P1_lt_186_n8), .INP(P1_N5429) );
  OR2X1 P1_lt_186_U7 ( .IN2(P1_N5114), .IN1(P1_lt_186_n8), .Q(P1_lt_186_n10)
         );
  NAND2X0 P1_lt_186_U6 ( .IN1(P1_lt_186_n9), .IN2(P1_lt_186_n10), 
        .QN(P1_lt_186_n6) );
  NAND2X0 P1_lt_186_U5 ( .IN1(P1_N5114), .IN2(P1_lt_186_n8), .QN(P1_lt_186_n7)
         );
  NAND2X0 P1_lt_186_U4 ( .IN1(P1_lt_186_n6), .IN2(P1_lt_186_n7), 
        .QN(P1_lt_186_n3) );
  NAND2X0 P1_lt_186_U3 ( .IN1(P1_N5115), .IN2(P1_lt_186_n5), .QN(P1_lt_186_n4)
         );
  NAND2X0 P1_lt_186_U2 ( .IN1(P1_lt_186_n3), .IN2(P1_lt_186_n4), 
        .QN(P1_lt_186_n2) );
  NAND2X0 P1_lt_186_U1 ( .IN1(P1_lt_186_n1), .IN2(P1_lt_186_n2), .QN(P1_N5281)
         );
  NOR2X0 P1_lt_186_U122 ( .QN(P1_lt_186_n152), .IN1(P1_lt_186_n153), 
        .IN2(P1_lt_186_n154) );
  NOR2X0 P1_lt_186_U121 ( .QN(P1_lt_186_n149), .IN1(P1_lt_186_n151), 
        .IN2(P1_lt_186_n152) );
  INVX0 P1_lt_186_U120 ( .ZN(P1_lt_186_n148), .INP(P1_N5401) );
  OR2X1 P1_lt_186_U119 ( .IN2(P1_N5086), .IN1(P1_lt_186_n148), 
        .Q(P1_lt_186_n150) );
  NAND2X0 P1_lt_186_U118 ( .IN1(P1_lt_186_n149), .IN2(P1_lt_186_n150), 
        .QN(P1_lt_186_n146) );
  NAND2X0 P1_lt_186_U117 ( .IN1(P1_N5086), .IN2(P1_lt_186_n148), 
        .QN(P1_lt_186_n147) );
  NAND2X0 P1_lt_186_U116 ( .IN1(P1_lt_186_n146), .IN2(P1_lt_186_n147), 
        .QN(P1_lt_186_n145) );
  NOR2X0 P1_lt_186_U115 ( .QN(P1_lt_186_n141), .IN1(P1_lt_186_n144), 
        .IN2(P1_lt_186_n145) );
  NOR2X0 P1_lt_186_U114 ( .QN(P1_lt_186_n142), .IN1(P1_N5087), 
        .IN2(P1_lt_186_n143) );
  NOR2X0 P1_lt_186_U113 ( .QN(P1_lt_186_n139), .IN1(P1_lt_186_n141), 
        .IN2(P1_lt_186_n142) );
  INVX0 P1_lt_186_U112 ( .ZN(P1_lt_186_n138), .INP(P1_N5403) );
  OR2X1 P1_lt_186_U111 ( .IN2(P1_N5088), .IN1(P1_lt_186_n138), 
        .Q(P1_lt_186_n140) );
  NAND2X0 P1_lt_186_U110 ( .IN1(P1_lt_186_n139), .IN2(P1_lt_186_n140), 
        .QN(P1_lt_186_n136) );
  NAND2X0 P1_lt_186_U109 ( .IN1(P1_N5088), .IN2(P1_lt_186_n138), 
        .QN(P1_lt_186_n137) );
  NAND2X0 P1_lt_186_U108 ( .IN1(P1_lt_186_n136), .IN2(P1_lt_186_n137), 
        .QN(P1_lt_186_n135) );
  NOR2X0 P1_lt_186_U107 ( .QN(P1_lt_186_n131), .IN1(P1_lt_186_n134), 
        .IN2(P1_lt_186_n135) );
  NOR2X0 P1_lt_186_U106 ( .QN(P1_lt_186_n132), .IN1(P1_N5089), 
        .IN2(P1_lt_186_n133) );
  NOR2X0 P1_lt_186_U105 ( .QN(P1_lt_186_n129), .IN1(P1_lt_186_n131), 
        .IN2(P1_lt_186_n132) );
  INVX0 P1_lt_186_U104 ( .ZN(P1_lt_186_n128), .INP(P1_N5405) );
  OR2X1 P1_lt_186_U103 ( .IN2(P1_N5090), .IN1(P1_lt_186_n128), 
        .Q(P1_lt_186_n130) );
  NAND2X0 P1_lt_186_U102 ( .IN1(P1_lt_186_n129), .IN2(P1_lt_186_n130), 
        .QN(P1_lt_186_n126) );
  NAND2X0 P1_lt_186_U101 ( .IN1(P1_N5090), .IN2(P1_lt_186_n128), 
        .QN(P1_lt_186_n127) );
  NAND2X0 P1_lt_186_U100 ( .IN1(P1_lt_186_n126), .IN2(P1_lt_186_n127), 
        .QN(P1_lt_186_n125) );
  NOR2X0 P1_lt_186_U99 ( .QN(P1_lt_186_n121), .IN1(P1_lt_186_n124), 
        .IN2(P1_lt_186_n125) );
  NOR2X0 P1_lt_186_U98 ( .QN(P1_lt_186_n122), .IN1(P1_N5091), 
        .IN2(P1_lt_186_n123) );
  NOR2X0 P1_lt_186_U97 ( .QN(P1_lt_186_n119), .IN1(P1_lt_186_n121), 
        .IN2(P1_lt_186_n122) );
  INVX0 P1_lt_186_U96 ( .ZN(P1_lt_186_n118), .INP(P1_N5407) );
  OR2X1 P1_lt_186_U95 ( .IN2(P1_N5092), .IN1(P1_lt_186_n118), 
        .Q(P1_lt_186_n120) );
  NAND2X0 P1_lt_186_U94 ( .IN1(P1_lt_186_n119), .IN2(P1_lt_186_n120), 
        .QN(P1_lt_186_n116) );
  NAND2X0 P1_lt_186_U93 ( .IN1(P1_N5092), .IN2(P1_lt_186_n118), 
        .QN(P1_lt_186_n117) );
  NAND2X0 P1_lt_186_U92 ( .IN1(P1_lt_186_n116), .IN2(P1_lt_186_n117), 
        .QN(P1_lt_186_n115) );
  NOR2X0 P1_lt_186_U91 ( .QN(P1_lt_186_n112), .IN1(P1_lt_186_n114), 
        .IN2(P1_lt_186_n115) );
  INVX0 P1_lt_186_U90 ( .ZN(P1_lt_186_n108), .INP(P1_N5409) );
  NOR2X0 P1_lt_186_U89 ( .QN(P1_lt_186_n113), .IN1(P1_N5094), 
        .IN2(P1_lt_186_n108) );
  NOR2X0 P1_lt_186_U88 ( .QN(P1_lt_186_n109), .IN1(P1_lt_186_n112), 
        .IN2(P1_lt_186_n113) );
  NAND2X0 P1_lt_186_U87 ( .IN1(P1_N5408), .IN2(n7273), .QN(P1_lt_186_n110) );
  NAND2X0 P1_lt_186_U86 ( .IN1(P1_lt_186_n109), .IN2(P1_lt_186_n110), 
        .QN(P1_lt_186_n106) );
  NAND2X0 P1_lt_186_U85 ( .IN1(P1_N5094), .IN2(P1_lt_186_n108), 
        .QN(P1_lt_186_n107) );
  NAND2X0 P1_lt_186_U84 ( .IN1(P1_lt_186_n106), .IN2(P1_lt_186_n107), 
        .QN(P1_lt_186_n105) );
  NOR2X0 P1_lt_186_U83 ( .QN(P1_lt_186_n101), .IN1(P1_lt_186_n104), 
        .IN2(P1_lt_186_n105) );
  NOR2X0 P1_lt_186_U82 ( .QN(P1_lt_186_n102), .IN1(P1_N5095), 
        .IN2(P1_lt_186_n103) );
  NOR2X0 P1_lt_186_U81 ( .QN(P1_lt_186_n99), .IN1(P1_lt_186_n101), 
        .IN2(P1_lt_186_n102) );
  INVX0 P1_lt_186_U80 ( .ZN(P1_lt_186_n98), .INP(P1_N5411) );
  OR2X1 P1_lt_186_U79 ( .IN2(P1_N5096), .IN1(P1_lt_186_n98), 
        .Q(P1_lt_186_n100) );
  NAND2X0 P1_lt_186_U78 ( .IN1(P1_lt_186_n99), .IN2(P1_lt_186_n100), 
        .QN(P1_lt_186_n96) );
  NAND2X0 P1_lt_186_U77 ( .IN1(P1_N5096), .IN2(P1_lt_186_n98), 
        .QN(P1_lt_186_n97) );
  NAND2X0 P1_lt_186_U76 ( .IN1(P1_lt_186_n96), .IN2(P1_lt_186_n97), 
        .QN(P1_lt_186_n95) );
  NOR2X0 P1_lt_186_U75 ( .QN(P1_lt_186_n91), .IN1(P1_lt_186_n94), 
        .IN2(P1_lt_186_n95) );
  NOR2X0 P1_lt_186_U74 ( .QN(P1_lt_186_n92), .IN1(P1_N5097), 
        .IN2(P1_lt_186_n93) );
  NOR2X0 P1_lt_186_U73 ( .QN(P1_lt_186_n89), .IN1(P1_lt_186_n91), 
        .IN2(P1_lt_186_n92) );
  INVX0 P1_lt_186_U72 ( .ZN(P1_lt_186_n88), .INP(P1_N5413) );
  OR2X1 P1_lt_186_U71 ( .IN2(P1_N5098), .IN1(P1_lt_186_n88), .Q(P1_lt_186_n90)
         );
  NAND2X0 P1_lt_186_U70 ( .IN1(P1_lt_186_n89), .IN2(P1_lt_186_n90), 
        .QN(P1_lt_186_n86) );
  NAND2X0 P1_lt_186_U69 ( .IN1(P1_N5098), .IN2(P1_lt_186_n88), 
        .QN(P1_lt_186_n87) );
  NAND2X0 P1_lt_186_U68 ( .IN1(P1_lt_186_n86), .IN2(P1_lt_186_n87), 
        .QN(P1_lt_186_n85) );
  NOR2X0 P1_lt_186_U67 ( .QN(P1_lt_186_n81), .IN1(P1_lt_186_n84), 
        .IN2(P1_lt_186_n85) );
  NOR2X0 P1_lt_186_U66 ( .QN(P1_lt_186_n82), .IN1(P1_N5099), 
        .IN2(P1_lt_186_n83) );
  NOR2X0 P1_lt_186_U65 ( .QN(P1_lt_186_n79), .IN1(P1_lt_186_n81), 
        .IN2(P1_lt_186_n82) );
  INVX0 P1_lt_186_U64 ( .ZN(P1_lt_186_n78), .INP(P1_N5415) );
  OR2X1 P1_lt_186_U63 ( .IN2(P1_N5100), .IN1(P1_lt_186_n78), .Q(P1_lt_186_n80)
         );
  NAND2X0 P1_lt_186_U62 ( .IN1(P1_lt_186_n79), .IN2(P1_lt_186_n80), 
        .QN(P1_lt_186_n76) );
  NAND2X0 P1_lt_186_U61 ( .IN1(P1_N5100), .IN2(P1_lt_186_n78), 
        .QN(P1_lt_186_n77) );
  NAND2X0 P1_lt_186_U60 ( .IN1(P1_lt_186_n76), .IN2(P1_lt_186_n77), 
        .QN(P1_lt_186_n75) );
  NOR2X0 P1_lt_186_U59 ( .QN(P1_lt_186_n71), .IN1(P1_lt_186_n74), 
        .IN2(P1_lt_186_n75) );
  NOR2X0 P1_lt_186_U58 ( .QN(P1_lt_186_n72), .IN1(P1_N5101), 
        .IN2(P1_lt_186_n73) );
  NOR2X0 P1_lt_186_U57 ( .QN(P1_lt_186_n69), .IN1(P1_lt_186_n71), 
        .IN2(P1_lt_186_n72) );
  INVX0 P1_lt_186_U56 ( .ZN(P1_lt_186_n68), .INP(P1_N5417) );
  OR2X1 P1_lt_186_U55 ( .IN2(P1_N5102), .IN1(P1_lt_186_n68), .Q(P1_lt_186_n70)
         );
  NAND2X0 P1_lt_186_U54 ( .IN1(P1_lt_186_n69), .IN2(P1_lt_186_n70), 
        .QN(P1_lt_186_n66) );
  NAND2X0 P1_lt_186_U53 ( .IN1(P1_N5102), .IN2(P1_lt_186_n68), 
        .QN(P1_lt_186_n67) );
  NAND2X0 P1_lt_186_U52 ( .IN1(P1_lt_186_n66), .IN2(P1_lt_186_n67), 
        .QN(P1_lt_186_n65) );
  NOR2X0 P1_lt_186_U51 ( .QN(P1_lt_186_n61), .IN1(P1_lt_186_n64), 
        .IN2(P1_lt_186_n65) );
  NOR2X0 P1_lt_186_U50 ( .QN(P1_lt_186_n62), .IN1(P1_N5103), 
        .IN2(P1_lt_186_n63) );
  NOR2X0 P1_lt_186_U49 ( .QN(P1_lt_186_n59), .IN1(P1_lt_186_n61), 
        .IN2(P1_lt_186_n62) );
  INVX0 P1_lt_186_U48 ( .ZN(P1_lt_186_n58), .INP(P1_N5419) );
  OR2X1 P1_lt_186_U47 ( .IN2(P1_N5104), .IN1(P1_lt_186_n58), .Q(P1_lt_186_n60)
         );
  NAND2X0 P1_lt_186_U46 ( .IN1(P1_lt_186_n59), .IN2(P1_lt_186_n60), 
        .QN(P1_lt_186_n56) );
  NAND2X0 P1_lt_186_U45 ( .IN1(P1_N5104), .IN2(P1_lt_186_n58), 
        .QN(P1_lt_186_n57) );
  NAND2X0 P1_lt_186_U44 ( .IN1(P1_lt_186_n56), .IN2(P1_lt_186_n57), 
        .QN(P1_lt_186_n55) );
  NOR2X0 P1_lt_186_U43 ( .QN(P1_lt_186_n51), .IN1(P1_lt_186_n54), 
        .IN2(P1_lt_186_n55) );
  NOR2X0 P1_lt_186_U42 ( .QN(P1_lt_186_n52), .IN1(P1_N5105), 
        .IN2(P1_lt_186_n53) );
  NOR2X0 P1_lt_186_U41 ( .QN(P1_lt_186_n49), .IN1(P1_lt_186_n51), 
        .IN2(P1_lt_186_n52) );
  INVX0 P1_lt_186_U40 ( .ZN(P1_lt_186_n48), .INP(P1_N5421) );
  OR2X1 P1_lt_186_U39 ( .IN2(P1_N5106), .IN1(P1_lt_186_n48), .Q(P1_lt_186_n50)
         );
  NAND2X0 P1_lt_186_U38 ( .IN1(P1_lt_186_n49), .IN2(P1_lt_186_n50), 
        .QN(P1_lt_186_n46) );
  NAND2X0 P1_lt_186_U37 ( .IN1(P1_N5106), .IN2(P1_lt_186_n48), 
        .QN(P1_lt_186_n47) );
  NAND2X0 P1_lt_186_U36 ( .IN1(P1_lt_186_n46), .IN2(P1_lt_186_n47), 
        .QN(P1_lt_186_n45) );
  NOR2X0 P1_lt_186_U35 ( .QN(P1_lt_186_n41), .IN1(P1_lt_186_n44), 
        .IN2(P1_lt_186_n45) );
  NOR2X0 P1_lt_186_U34 ( .QN(P1_lt_186_n42), .IN1(P1_N5107), 
        .IN2(P1_lt_186_n43) );
  NOR2X0 P1_lt_186_U33 ( .QN(P1_lt_186_n39), .IN1(P1_lt_186_n41), 
        .IN2(P1_lt_186_n42) );
  INVX0 P1_lt_186_U32 ( .ZN(P1_lt_186_n38), .INP(P1_N5423) );
  OR2X1 P1_lt_186_U31 ( .IN2(P1_N5108), .IN1(P1_lt_186_n38), .Q(P1_lt_186_n40)
         );
  NAND2X0 P1_lt_186_U30 ( .IN1(P1_lt_186_n39), .IN2(P1_lt_186_n40), 
        .QN(P1_lt_186_n36) );
  INVX0 P1_lt_186_U157 ( .ZN(P1_lt_186_n5), .INP(P1_N5430) );
  OR2X1 P1_lt_186_U156 ( .IN2(P1_N5115), .IN1(P1_lt_186_n5), .Q(P1_lt_186_n1)
         );
  INVX0 P1_lt_186_U155 ( .ZN(P1_lt_186_n13), .INP(P1_N5428) );
  AND2X1 P1_lt_186_U154 ( .IN1(P1_lt_186_n13), .IN2(P1_N5113), 
        .Q(P1_lt_186_n14) );
  INVX0 P1_lt_186_U153 ( .ZN(P1_lt_186_n23), .INP(P1_N5426) );
  AND2X1 P1_lt_186_U152 ( .IN1(P1_lt_186_n23), .IN2(P1_N5111), 
        .Q(P1_lt_186_n24) );
  INVX0 P1_lt_186_U151 ( .ZN(P1_lt_186_n33), .INP(P1_N5424) );
  AND2X1 P1_lt_186_U150 ( .IN1(P1_lt_186_n33), .IN2(P1_N5109), 
        .Q(P1_lt_186_n34) );
  INVX0 P1_lt_186_U149 ( .ZN(P1_lt_186_n43), .INP(P1_N5422) );
  AND2X1 P1_lt_186_U148 ( .IN1(P1_lt_186_n43), .IN2(P1_N5107), 
        .Q(P1_lt_186_n44) );
  INVX0 P1_lt_186_U147 ( .ZN(P1_lt_186_n53), .INP(P1_N5420) );
  AND2X1 P1_lt_186_U146 ( .IN1(P1_lt_186_n53), .IN2(P1_N5105), 
        .Q(P1_lt_186_n54) );
  INVX0 P1_lt_186_U145 ( .ZN(P1_lt_186_n63), .INP(P1_N5418) );
  AND2X1 P1_lt_186_U144 ( .IN1(P1_lt_186_n63), .IN2(P1_N5103), 
        .Q(P1_lt_186_n64) );
  INVX0 P1_lt_186_U143 ( .ZN(P1_lt_186_n73), .INP(P1_N5416) );
  AND2X1 P1_lt_186_U142 ( .IN1(P1_lt_186_n73), .IN2(P1_N5101), 
        .Q(P1_lt_186_n74) );
  INVX0 P1_lt_186_U141 ( .ZN(P1_lt_186_n83), .INP(P1_N5414) );
  AND2X1 P1_lt_186_U140 ( .IN1(P1_lt_186_n83), .IN2(P1_N5099), 
        .Q(P1_lt_186_n84) );
  INVX0 P1_lt_186_U139 ( .ZN(P1_lt_186_n93), .INP(P1_N5412) );
  AND2X1 P1_lt_186_U138 ( .IN1(P1_lt_186_n93), .IN2(P1_N5097), 
        .Q(P1_lt_186_n94) );
  INVX0 P1_lt_186_U137 ( .ZN(P1_lt_186_n103), .INP(P1_N5410) );
  AND2X1 P1_lt_186_U136 ( .IN1(P1_lt_186_n103), .IN2(P1_N5095), 
        .Q(P1_lt_186_n104) );
  NOR2X0 P1_lt_186_U134 ( .QN(P1_lt_186_n114), .IN1(P1_N5408), .IN2(n7273) );
  INVX0 P1_lt_186_U133 ( .ZN(P1_lt_186_n123), .INP(P1_N5406) );
  AND2X1 P1_lt_186_U132 ( .IN1(P1_lt_186_n123), .IN2(P1_N5091), 
        .Q(P1_lt_186_n124) );
  INVX0 P1_lt_186_U131 ( .ZN(P1_lt_186_n133), .INP(P1_N5404) );
  AND2X1 P1_lt_186_U130 ( .IN1(P1_lt_186_n133), .IN2(P1_N5089), 
        .Q(P1_lt_186_n134) );
  INVX0 P1_lt_186_U129 ( .ZN(P1_lt_186_n143), .INP(P1_N5402) );
  AND2X1 P1_lt_186_U128 ( .IN1(P1_lt_186_n143), .IN2(P1_N5087), 
        .Q(P1_lt_186_n144) );
  INVX0 P1_lt_186_U127 ( .ZN(P1_lt_186_n154), .INP(P1_N5400) );
  INVX0 P1_lt_186_U126 ( .ZN(P1_lt_186_n156), .INP(P1_N5084) );
  NOR2X0 P1_lt_186_U125 ( .QN(P1_lt_186_n153), .IN1(P1_lt_186_n156), 
        .IN2(P1_N5399) );
  AND2X1 P1_lt_186_U124 ( .IN1(P1_lt_186_n154), .IN2(P1_lt_186_n153), 
        .Q(P1_lt_186_n155) );
  NOR2X0 P1_lt_186_U123 ( .QN(P1_lt_186_n151), .IN1(P1_N5085), 
        .IN2(P1_lt_186_n155) );
  NAND2X0 P1_lt_224_U93 ( .IN1(P1_N5092), .IN2(P1_lt_224_n118), 
        .QN(P1_lt_224_n117) );
  NAND2X0 P1_lt_224_U92 ( .IN1(P1_lt_224_n116), .IN2(P1_lt_224_n117), 
        .QN(P1_lt_224_n115) );
  NOR2X0 P1_lt_224_U91 ( .QN(P1_lt_224_n112), .IN1(P1_lt_224_n114), 
        .IN2(P1_lt_224_n115) );
  INVX0 P1_lt_224_U90 ( .ZN(P1_lt_224_n108), .INP(P1_N5409) );
  NOR2X0 P1_lt_224_U89 ( .QN(P1_lt_224_n113), .IN1(P1_N5094), 
        .IN2(P1_lt_224_n108) );
  NOR2X0 P1_lt_224_U88 ( .QN(P1_lt_224_n109), .IN1(P1_lt_224_n112), 
        .IN2(P1_lt_224_n113) );
  NAND2X0 P1_lt_224_U87 ( .IN1(P1_N5408), .IN2(n7273), .QN(P1_lt_224_n110) );
  NAND2X0 P1_lt_224_U86 ( .IN1(P1_lt_224_n109), .IN2(P1_lt_224_n110), 
        .QN(P1_lt_224_n106) );
  NAND2X0 P1_lt_224_U85 ( .IN1(P1_N5094), .IN2(P1_lt_224_n108), 
        .QN(P1_lt_224_n107) );
  NAND2X0 P1_lt_224_U84 ( .IN1(P1_lt_224_n106), .IN2(P1_lt_224_n107), 
        .QN(P1_lt_224_n105) );
  NOR2X0 P1_lt_224_U83 ( .QN(P1_lt_224_n101), .IN1(P1_lt_224_n104), 
        .IN2(P1_lt_224_n105) );
  NOR2X0 P1_lt_224_U82 ( .QN(P1_lt_224_n102), .IN1(P1_N5095), 
        .IN2(P1_lt_224_n103) );
  NOR2X0 P1_lt_224_U81 ( .QN(P1_lt_224_n99), .IN1(P1_lt_224_n101), 
        .IN2(P1_lt_224_n102) );
  INVX0 P1_lt_224_U80 ( .ZN(P1_lt_224_n98), .INP(P1_N5411) );
  OR2X1 P1_lt_224_U79 ( .IN2(P1_N5096), .IN1(P1_lt_224_n98), 
        .Q(P1_lt_224_n100) );
  NAND2X0 P1_lt_224_U78 ( .IN1(P1_lt_224_n99), .IN2(P1_lt_224_n100), 
        .QN(P1_lt_224_n96) );
  NAND2X0 P1_lt_224_U77 ( .IN1(P1_N5096), .IN2(P1_lt_224_n98), 
        .QN(P1_lt_224_n97) );
  NAND2X0 P1_lt_224_U76 ( .IN1(P1_lt_224_n96), .IN2(P1_lt_224_n97), 
        .QN(P1_lt_224_n95) );
  NOR2X0 P1_lt_224_U75 ( .QN(P1_lt_224_n91), .IN1(P1_lt_224_n94), 
        .IN2(P1_lt_224_n95) );
  NOR2X0 P1_lt_224_U74 ( .QN(P1_lt_224_n92), .IN1(P1_N5097), 
        .IN2(P1_lt_224_n93) );
  NOR2X0 P1_lt_224_U73 ( .QN(P1_lt_224_n89), .IN1(P1_lt_224_n91), 
        .IN2(P1_lt_224_n92) );
  INVX0 P1_lt_224_U72 ( .ZN(P1_lt_224_n88), .INP(P1_N5413) );
  OR2X1 P1_lt_224_U71 ( .IN2(P1_N5098), .IN1(P1_lt_224_n88), .Q(P1_lt_224_n90)
         );
  NAND2X0 P1_lt_224_U70 ( .IN1(P1_lt_224_n89), .IN2(P1_lt_224_n90), 
        .QN(P1_lt_224_n86) );
  NAND2X0 P1_lt_224_U69 ( .IN1(P1_N5098), .IN2(P1_lt_224_n88), 
        .QN(P1_lt_224_n87) );
  NAND2X0 P1_lt_224_U68 ( .IN1(P1_lt_224_n86), .IN2(P1_lt_224_n87), 
        .QN(P1_lt_224_n85) );
  NOR2X0 P1_lt_224_U67 ( .QN(P1_lt_224_n81), .IN1(P1_lt_224_n84), 
        .IN2(P1_lt_224_n85) );
  NOR2X0 P1_lt_224_U66 ( .QN(P1_lt_224_n82), .IN1(P1_N5099), 
        .IN2(P1_lt_224_n83) );
  NOR2X0 P1_lt_224_U65 ( .QN(P1_lt_224_n79), .IN1(P1_lt_224_n81), 
        .IN2(P1_lt_224_n82) );
  INVX0 P1_lt_224_U64 ( .ZN(P1_lt_224_n78), .INP(P1_N5415) );
  OR2X1 P1_lt_224_U63 ( .IN2(P1_N5100), .IN1(P1_lt_224_n78), .Q(P1_lt_224_n80)
         );
  NAND2X0 P1_lt_224_U62 ( .IN1(P1_lt_224_n79), .IN2(P1_lt_224_n80), 
        .QN(P1_lt_224_n76) );
  NAND2X0 P1_lt_224_U61 ( .IN1(P1_N5100), .IN2(P1_lt_224_n78), 
        .QN(P1_lt_224_n77) );
  NAND2X0 P1_lt_224_U60 ( .IN1(P1_lt_224_n76), .IN2(P1_lt_224_n77), 
        .QN(P1_lt_224_n75) );
  NOR2X0 P1_lt_224_U59 ( .QN(P1_lt_224_n71), .IN1(P1_lt_224_n74), 
        .IN2(P1_lt_224_n75) );
  NOR2X0 P1_lt_224_U58 ( .QN(P1_lt_224_n72), .IN1(P1_N5101), 
        .IN2(P1_lt_224_n73) );
  NOR2X0 P1_lt_224_U57 ( .QN(P1_lt_224_n69), .IN1(P1_lt_224_n71), 
        .IN2(P1_lt_224_n72) );
  INVX0 P1_lt_224_U56 ( .ZN(P1_lt_224_n68), .INP(P1_N5417) );
  OR2X1 P1_lt_224_U55 ( .IN2(P1_N5102), .IN1(P1_lt_224_n68), .Q(P1_lt_224_n70)
         );
  NAND2X0 P1_lt_224_U54 ( .IN1(P1_lt_224_n69), .IN2(P1_lt_224_n70), 
        .QN(P1_lt_224_n66) );
  NAND2X0 P1_lt_224_U53 ( .IN1(P1_N5102), .IN2(P1_lt_224_n68), 
        .QN(P1_lt_224_n67) );
  NAND2X0 P1_lt_224_U52 ( .IN1(P1_lt_224_n66), .IN2(P1_lt_224_n67), 
        .QN(P1_lt_224_n65) );
  NOR2X0 P1_lt_224_U51 ( .QN(P1_lt_224_n61), .IN1(P1_lt_224_n64), 
        .IN2(P1_lt_224_n65) );
  NOR2X0 P1_lt_224_U50 ( .QN(P1_lt_224_n62), .IN1(P1_N5103), 
        .IN2(P1_lt_224_n63) );
  NOR2X0 P1_lt_224_U49 ( .QN(P1_lt_224_n59), .IN1(P1_lt_224_n61), 
        .IN2(P1_lt_224_n62) );
  INVX0 P1_lt_224_U48 ( .ZN(P1_lt_224_n58), .INP(P1_N5419) );
  OR2X1 P1_lt_224_U47 ( .IN2(P1_N5104), .IN1(P1_lt_224_n58), .Q(P1_lt_224_n60)
         );
  NAND2X0 P1_lt_224_U46 ( .IN1(P1_lt_224_n59), .IN2(P1_lt_224_n60), 
        .QN(P1_lt_224_n56) );
  NAND2X0 P1_lt_224_U45 ( .IN1(P1_N5104), .IN2(P1_lt_224_n58), 
        .QN(P1_lt_224_n57) );
  NAND2X0 P1_lt_224_U44 ( .IN1(P1_lt_224_n56), .IN2(P1_lt_224_n57), 
        .QN(P1_lt_224_n55) );
  NOR2X0 P1_lt_224_U43 ( .QN(P1_lt_224_n51), .IN1(P1_lt_224_n54), 
        .IN2(P1_lt_224_n55) );
  NOR2X0 P1_lt_224_U42 ( .QN(P1_lt_224_n52), .IN1(P1_N5105), 
        .IN2(P1_lt_224_n53) );
  NOR2X0 P1_lt_224_U41 ( .QN(P1_lt_224_n49), .IN1(P1_lt_224_n51), 
        .IN2(P1_lt_224_n52) );
  INVX0 P1_lt_224_U40 ( .ZN(P1_lt_224_n48), .INP(P1_N5421) );
  OR2X1 P1_lt_224_U39 ( .IN2(P1_N5106), .IN1(P1_lt_224_n48), .Q(P1_lt_224_n50)
         );
  NAND2X0 P1_lt_224_U38 ( .IN1(P1_lt_224_n49), .IN2(P1_lt_224_n50), 
        .QN(P1_lt_224_n46) );
  NAND2X0 P1_lt_224_U37 ( .IN1(P1_N5106), .IN2(P1_lt_224_n48), 
        .QN(P1_lt_224_n47) );
  NAND2X0 P1_lt_224_U36 ( .IN1(P1_lt_224_n46), .IN2(P1_lt_224_n47), 
        .QN(P1_lt_224_n45) );
  NOR2X0 P1_lt_224_U35 ( .QN(P1_lt_224_n41), .IN1(P1_lt_224_n44), 
        .IN2(P1_lt_224_n45) );
  NOR2X0 P1_lt_224_U34 ( .QN(P1_lt_224_n42), .IN1(P1_N5107), 
        .IN2(P1_lt_224_n43) );
  NOR2X0 P1_lt_224_U33 ( .QN(P1_lt_224_n39), .IN1(P1_lt_224_n41), 
        .IN2(P1_lt_224_n42) );
  INVX0 P1_lt_224_U32 ( .ZN(P1_lt_224_n38), .INP(P1_N5423) );
  OR2X1 P1_lt_224_U31 ( .IN2(P1_N5108), .IN1(P1_lt_224_n38), .Q(P1_lt_224_n40)
         );
  NAND2X0 P1_lt_224_U30 ( .IN1(P1_lt_224_n39), .IN2(P1_lt_224_n40), 
        .QN(P1_lt_224_n36) );
  NAND2X0 P1_lt_224_U29 ( .IN1(P1_N5108), .IN2(P1_lt_224_n38), 
        .QN(P1_lt_224_n37) );
  NAND2X0 P1_lt_224_U28 ( .IN1(P1_lt_224_n36), .IN2(P1_lt_224_n37), 
        .QN(P1_lt_224_n35) );
  NOR2X0 P1_lt_224_U27 ( .QN(P1_lt_224_n31), .IN1(P1_lt_224_n34), 
        .IN2(P1_lt_224_n35) );
  NOR2X0 P1_lt_224_U26 ( .QN(P1_lt_224_n32), .IN1(P1_N5109), 
        .IN2(P1_lt_224_n33) );
  NOR2X0 P1_lt_224_U25 ( .QN(P1_lt_224_n29), .IN1(P1_lt_224_n31), 
        .IN2(P1_lt_224_n32) );
  INVX0 P1_lt_224_U24 ( .ZN(P1_lt_224_n28), .INP(P1_N5425) );
  OR2X1 P1_lt_224_U23 ( .IN2(P1_N5110), .IN1(P1_lt_224_n28), .Q(P1_lt_224_n30)
         );
  NAND2X0 P1_lt_224_U22 ( .IN1(P1_lt_224_n29), .IN2(P1_lt_224_n30), 
        .QN(P1_lt_224_n26) );
  NAND2X0 P1_lt_224_U21 ( .IN1(P1_N5110), .IN2(P1_lt_224_n28), 
        .QN(P1_lt_224_n27) );
  NAND2X0 P1_lt_224_U20 ( .IN1(P1_lt_224_n26), .IN2(P1_lt_224_n27), 
        .QN(P1_lt_224_n25) );
  NOR2X0 P1_lt_224_U19 ( .QN(P1_lt_224_n21), .IN1(P1_lt_224_n24), 
        .IN2(P1_lt_224_n25) );
  NOR2X0 P1_lt_224_U18 ( .QN(P1_lt_224_n22), .IN1(P1_N5111), 
        .IN2(P1_lt_224_n23) );
  NOR2X0 P1_lt_224_U17 ( .QN(P1_lt_224_n19), .IN1(P1_lt_224_n21), 
        .IN2(P1_lt_224_n22) );
  INVX0 P1_lt_224_U16 ( .ZN(P1_lt_224_n18), .INP(P1_N5427) );
  OR2X1 P1_lt_224_U15 ( .IN2(P1_N5112), .IN1(P1_lt_224_n18), .Q(P1_lt_224_n20)
         );
  NAND2X0 P1_lt_224_U14 ( .IN1(P1_lt_224_n19), .IN2(P1_lt_224_n20), 
        .QN(P1_lt_224_n16) );
  NAND2X0 P1_lt_224_U13 ( .IN1(P1_N5112), .IN2(P1_lt_224_n18), 
        .QN(P1_lt_224_n17) );
  NAND2X0 P1_lt_224_U12 ( .IN1(P1_lt_224_n16), .IN2(P1_lt_224_n17), 
        .QN(P1_lt_224_n15) );
  NOR2X0 P1_lt_224_U11 ( .QN(P1_lt_224_n11), .IN1(P1_lt_224_n14), 
        .IN2(P1_lt_224_n15) );
  NOR2X0 P1_lt_224_U10 ( .QN(P1_lt_224_n12), .IN1(P1_N5113), 
        .IN2(P1_lt_224_n13) );
  NOR2X0 P1_lt_224_U9 ( .QN(P1_lt_224_n9), .IN1(P1_lt_224_n11), 
        .IN2(P1_lt_224_n12) );
  INVX0 P1_lt_224_U8 ( .ZN(P1_lt_224_n8), .INP(P1_N5429) );
  OR2X1 P1_lt_224_U7 ( .IN2(P1_N5114), .IN1(P1_lt_224_n8), .Q(P1_lt_224_n10)
         );
  NAND2X0 P1_lt_224_U6 ( .IN1(P1_lt_224_n9), .IN2(P1_lt_224_n10), 
        .QN(P1_lt_224_n6) );
  NAND2X0 P1_lt_224_U5 ( .IN1(P1_N5114), .IN2(P1_lt_224_n8), .QN(P1_lt_224_n7)
         );
  NAND2X0 P1_lt_224_U4 ( .IN1(P1_lt_224_n6), .IN2(P1_lt_224_n7), 
        .QN(P1_lt_224_n3) );
  NAND2X0 P1_lt_224_U3 ( .IN1(P1_N5115), .IN2(P1_lt_224_n5), .QN(P1_lt_224_n4)
         );
  NAND2X0 P1_lt_224_U2 ( .IN1(P1_lt_224_n3), .IN2(P1_lt_224_n4), 
        .QN(P1_lt_224_n2) );
  NAND2X0 P1_lt_224_U1 ( .IN1(P1_lt_224_n1), .IN2(P1_lt_224_n2), .QN(P1_N5362)
         );
  INVX0 P1_lt_224_U157 ( .ZN(P1_lt_224_n5), .INP(P1_N5430) );
  OR2X1 P1_lt_224_U156 ( .IN2(P1_N5115), .IN1(P1_lt_224_n5), .Q(P1_lt_224_n1)
         );
  INVX0 P1_lt_224_U155 ( .ZN(P1_lt_224_n13), .INP(P1_N5428) );
  AND2X1 P1_lt_224_U154 ( .IN1(P1_lt_224_n13), .IN2(P1_N5113), 
        .Q(P1_lt_224_n14) );
  INVX0 P1_lt_224_U153 ( .ZN(P1_lt_224_n23), .INP(P1_N5426) );
  AND2X1 P1_lt_224_U152 ( .IN1(P1_lt_224_n23), .IN2(P1_N5111), 
        .Q(P1_lt_224_n24) );
  INVX0 P1_lt_224_U151 ( .ZN(P1_lt_224_n33), .INP(P1_N5424) );
  AND2X1 P1_lt_224_U150 ( .IN1(P1_lt_224_n33), .IN2(P1_N5109), 
        .Q(P1_lt_224_n34) );
  INVX0 P1_lt_224_U149 ( .ZN(P1_lt_224_n43), .INP(P1_N5422) );
  AND2X1 P1_lt_224_U148 ( .IN1(P1_lt_224_n43), .IN2(P1_N5107), 
        .Q(P1_lt_224_n44) );
  INVX0 P1_lt_224_U147 ( .ZN(P1_lt_224_n53), .INP(P1_N5420) );
  AND2X1 P1_lt_224_U146 ( .IN1(P1_lt_224_n53), .IN2(P1_N5105), 
        .Q(P1_lt_224_n54) );
  INVX0 P1_lt_224_U145 ( .ZN(P1_lt_224_n63), .INP(P1_N5418) );
  AND2X1 P1_lt_224_U144 ( .IN1(P1_lt_224_n63), .IN2(P1_N5103), 
        .Q(P1_lt_224_n64) );
  INVX0 P1_lt_224_U143 ( .ZN(P1_lt_224_n73), .INP(P1_N5416) );
  AND2X1 P1_lt_224_U142 ( .IN1(P1_lt_224_n73), .IN2(P1_N5101), 
        .Q(P1_lt_224_n74) );
  INVX0 P1_lt_224_U141 ( .ZN(P1_lt_224_n83), .INP(P1_N5414) );
  AND2X1 P1_lt_224_U140 ( .IN1(P1_lt_224_n83), .IN2(P1_N5099), 
        .Q(P1_lt_224_n84) );
  INVX0 P1_lt_224_U139 ( .ZN(P1_lt_224_n93), .INP(P1_N5412) );
  AND2X1 P1_lt_224_U138 ( .IN1(P1_lt_224_n93), .IN2(P1_N5097), 
        .Q(P1_lt_224_n94) );
  INVX0 P1_lt_224_U137 ( .ZN(P1_lt_224_n103), .INP(P1_N5410) );
  AND2X1 P1_lt_224_U136 ( .IN1(P1_lt_224_n103), .IN2(P1_N5095), 
        .Q(P1_lt_224_n104) );
  NOR2X0 P1_lt_224_U134 ( .QN(P1_lt_224_n114), .IN1(P1_N5408), .IN2(n7273) );
  INVX0 P1_lt_224_U133 ( .ZN(P1_lt_224_n123), .INP(P1_N5406) );
  AND2X1 P1_lt_224_U132 ( .IN1(P1_lt_224_n123), .IN2(P1_N5091), 
        .Q(P1_lt_224_n124) );
  INVX0 P1_lt_224_U131 ( .ZN(P1_lt_224_n133), .INP(P1_N5404) );
  AND2X1 P1_lt_224_U130 ( .IN1(P1_lt_224_n133), .IN2(P1_N5089), 
        .Q(P1_lt_224_n134) );
  INVX0 P1_lt_224_U129 ( .ZN(P1_lt_224_n143), .INP(P1_N5402) );
  AND2X1 P1_lt_224_U128 ( .IN1(P1_lt_224_n143), .IN2(P1_N5087), 
        .Q(P1_lt_224_n144) );
  INVX0 P1_lt_224_U127 ( .ZN(P1_lt_224_n154), .INP(P1_N5400) );
  INVX0 P1_lt_224_U126 ( .ZN(P1_lt_224_n156), .INP(P1_N5084) );
  NOR2X0 P1_lt_224_U125 ( .QN(P1_lt_224_n153), .IN1(P1_lt_224_n156), 
        .IN2(P1_N5399) );
  AND2X1 P1_lt_224_U124 ( .IN1(P1_lt_224_n154), .IN2(P1_lt_224_n153), 
        .Q(P1_lt_224_n155) );
  NOR2X0 P1_lt_224_U123 ( .QN(P1_lt_224_n151), .IN1(P1_N5085), 
        .IN2(P1_lt_224_n155) );
  NOR2X0 P1_lt_224_U122 ( .QN(P1_lt_224_n152), .IN1(P1_lt_224_n153), 
        .IN2(P1_lt_224_n154) );
  NOR2X0 P1_lt_224_U121 ( .QN(P1_lt_224_n149), .IN1(P1_lt_224_n151), 
        .IN2(P1_lt_224_n152) );
  INVX0 P1_lt_224_U120 ( .ZN(P1_lt_224_n148), .INP(P1_N5401) );
  OR2X1 P1_lt_224_U119 ( .IN2(P1_N5086), .IN1(P1_lt_224_n148), 
        .Q(P1_lt_224_n150) );
  NAND2X0 P1_lt_224_U118 ( .IN1(P1_lt_224_n149), .IN2(P1_lt_224_n150), 
        .QN(P1_lt_224_n146) );
  NAND2X0 P1_lt_224_U117 ( .IN1(P1_N5086), .IN2(P1_lt_224_n148), 
        .QN(P1_lt_224_n147) );
  NAND2X0 P1_lt_224_U116 ( .IN1(P1_lt_224_n146), .IN2(P1_lt_224_n147), 
        .QN(P1_lt_224_n145) );
  NOR2X0 P1_lt_224_U115 ( .QN(P1_lt_224_n141), .IN1(P1_lt_224_n144), 
        .IN2(P1_lt_224_n145) );
  NOR2X0 P1_lt_224_U114 ( .QN(P1_lt_224_n142), .IN1(P1_N5087), 
        .IN2(P1_lt_224_n143) );
  NOR2X0 P1_lt_224_U113 ( .QN(P1_lt_224_n139), .IN1(P1_lt_224_n141), 
        .IN2(P1_lt_224_n142) );
  INVX0 P1_lt_224_U112 ( .ZN(P1_lt_224_n138), .INP(P1_N5403) );
  OR2X1 P1_lt_224_U111 ( .IN2(P1_N5088), .IN1(P1_lt_224_n138), 
        .Q(P1_lt_224_n140) );
  NAND2X0 P1_lt_224_U110 ( .IN1(P1_lt_224_n139), .IN2(P1_lt_224_n140), 
        .QN(P1_lt_224_n136) );
  NAND2X0 P1_lt_224_U109 ( .IN1(P1_N5088), .IN2(P1_lt_224_n138), 
        .QN(P1_lt_224_n137) );
  NAND2X0 P1_lt_224_U108 ( .IN1(P1_lt_224_n136), .IN2(P1_lt_224_n137), 
        .QN(P1_lt_224_n135) );
  NOR2X0 P1_lt_224_U107 ( .QN(P1_lt_224_n131), .IN1(P1_lt_224_n134), 
        .IN2(P1_lt_224_n135) );
  NOR2X0 P1_lt_224_U106 ( .QN(P1_lt_224_n132), .IN1(P1_N5089), 
        .IN2(P1_lt_224_n133) );
  NOR2X0 P1_lt_224_U105 ( .QN(P1_lt_224_n129), .IN1(P1_lt_224_n131), 
        .IN2(P1_lt_224_n132) );
  INVX0 P1_lt_224_U104 ( .ZN(P1_lt_224_n128), .INP(P1_N5405) );
  OR2X1 P1_lt_224_U103 ( .IN2(P1_N5090), .IN1(P1_lt_224_n128), 
        .Q(P1_lt_224_n130) );
  NAND2X0 P1_lt_224_U102 ( .IN1(P1_lt_224_n129), .IN2(P1_lt_224_n130), 
        .QN(P1_lt_224_n126) );
  NAND2X0 P1_lt_224_U101 ( .IN1(P1_N5090), .IN2(P1_lt_224_n128), 
        .QN(P1_lt_224_n127) );
  NAND2X0 P1_lt_224_U100 ( .IN1(P1_lt_224_n126), .IN2(P1_lt_224_n127), 
        .QN(P1_lt_224_n125) );
  NOR2X0 P1_lt_224_U99 ( .QN(P1_lt_224_n121), .IN1(P1_lt_224_n124), 
        .IN2(P1_lt_224_n125) );
  NOR2X0 P1_lt_224_U98 ( .QN(P1_lt_224_n122), .IN1(P1_N5091), 
        .IN2(P1_lt_224_n123) );
  NOR2X0 P1_lt_224_U97 ( .QN(P1_lt_224_n119), .IN1(P1_lt_224_n121), 
        .IN2(P1_lt_224_n122) );
  INVX0 P1_lt_224_U96 ( .ZN(P1_lt_224_n118), .INP(P1_N5407) );
  OR2X1 P1_lt_224_U95 ( .IN2(P1_N5092), .IN1(P1_lt_224_n118), 
        .Q(P1_lt_224_n120) );
  NAND2X0 P1_lt_224_U94 ( .IN1(P1_lt_224_n119), .IN2(P1_lt_224_n120), 
        .QN(P1_lt_224_n116) );
  INVX0 P1_lt_232_U64 ( .ZN(P1_lt_232_n78), .INP(P1_N5415) );
  OR2X1 P1_lt_232_U63 ( .IN2(P1_N5100), .IN1(P1_lt_232_n78), .Q(P1_lt_232_n80)
         );
  NAND2X0 P1_lt_232_U62 ( .IN1(P1_lt_232_n79), .IN2(P1_lt_232_n80), 
        .QN(P1_lt_232_n76) );
  NAND2X0 P1_lt_232_U61 ( .IN1(P1_N5100), .IN2(P1_lt_232_n78), 
        .QN(P1_lt_232_n77) );
  NAND2X0 P1_lt_232_U60 ( .IN1(P1_lt_232_n76), .IN2(P1_lt_232_n77), 
        .QN(P1_lt_232_n75) );
  NOR2X0 P1_lt_232_U59 ( .QN(P1_lt_232_n71), .IN1(P1_lt_232_n74), 
        .IN2(P1_lt_232_n75) );
  NOR2X0 P1_lt_232_U58 ( .QN(P1_lt_232_n72), .IN1(P1_N5101), 
        .IN2(P1_lt_232_n73) );
  NOR2X0 P1_lt_232_U57 ( .QN(P1_lt_232_n69), .IN1(P1_lt_232_n71), 
        .IN2(P1_lt_232_n72) );
  INVX0 P1_lt_232_U56 ( .ZN(P1_lt_232_n68), .INP(P1_N5417) );
  OR2X1 P1_lt_232_U55 ( .IN2(P1_N5102), .IN1(P1_lt_232_n68), .Q(P1_lt_232_n70)
         );
  NAND2X0 P1_lt_232_U54 ( .IN1(P1_lt_232_n69), .IN2(P1_lt_232_n70), 
        .QN(P1_lt_232_n66) );
  NAND2X0 P1_lt_232_U53 ( .IN1(P1_N5102), .IN2(P1_lt_232_n68), 
        .QN(P1_lt_232_n67) );
  NAND2X0 P1_lt_232_U52 ( .IN1(P1_lt_232_n66), .IN2(P1_lt_232_n67), 
        .QN(P1_lt_232_n65) );
  NOR2X0 P1_lt_232_U51 ( .QN(P1_lt_232_n61), .IN1(P1_lt_232_n64), 
        .IN2(P1_lt_232_n65) );
  NOR2X0 P1_lt_232_U50 ( .QN(P1_lt_232_n62), .IN1(P1_N5103), 
        .IN2(P1_lt_232_n63) );
  NOR2X0 P1_lt_232_U49 ( .QN(P1_lt_232_n59), .IN1(P1_lt_232_n61), 
        .IN2(P1_lt_232_n62) );
  INVX0 P1_lt_232_U48 ( .ZN(P1_lt_232_n58), .INP(P1_N5419) );
  OR2X1 P1_lt_232_U47 ( .IN2(P1_N5104), .IN1(P1_lt_232_n58), .Q(P1_lt_232_n60)
         );
  NAND2X0 P1_lt_232_U46 ( .IN1(P1_lt_232_n59), .IN2(P1_lt_232_n60), 
        .QN(P1_lt_232_n56) );
  NAND2X0 P1_lt_232_U45 ( .IN1(P1_N5104), .IN2(P1_lt_232_n58), 
        .QN(P1_lt_232_n57) );
  NAND2X0 P1_lt_232_U44 ( .IN1(P1_lt_232_n56), .IN2(P1_lt_232_n57), 
        .QN(P1_lt_232_n55) );
  NOR2X0 P1_lt_232_U43 ( .QN(P1_lt_232_n51), .IN1(P1_lt_232_n54), 
        .IN2(P1_lt_232_n55) );
  NOR2X0 P1_lt_232_U42 ( .QN(P1_lt_232_n52), .IN1(P1_N5105), 
        .IN2(P1_lt_232_n53) );
  NOR2X0 P1_lt_232_U41 ( .QN(P1_lt_232_n49), .IN1(P1_lt_232_n51), 
        .IN2(P1_lt_232_n52) );
  INVX0 P1_lt_232_U40 ( .ZN(P1_lt_232_n48), .INP(P1_N5421) );
  OR2X1 P1_lt_232_U39 ( .IN2(P1_N5106), .IN1(P1_lt_232_n48), .Q(P1_lt_232_n50)
         );
  NAND2X0 P1_lt_232_U38 ( .IN1(P1_lt_232_n49), .IN2(P1_lt_232_n50), 
        .QN(P1_lt_232_n46) );
  NAND2X0 P1_lt_232_U37 ( .IN1(P1_N5106), .IN2(P1_lt_232_n48), 
        .QN(P1_lt_232_n47) );
  NAND2X0 P1_lt_232_U36 ( .IN1(P1_lt_232_n46), .IN2(P1_lt_232_n47), 
        .QN(P1_lt_232_n45) );
  NOR2X0 P1_lt_232_U35 ( .QN(P1_lt_232_n41), .IN1(P1_lt_232_n44), 
        .IN2(P1_lt_232_n45) );
  NOR2X0 P1_lt_232_U34 ( .QN(P1_lt_232_n42), .IN1(P1_N5107), 
        .IN2(P1_lt_232_n43) );
  NOR2X0 P1_lt_232_U33 ( .QN(P1_lt_232_n39), .IN1(P1_lt_232_n41), 
        .IN2(P1_lt_232_n42) );
  INVX0 P1_lt_232_U32 ( .ZN(P1_lt_232_n38), .INP(P1_N5423) );
  OR2X1 P1_lt_232_U31 ( .IN2(P1_N5108), .IN1(P1_lt_232_n38), .Q(P1_lt_232_n40)
         );
  NAND2X0 P1_lt_232_U30 ( .IN1(P1_lt_232_n39), .IN2(P1_lt_232_n40), 
        .QN(P1_lt_232_n36) );
  NAND2X0 P1_lt_232_U29 ( .IN1(P1_N5108), .IN2(P1_lt_232_n38), 
        .QN(P1_lt_232_n37) );
  NAND2X0 P1_lt_232_U28 ( .IN1(P1_lt_232_n36), .IN2(P1_lt_232_n37), 
        .QN(P1_lt_232_n35) );
  NOR2X0 P1_lt_232_U27 ( .QN(P1_lt_232_n31), .IN1(P1_lt_232_n34), 
        .IN2(P1_lt_232_n35) );
  NOR2X0 P1_lt_232_U26 ( .QN(P1_lt_232_n32), .IN1(P1_N5109), 
        .IN2(P1_lt_232_n33) );
  NOR2X0 P1_lt_232_U25 ( .QN(P1_lt_232_n29), .IN1(P1_lt_232_n31), 
        .IN2(P1_lt_232_n32) );
  INVX0 P1_lt_232_U24 ( .ZN(P1_lt_232_n28), .INP(P1_N5425) );
  OR2X1 P1_lt_232_U23 ( .IN2(P1_N5110), .IN1(P1_lt_232_n28), .Q(P1_lt_232_n30)
         );
  NAND2X0 P1_lt_232_U22 ( .IN1(P1_lt_232_n29), .IN2(P1_lt_232_n30), 
        .QN(P1_lt_232_n26) );
  NAND2X0 P1_lt_232_U21 ( .IN1(P1_N5110), .IN2(P1_lt_232_n28), 
        .QN(P1_lt_232_n27) );
  NAND2X0 P1_lt_232_U20 ( .IN1(P1_lt_232_n26), .IN2(P1_lt_232_n27), 
        .QN(P1_lt_232_n25) );
  NOR2X0 P1_lt_232_U19 ( .QN(P1_lt_232_n21), .IN1(P1_lt_232_n24), 
        .IN2(P1_lt_232_n25) );
  NOR2X0 P1_lt_232_U18 ( .QN(P1_lt_232_n22), .IN1(P1_N5111), 
        .IN2(P1_lt_232_n23) );
  NOR2X0 P1_lt_232_U17 ( .QN(P1_lt_232_n19), .IN1(P1_lt_232_n21), 
        .IN2(P1_lt_232_n22) );
  INVX0 P1_lt_232_U16 ( .ZN(P1_lt_232_n18), .INP(P1_N5427) );
  OR2X1 P1_lt_232_U15 ( .IN2(P1_N5112), .IN1(P1_lt_232_n18), .Q(P1_lt_232_n20)
         );
  NAND2X0 P1_lt_232_U14 ( .IN1(P1_lt_232_n19), .IN2(P1_lt_232_n20), 
        .QN(P1_lt_232_n16) );
  NAND2X0 P1_lt_232_U13 ( .IN1(P1_N5112), .IN2(P1_lt_232_n18), 
        .QN(P1_lt_232_n17) );
  NAND2X0 P1_lt_232_U12 ( .IN1(P1_lt_232_n16), .IN2(P1_lt_232_n17), 
        .QN(P1_lt_232_n15) );
  NOR2X0 P1_lt_232_U11 ( .QN(P1_lt_232_n11), .IN1(P1_lt_232_n14), 
        .IN2(P1_lt_232_n15) );
  NOR2X0 P1_lt_232_U10 ( .QN(P1_lt_232_n12), .IN1(P1_N5113), 
        .IN2(P1_lt_232_n13) );
  NOR2X0 P1_lt_232_U9 ( .QN(P1_lt_232_n9), .IN1(P1_lt_232_n11), 
        .IN2(P1_lt_232_n12) );
  INVX0 P1_lt_232_U8 ( .ZN(P1_lt_232_n8), .INP(P1_N5429) );
  OR2X1 P1_lt_232_U7 ( .IN2(P1_N5114), .IN1(P1_lt_232_n8), .Q(P1_lt_232_n10)
         );
  NAND2X0 P1_lt_232_U6 ( .IN1(P1_lt_232_n9), .IN2(P1_lt_232_n10), 
        .QN(P1_lt_232_n6) );
  NAND2X0 P1_lt_232_U5 ( .IN1(P1_N5114), .IN2(P1_lt_232_n8), .QN(P1_lt_232_n7)
         );
  NAND2X0 P1_lt_232_U4 ( .IN1(P1_lt_232_n6), .IN2(P1_lt_232_n7), 
        .QN(P1_lt_232_n3) );
  NAND2X0 P1_lt_232_U3 ( .IN1(P1_N5115), .IN2(P1_lt_232_n5), .QN(P1_lt_232_n4)
         );
  NAND2X0 P1_lt_232_U2 ( .IN1(P1_lt_232_n3), .IN2(P1_lt_232_n4), 
        .QN(P1_lt_232_n2) );
  NAND2X0 P1_lt_232_U1 ( .IN1(P1_lt_232_n1), .IN2(P1_lt_232_n2), .QN(P1_N5431)
         );
  INVX0 P1_lt_232_U157 ( .ZN(P1_lt_232_n5), .INP(P1_N5430) );
  OR2X1 P1_lt_232_U156 ( .IN2(P1_N5115), .IN1(P1_lt_232_n5), .Q(P1_lt_232_n1)
         );
  INVX0 P1_lt_232_U155 ( .ZN(P1_lt_232_n13), .INP(P1_N5428) );
  AND2X1 P1_lt_232_U154 ( .IN1(P1_lt_232_n13), .IN2(P1_N5113), 
        .Q(P1_lt_232_n14) );
  INVX0 P1_lt_232_U153 ( .ZN(P1_lt_232_n23), .INP(P1_N5426) );
  AND2X1 P1_lt_232_U152 ( .IN1(P1_lt_232_n23), .IN2(P1_N5111), 
        .Q(P1_lt_232_n24) );
  INVX0 P1_lt_232_U151 ( .ZN(P1_lt_232_n33), .INP(P1_N5424) );
  AND2X1 P1_lt_232_U150 ( .IN1(P1_lt_232_n33), .IN2(P1_N5109), 
        .Q(P1_lt_232_n34) );
  INVX0 P1_lt_232_U149 ( .ZN(P1_lt_232_n43), .INP(P1_N5422) );
  AND2X1 P1_lt_232_U148 ( .IN1(P1_lt_232_n43), .IN2(P1_N5107), 
        .Q(P1_lt_232_n44) );
  INVX0 P1_lt_232_U147 ( .ZN(P1_lt_232_n53), .INP(P1_N5420) );
  AND2X1 P1_lt_232_U146 ( .IN1(P1_lt_232_n53), .IN2(P1_N5105), 
        .Q(P1_lt_232_n54) );
  INVX0 P1_lt_232_U145 ( .ZN(P1_lt_232_n63), .INP(P1_N5418) );
  AND2X1 P1_lt_232_U144 ( .IN1(P1_lt_232_n63), .IN2(P1_N5103), 
        .Q(P1_lt_232_n64) );
  INVX0 P1_lt_232_U143 ( .ZN(P1_lt_232_n73), .INP(P1_N5416) );
  AND2X1 P1_lt_232_U142 ( .IN1(P1_lt_232_n73), .IN2(P1_N5101), 
        .Q(P1_lt_232_n74) );
  INVX0 P1_lt_232_U141 ( .ZN(P1_lt_232_n83), .INP(P1_N5414) );
  AND2X1 P1_lt_232_U140 ( .IN1(P1_lt_232_n83), .IN2(P1_N5099), 
        .Q(P1_lt_232_n84) );
  INVX0 P1_lt_232_U139 ( .ZN(P1_lt_232_n93), .INP(P1_N5412) );
  AND2X1 P1_lt_232_U138 ( .IN1(P1_lt_232_n93), .IN2(P1_N5097), 
        .Q(P1_lt_232_n94) );
  INVX0 P1_lt_232_U137 ( .ZN(P1_lt_232_n103), .INP(P1_N5410) );
  AND2X1 P1_lt_232_U136 ( .IN1(P1_lt_232_n103), .IN2(P1_N5095), 
        .Q(P1_lt_232_n104) );
  NOR2X0 P1_lt_232_U134 ( .QN(P1_lt_232_n114), .IN1(P1_N5408), .IN2(n7273) );
  INVX0 P1_lt_232_U133 ( .ZN(P1_lt_232_n123), .INP(P1_N5406) );
  AND2X1 P1_lt_232_U132 ( .IN1(P1_lt_232_n123), .IN2(P1_N5091), 
        .Q(P1_lt_232_n124) );
  INVX0 P1_lt_232_U131 ( .ZN(P1_lt_232_n133), .INP(P1_N5404) );
  AND2X1 P1_lt_232_U130 ( .IN1(P1_lt_232_n133), .IN2(P1_N5089), 
        .Q(P1_lt_232_n134) );
  INVX0 P1_lt_232_U129 ( .ZN(P1_lt_232_n143), .INP(P1_N5402) );
  AND2X1 P1_lt_232_U128 ( .IN1(P1_lt_232_n143), .IN2(P1_N5087), 
        .Q(P1_lt_232_n144) );
  INVX0 P1_lt_232_U127 ( .ZN(P1_lt_232_n154), .INP(P1_N5400) );
  INVX0 P1_lt_232_U126 ( .ZN(P1_lt_232_n156), .INP(P1_N5084) );
  NOR2X0 P1_lt_232_U125 ( .QN(P1_lt_232_n153), .IN1(P1_lt_232_n156), 
        .IN2(P1_N5399) );
  AND2X1 P1_lt_232_U124 ( .IN1(P1_lt_232_n154), .IN2(P1_lt_232_n153), 
        .Q(P1_lt_232_n155) );
  NOR2X0 P1_lt_232_U123 ( .QN(P1_lt_232_n151), .IN1(P1_N5085), 
        .IN2(P1_lt_232_n155) );
  NOR2X0 P1_lt_232_U122 ( .QN(P1_lt_232_n152), .IN1(P1_lt_232_n153), 
        .IN2(P1_lt_232_n154) );
  NOR2X0 P1_lt_232_U121 ( .QN(P1_lt_232_n149), .IN1(P1_lt_232_n151), 
        .IN2(P1_lt_232_n152) );
  INVX0 P1_lt_232_U120 ( .ZN(P1_lt_232_n148), .INP(P1_N5401) );
  OR2X1 P1_lt_232_U119 ( .IN2(P1_N5086), .IN1(P1_lt_232_n148), 
        .Q(P1_lt_232_n150) );
  NAND2X0 P1_lt_232_U118 ( .IN1(P1_lt_232_n149), .IN2(P1_lt_232_n150), 
        .QN(P1_lt_232_n146) );
  NAND2X0 P1_lt_232_U117 ( .IN1(P1_N5086), .IN2(P1_lt_232_n148), 
        .QN(P1_lt_232_n147) );
  NAND2X0 P1_lt_232_U116 ( .IN1(P1_lt_232_n146), .IN2(P1_lt_232_n147), 
        .QN(P1_lt_232_n145) );
  NOR2X0 P1_lt_232_U115 ( .QN(P1_lt_232_n141), .IN1(P1_lt_232_n144), 
        .IN2(P1_lt_232_n145) );
  NOR2X0 P1_lt_232_U114 ( .QN(P1_lt_232_n142), .IN1(P1_N5087), 
        .IN2(P1_lt_232_n143) );
  NOR2X0 P1_lt_232_U113 ( .QN(P1_lt_232_n139), .IN1(P1_lt_232_n141), 
        .IN2(P1_lt_232_n142) );
  INVX0 P1_lt_232_U112 ( .ZN(P1_lt_232_n138), .INP(P1_N5403) );
  OR2X1 P1_lt_232_U111 ( .IN2(P1_N5088), .IN1(P1_lt_232_n138), 
        .Q(P1_lt_232_n140) );
  NAND2X0 P1_lt_232_U110 ( .IN1(P1_lt_232_n139), .IN2(P1_lt_232_n140), 
        .QN(P1_lt_232_n136) );
  NAND2X0 P1_lt_232_U109 ( .IN1(P1_N5088), .IN2(P1_lt_232_n138), 
        .QN(P1_lt_232_n137) );
  NAND2X0 P1_lt_232_U108 ( .IN1(P1_lt_232_n136), .IN2(P1_lt_232_n137), 
        .QN(P1_lt_232_n135) );
  NOR2X0 P1_lt_232_U107 ( .QN(P1_lt_232_n131), .IN1(P1_lt_232_n134), 
        .IN2(P1_lt_232_n135) );
  NOR2X0 P1_lt_232_U106 ( .QN(P1_lt_232_n132), .IN1(P1_N5089), 
        .IN2(P1_lt_232_n133) );
  NOR2X0 P1_lt_232_U105 ( .QN(P1_lt_232_n129), .IN1(P1_lt_232_n131), 
        .IN2(P1_lt_232_n132) );
  INVX0 P1_lt_232_U104 ( .ZN(P1_lt_232_n128), .INP(P1_N5405) );
  OR2X1 P1_lt_232_U103 ( .IN2(P1_N5090), .IN1(P1_lt_232_n128), 
        .Q(P1_lt_232_n130) );
  NAND2X0 P1_lt_232_U102 ( .IN1(P1_lt_232_n129), .IN2(P1_lt_232_n130), 
        .QN(P1_lt_232_n126) );
  NAND2X0 P1_lt_232_U101 ( .IN1(P1_N5090), .IN2(P1_lt_232_n128), 
        .QN(P1_lt_232_n127) );
  NAND2X0 P1_lt_232_U100 ( .IN1(P1_lt_232_n126), .IN2(P1_lt_232_n127), 
        .QN(P1_lt_232_n125) );
  NOR2X0 P1_lt_232_U99 ( .QN(P1_lt_232_n121), .IN1(P1_lt_232_n124), 
        .IN2(P1_lt_232_n125) );
  NOR2X0 P1_lt_232_U98 ( .QN(P1_lt_232_n122), .IN1(P1_N5091), 
        .IN2(P1_lt_232_n123) );
  NOR2X0 P1_lt_232_U97 ( .QN(P1_lt_232_n119), .IN1(P1_lt_232_n121), 
        .IN2(P1_lt_232_n122) );
  INVX0 P1_lt_232_U96 ( .ZN(P1_lt_232_n118), .INP(P1_N5407) );
  OR2X1 P1_lt_232_U95 ( .IN2(P1_N5092), .IN1(P1_lt_232_n118), 
        .Q(P1_lt_232_n120) );
  NAND2X0 P1_lt_232_U94 ( .IN1(P1_lt_232_n119), .IN2(P1_lt_232_n120), 
        .QN(P1_lt_232_n116) );
  NAND2X0 P1_lt_232_U93 ( .IN1(P1_N5092), .IN2(P1_lt_232_n118), 
        .QN(P1_lt_232_n117) );
  NAND2X0 P1_lt_232_U92 ( .IN1(P1_lt_232_n116), .IN2(P1_lt_232_n117), 
        .QN(P1_lt_232_n115) );
  NOR2X0 P1_lt_232_U91 ( .QN(P1_lt_232_n112), .IN1(P1_lt_232_n114), 
        .IN2(P1_lt_232_n115) );
  INVX0 P1_lt_232_U90 ( .ZN(P1_lt_232_n108), .INP(P1_N5409) );
  NOR2X0 P1_lt_232_U89 ( .QN(P1_lt_232_n113), .IN1(P1_N5094), 
        .IN2(P1_lt_232_n108) );
  NOR2X0 P1_lt_232_U88 ( .QN(P1_lt_232_n109), .IN1(P1_lt_232_n112), 
        .IN2(P1_lt_232_n113) );
  NAND2X0 P1_lt_232_U87 ( .IN1(P1_N5408), .IN2(n7273), .QN(P1_lt_232_n110) );
  NAND2X0 P1_lt_232_U86 ( .IN1(P1_lt_232_n109), .IN2(P1_lt_232_n110), 
        .QN(P1_lt_232_n106) );
  NAND2X0 P1_lt_232_U85 ( .IN1(P1_N5094), .IN2(P1_lt_232_n108), 
        .QN(P1_lt_232_n107) );
  NAND2X0 P1_lt_232_U84 ( .IN1(P1_lt_232_n106), .IN2(P1_lt_232_n107), 
        .QN(P1_lt_232_n105) );
  NOR2X0 P1_lt_232_U83 ( .QN(P1_lt_232_n101), .IN1(P1_lt_232_n104), 
        .IN2(P1_lt_232_n105) );
  NOR2X0 P1_lt_232_U82 ( .QN(P1_lt_232_n102), .IN1(P1_N5095), 
        .IN2(P1_lt_232_n103) );
  NOR2X0 P1_lt_232_U81 ( .QN(P1_lt_232_n99), .IN1(P1_lt_232_n101), 
        .IN2(P1_lt_232_n102) );
  INVX0 P1_lt_232_U80 ( .ZN(P1_lt_232_n98), .INP(P1_N5411) );
  OR2X1 P1_lt_232_U79 ( .IN2(P1_N5096), .IN1(P1_lt_232_n98), 
        .Q(P1_lt_232_n100) );
  NAND2X0 P1_lt_232_U78 ( .IN1(P1_lt_232_n99), .IN2(P1_lt_232_n100), 
        .QN(P1_lt_232_n96) );
  NAND2X0 P1_lt_232_U77 ( .IN1(P1_N5096), .IN2(P1_lt_232_n98), 
        .QN(P1_lt_232_n97) );
  NAND2X0 P1_lt_232_U76 ( .IN1(P1_lt_232_n96), .IN2(P1_lt_232_n97), 
        .QN(P1_lt_232_n95) );
  NOR2X0 P1_lt_232_U75 ( .QN(P1_lt_232_n91), .IN1(P1_lt_232_n94), 
        .IN2(P1_lt_232_n95) );
  NOR2X0 P1_lt_232_U74 ( .QN(P1_lt_232_n92), .IN1(P1_N5097), 
        .IN2(P1_lt_232_n93) );
  NOR2X0 P1_lt_232_U73 ( .QN(P1_lt_232_n89), .IN1(P1_lt_232_n91), 
        .IN2(P1_lt_232_n92) );
  INVX0 P1_lt_232_U72 ( .ZN(P1_lt_232_n88), .INP(P1_N5413) );
  OR2X1 P1_lt_232_U71 ( .IN2(P1_N5098), .IN1(P1_lt_232_n88), .Q(P1_lt_232_n90)
         );
  NAND2X0 P1_lt_232_U70 ( .IN1(P1_lt_232_n89), .IN2(P1_lt_232_n90), 
        .QN(P1_lt_232_n86) );
  NAND2X0 P1_lt_232_U69 ( .IN1(P1_N5098), .IN2(P1_lt_232_n88), 
        .QN(P1_lt_232_n87) );
  NAND2X0 P1_lt_232_U68 ( .IN1(P1_lt_232_n86), .IN2(P1_lt_232_n87), 
        .QN(P1_lt_232_n85) );
  NOR2X0 P1_lt_232_U67 ( .QN(P1_lt_232_n81), .IN1(P1_lt_232_n84), 
        .IN2(P1_lt_232_n85) );
  NOR2X0 P1_lt_232_U66 ( .QN(P1_lt_232_n82), .IN1(P1_N5099), 
        .IN2(P1_lt_232_n83) );
  NOR2X0 P1_lt_232_U65 ( .QN(P1_lt_232_n79), .IN1(P1_lt_232_n81), 
        .IN2(P1_lt_232_n82) );
  OR2X1 P2_sub_858_U2 ( .IN2(P2_sub_858_n4), .IN1(P2_sub_858_n3), 
        .Q(P2_sub_858_n2) );
  NAND2X0 P2_sub_858_U1 ( .IN1(P2_sub_858_n1), .IN2(P2_sub_858_n2), 
        .QN(P2_N1737) );
  NAND2X0 P2_sub_858_U95 ( .IN1(P2_sub_858_n101), .IN2(P2_sub_858_n96), 
        .QN(P2_sub_858_n99) );
  OR2X1 P2_sub_858_U94 ( .IN2(P2_sub_858_n96), .IN1(P2_sub_858_n101), 
        .Q(P2_sub_858_n100) );
  NAND2X0 P2_sub_858_U93 ( .IN1(P2_sub_858_n99), .IN2(P2_sub_858_n100), 
        .QN(P2_N1752) );
  INVX0 P2_sub_858_U92 ( .ZN(P2_sub_858_n85), .INP(P2_N1511) );
  NAND2X0 P2_sub_858_U91 ( .IN1(n7237), .IN2(P2_sub_858_n85), 
        .QN(P2_sub_858_n97) );
  OR2X1 P2_sub_858_U90 ( .IN2(n7237), .IN1(P2_sub_858_n85), .Q(P2_sub_858_n98)
         );
  NAND2X0 P2_sub_858_U89 ( .IN1(P2_sub_858_n97), .IN2(P2_sub_858_n98), 
        .QN(P2_sub_858_n91) );
  NAND2X0 P2_sub_858_U88 ( .IN1(P2_N5095), .IN2(P2_sub_858_n96), 
        .QN(P2_sub_858_n92) );
  OR2X1 P2_sub_858_U87 ( .IN2(P2_N5095), .IN1(P2_sub_858_n96), 
        .Q(P2_sub_858_n94) );
  NAND2X0 P2_sub_858_U86 ( .IN1(P2_sub_858_n94), .IN2(P2_sub_858_n95), 
        .QN(P2_sub_858_n93) );
  NAND2X0 P2_sub_858_U85 ( .IN1(P2_sub_858_n92), .IN2(P2_sub_858_n93), 
        .QN(P2_sub_858_n86) );
  NAND2X0 P2_sub_858_U84 ( .IN1(P2_sub_858_n91), .IN2(P2_sub_858_n86), 
        .QN(P2_sub_858_n89) );
  OR2X1 P2_sub_858_U83 ( .IN2(P2_sub_858_n86), .IN1(P2_sub_858_n91), 
        .Q(P2_sub_858_n90) );
  NAND2X0 P2_sub_858_U82 ( .IN1(P2_sub_858_n89), .IN2(P2_sub_858_n90), 
        .QN(P2_N1753) );
  INVX0 P2_sub_858_U81 ( .ZN(P2_sub_858_n75), .INP(P2_N1512) );
  NAND2X0 P2_sub_858_U80 ( .IN1(n7231), .IN2(P2_sub_858_n75), 
        .QN(P2_sub_858_n87) );
  OR2X1 P2_sub_858_U79 ( .IN2(n7231), .IN1(P2_sub_858_n75), .Q(P2_sub_858_n88)
         );
  NAND2X0 P2_sub_858_U78 ( .IN1(P2_sub_858_n87), .IN2(P2_sub_858_n88), 
        .QN(P2_sub_858_n81) );
  NAND2X0 P2_sub_858_U77 ( .IN1(n7237), .IN2(P2_sub_858_n86), 
        .QN(P2_sub_858_n82) );
  OR2X1 P2_sub_858_U76 ( .IN2(n7237), .IN1(P2_sub_858_n86), .Q(P2_sub_858_n84)
         );
  NAND2X0 P2_sub_858_U75 ( .IN1(P2_sub_858_n84), .IN2(P2_sub_858_n85), 
        .QN(P2_sub_858_n83) );
  NAND2X0 P2_sub_858_U74 ( .IN1(P2_sub_858_n82), .IN2(P2_sub_858_n83), 
        .QN(P2_sub_858_n76) );
  NAND2X0 P2_sub_858_U73 ( .IN1(P2_sub_858_n81), .IN2(P2_sub_858_n76), 
        .QN(P2_sub_858_n79) );
  OR2X1 P2_sub_858_U72 ( .IN2(P2_sub_858_n76), .IN1(P2_sub_858_n81), 
        .Q(P2_sub_858_n80) );
  NAND2X0 P2_sub_858_U71 ( .IN1(P2_sub_858_n79), .IN2(P2_sub_858_n80), 
        .QN(P2_N1754) );
  INVX0 P2_sub_858_U70 ( .ZN(P2_sub_858_n64), .INP(P2_N1513) );
  NAND2X0 P2_sub_858_U69 ( .IN1(P2_N5098), .IN2(P2_sub_858_n64), 
        .QN(P2_sub_858_n77) );
  OR2X1 P2_sub_858_U68 ( .IN2(P2_N5098), .IN1(P2_sub_858_n64), 
        .Q(P2_sub_858_n78) );
  NAND2X0 P2_sub_858_U67 ( .IN1(P2_sub_858_n77), .IN2(P2_sub_858_n78), 
        .QN(P2_sub_858_n71) );
  NAND2X0 P2_sub_858_U66 ( .IN1(n7231), .IN2(P2_sub_858_n76), 
        .QN(P2_sub_858_n72) );
  OR2X1 P2_sub_858_U65 ( .IN2(n7231), .IN1(P2_sub_858_n76), .Q(P2_sub_858_n74)
         );
  NAND2X0 P2_sub_858_U64 ( .IN1(P2_sub_858_n74), .IN2(P2_sub_858_n75), 
        .QN(P2_sub_858_n73) );
  NAND2X0 P2_sub_858_U63 ( .IN1(P2_sub_858_n72), .IN2(P2_sub_858_n73), 
        .QN(P2_sub_858_n65) );
  NAND2X0 P2_sub_858_U62 ( .IN1(P2_sub_858_n71), .IN2(P2_sub_858_n65), 
        .QN(P2_sub_858_n69) );
  OR2X1 P2_sub_858_U61 ( .IN2(P2_sub_858_n65), .IN1(P2_sub_858_n71), 
        .Q(P2_sub_858_n70) );
  NAND2X0 P2_sub_858_U60 ( .IN1(P2_sub_858_n69), .IN2(P2_sub_858_n70), 
        .QN(P2_N1755) );
  OR2X1 P2_sub_858_U58 ( .IN2(P2_N1514), .IN1(n7222), .Q(P2_sub_858_n66) );
  NAND2X0 P2_sub_858_U57 ( .IN1(P2_N1514), .IN2(n7222), .QN(P2_sub_858_n67) );
  NAND2X0 P2_sub_858_U56 ( .IN1(P2_sub_858_n66), .IN2(P2_sub_858_n67), 
        .QN(P2_sub_858_n60) );
  NAND2X0 P2_sub_858_U55 ( .IN1(P2_N5098), .IN2(P2_sub_858_n65), 
        .QN(P2_sub_858_n61) );
  OR2X1 P2_sub_858_U54 ( .IN2(P2_N5098), .IN1(P2_sub_858_n65), 
        .Q(P2_sub_858_n63) );
  NAND2X0 P2_sub_858_U53 ( .IN1(P2_sub_858_n63), .IN2(P2_sub_858_n64), 
        .QN(P2_sub_858_n62) );
  NAND2X0 P2_sub_858_U52 ( .IN1(P2_sub_858_n61), .IN2(P2_sub_858_n62), 
        .QN(P2_sub_858_n59) );
  NAND2X0 P2_sub_858_U51 ( .IN1(P2_sub_858_n60), .IN2(P2_sub_858_n59), 
        .QN(P2_sub_858_n57) );
  OR2X1 P2_sub_858_U50 ( .IN2(P2_sub_858_n60), .IN1(P2_sub_858_n59), 
        .Q(P2_sub_858_n58) );
  NAND2X0 P2_sub_858_U49 ( .IN1(P2_sub_858_n57), .IN2(P2_sub_858_n58), 
        .QN(P2_N1756) );
  NAND2X0 P2_sub_858_U48 ( .IN1(P2_N5073), .IN2(P2_sub_858_n56), 
        .QN(P2_sub_858_n54) );
  OR2X1 P2_sub_858_U47 ( .IN2(P2_N5073), .IN1(P2_sub_858_n56), 
        .Q(P2_sub_858_n55) );
  NAND2X0 P2_sub_858_U46 ( .IN1(P2_sub_858_n54), .IN2(P2_sub_858_n55), 
        .QN(P2_sub_858_n52) );
  NAND2X0 P2_sub_858_U45 ( .IN1(P2_sub_858_n52), .IN2(P2_sub_858_n53), 
        .QN(P2_sub_858_n50) );
  OR2X1 P2_sub_858_U44 ( .IN2(P2_sub_858_n53), .IN1(P2_sub_858_n52), 
        .Q(P2_sub_858_n51) );
  NAND2X0 P2_sub_858_U43 ( .IN1(P2_sub_858_n50), .IN2(P2_sub_858_n51), 
        .QN(P2_N1730) );
  NAND2X0 P2_sub_858_U42 ( .IN1(P2_N5074), .IN2(P2_sub_858_n49), 
        .QN(P2_sub_858_n47) );
  OR2X1 P2_sub_858_U41 ( .IN2(P2_N5074), .IN1(P2_sub_858_n49), 
        .Q(P2_sub_858_n48) );
  NAND2X0 P2_sub_858_U40 ( .IN1(P2_sub_858_n47), .IN2(P2_sub_858_n48), 
        .QN(P2_sub_858_n45) );
  NAND2X0 P2_sub_858_U39 ( .IN1(P2_sub_858_n45), .IN2(P2_sub_858_n46), 
        .QN(P2_sub_858_n43) );
  OR2X1 P2_sub_858_U38 ( .IN2(P2_sub_858_n46), .IN1(P2_sub_858_n45), 
        .Q(P2_sub_858_n44) );
  NAND2X0 P2_sub_858_U37 ( .IN1(P2_sub_858_n43), .IN2(P2_sub_858_n44), 
        .QN(P2_N1731) );
  NAND2X0 P2_sub_858_U36 ( .IN1(P2_N5075), .IN2(P2_sub_858_n42), 
        .QN(P2_sub_858_n40) );
  OR2X1 P2_sub_858_U35 ( .IN2(P2_N5075), .IN1(P2_sub_858_n42), 
        .Q(P2_sub_858_n41) );
  NAND2X0 P2_sub_858_U34 ( .IN1(P2_sub_858_n40), .IN2(P2_sub_858_n41), 
        .QN(P2_sub_858_n38) );
  NAND2X0 P2_sub_858_U33 ( .IN1(P2_sub_858_n38), .IN2(P2_sub_858_n39), 
        .QN(P2_sub_858_n36) );
  OR2X1 P2_sub_858_U32 ( .IN2(P2_sub_858_n39), .IN1(P2_sub_858_n38), 
        .Q(P2_sub_858_n37) );
  NAND2X0 P2_sub_858_U31 ( .IN1(P2_sub_858_n36), .IN2(P2_sub_858_n37), 
        .QN(P2_N1732) );
  NAND2X0 P2_sub_858_U30 ( .IN1(n7165), .IN2(P2_sub_858_n35), 
        .QN(P2_sub_858_n33) );
  OR2X1 P2_sub_858_U29 ( .IN2(n7165), .IN1(P2_sub_858_n35), .Q(P2_sub_858_n34)
         );
  NAND2X0 P2_sub_858_U28 ( .IN1(P2_sub_858_n33), .IN2(P2_sub_858_n34), 
        .QN(P2_sub_858_n31) );
  NAND2X0 P2_sub_858_U27 ( .IN1(P2_sub_858_n31), .IN2(P2_sub_858_n32), 
        .QN(P2_sub_858_n29) );
  OR2X1 P2_sub_858_U26 ( .IN2(P2_sub_858_n32), .IN1(P2_sub_858_n31), 
        .Q(P2_sub_858_n30) );
  NAND2X0 P2_sub_858_U25 ( .IN1(P2_sub_858_n29), .IN2(P2_sub_858_n30), 
        .QN(P2_N1733) );
  NAND2X0 P2_sub_858_U24 ( .IN1(P2_N5077), .IN2(P2_sub_858_n28), 
        .QN(P2_sub_858_n26) );
  OR2X1 P2_sub_858_U23 ( .IN2(P2_N5077), .IN1(P2_sub_858_n28), 
        .Q(P2_sub_858_n27) );
  NAND2X0 P2_sub_858_U22 ( .IN1(P2_sub_858_n26), .IN2(P2_sub_858_n27), 
        .QN(P2_sub_858_n24) );
  NAND2X0 P2_sub_858_U21 ( .IN1(P2_sub_858_n24), .IN2(P2_sub_858_n25), 
        .QN(P2_sub_858_n22) );
  OR2X1 P2_sub_858_U20 ( .IN2(P2_sub_858_n25), .IN1(P2_sub_858_n24), 
        .Q(P2_sub_858_n23) );
  NAND2X0 P2_sub_858_U19 ( .IN1(P2_sub_858_n22), .IN2(P2_sub_858_n23), 
        .QN(P2_N1734) );
  NAND2X0 P2_sub_858_U18 ( .IN1(n7158), .IN2(P2_sub_858_n21), 
        .QN(P2_sub_858_n19) );
  OR2X1 P2_sub_858_U17 ( .IN2(n7158), .IN1(P2_sub_858_n21), .Q(P2_sub_858_n20)
         );
  NAND2X0 P2_sub_858_U16 ( .IN1(P2_sub_858_n19), .IN2(P2_sub_858_n20), 
        .QN(P2_sub_858_n17) );
  NAND2X0 P2_sub_858_U15 ( .IN1(P2_sub_858_n17), .IN2(P2_sub_858_n18), 
        .QN(P2_sub_858_n15) );
  OR2X1 P2_sub_858_U14 ( .IN2(P2_sub_858_n18), .IN1(P2_sub_858_n17), 
        .Q(P2_sub_858_n16) );
  NAND2X0 P2_sub_858_U13 ( .IN1(P2_sub_858_n15), .IN2(P2_sub_858_n16), 
        .QN(P2_N1735) );
  NAND2X0 P2_sub_858_U12 ( .IN1(n7154), .IN2(P2_sub_858_n14), 
        .QN(P2_sub_858_n12) );
  OR2X1 P2_sub_858_U11 ( .IN2(n7154), .IN1(P2_sub_858_n14), .Q(P2_sub_858_n13)
         );
  NAND2X0 P2_sub_858_U10 ( .IN1(P2_sub_858_n12), .IN2(P2_sub_858_n13), 
        .QN(P2_sub_858_n10) );
  NAND2X0 P2_sub_858_U9 ( .IN1(P2_sub_858_n10), .IN2(P2_sub_858_n11), 
        .QN(P2_sub_858_n8) );
  OR2X1 P2_sub_858_U8 ( .IN2(P2_sub_858_n11), .IN1(P2_sub_858_n10), 
        .Q(P2_sub_858_n9) );
  NAND2X0 P2_sub_858_U7 ( .IN1(P2_sub_858_n8), .IN2(P2_sub_858_n9), 
        .QN(P2_N1736) );
  NAND2X0 P2_sub_858_U6 ( .IN1(n7151), .IN2(P2_sub_858_n7), .QN(P2_sub_858_n5)
         );
  OR2X1 P2_sub_858_U5 ( .IN2(n7151), .IN1(P2_sub_858_n7), .Q(P2_sub_858_n6) );
  NAND2X0 P2_sub_858_U4 ( .IN1(P2_sub_858_n5), .IN2(P2_sub_858_n6), 
        .QN(P2_sub_858_n3) );
  NAND2X0 P2_sub_858_U3 ( .IN1(P2_sub_858_n3), .IN2(P2_sub_858_n4), 
        .QN(P2_sub_858_n1) );
  OR2X1 P2_sub_858_U188 ( .IN2(P2_sub_858_n184), .IN1(P2_sub_858_n189), 
        .Q(P2_sub_858_n188) );
  NAND2X0 P2_sub_858_U187 ( .IN1(P2_sub_858_n187), .IN2(P2_sub_858_n188), 
        .QN(P2_N1744) );
  INVX0 P2_sub_858_U186 ( .ZN(P2_sub_858_n173), .INP(P2_N1503) );
  NAND2X0 P2_sub_858_U185 ( .IN1(n7194), .IN2(P2_sub_858_n173), 
        .QN(P2_sub_858_n185) );
  OR2X1 P2_sub_858_U184 ( .IN2(n7194), .IN1(P2_sub_858_n173), 
        .Q(P2_sub_858_n186) );
  NAND2X0 P2_sub_858_U183 ( .IN1(P2_sub_858_n185), .IN2(P2_sub_858_n186), 
        .QN(P2_sub_858_n179) );
  NAND2X0 P2_sub_858_U182 ( .IN1(P2_N5087), .IN2(P2_sub_858_n184), 
        .QN(P2_sub_858_n180) );
  OR2X1 P2_sub_858_U181 ( .IN2(P2_N5087), .IN1(P2_sub_858_n184), 
        .Q(P2_sub_858_n182) );
  NAND2X0 P2_sub_858_U180 ( .IN1(P2_sub_858_n182), .IN2(P2_sub_858_n183), 
        .QN(P2_sub_858_n181) );
  NAND2X0 P2_sub_858_U179 ( .IN1(P2_sub_858_n180), .IN2(P2_sub_858_n181), 
        .QN(P2_sub_858_n174) );
  NAND2X0 P2_sub_858_U178 ( .IN1(P2_sub_858_n179), .IN2(P2_sub_858_n174), 
        .QN(P2_sub_858_n177) );
  OR2X1 P2_sub_858_U177 ( .IN2(P2_sub_858_n174), .IN1(P2_sub_858_n179), 
        .Q(P2_sub_858_n178) );
  NAND2X0 P2_sub_858_U176 ( .IN1(P2_sub_858_n177), .IN2(P2_sub_858_n178), 
        .QN(P2_N1745) );
  INVX0 P2_sub_858_U175 ( .ZN(P2_sub_858_n163), .INP(P2_N1504) );
  NAND2X0 P2_sub_858_U174 ( .IN1(n7187), .IN2(P2_sub_858_n163), 
        .QN(P2_sub_858_n175) );
  OR2X1 P2_sub_858_U173 ( .IN2(n7187), .IN1(P2_sub_858_n163), 
        .Q(P2_sub_858_n176) );
  NAND2X0 P2_sub_858_U172 ( .IN1(P2_sub_858_n175), .IN2(P2_sub_858_n176), 
        .QN(P2_sub_858_n169) );
  NAND2X0 P2_sub_858_U171 ( .IN1(n7194), .IN2(P2_sub_858_n174), 
        .QN(P2_sub_858_n170) );
  OR2X1 P2_sub_858_U170 ( .IN2(n7194), .IN1(P2_sub_858_n174), 
        .Q(P2_sub_858_n172) );
  NAND2X0 P2_sub_858_U169 ( .IN1(P2_sub_858_n172), .IN2(P2_sub_858_n173), 
        .QN(P2_sub_858_n171) );
  NAND2X0 P2_sub_858_U168 ( .IN1(P2_sub_858_n170), .IN2(P2_sub_858_n171), 
        .QN(P2_sub_858_n164) );
  NAND2X0 P2_sub_858_U167 ( .IN1(P2_sub_858_n169), .IN2(P2_sub_858_n164), 
        .QN(P2_sub_858_n167) );
  OR2X1 P2_sub_858_U166 ( .IN2(P2_sub_858_n164), .IN1(P2_sub_858_n169), 
        .Q(P2_sub_858_n168) );
  NAND2X0 P2_sub_858_U165 ( .IN1(P2_sub_858_n167), .IN2(P2_sub_858_n168), 
        .QN(P2_N1746) );
  INVX0 P2_sub_858_U164 ( .ZN(P2_sub_858_n145), .INP(P2_N1505) );
  NAND2X0 P2_sub_858_U163 ( .IN1(n7263), .IN2(P2_sub_858_n145), 
        .QN(P2_sub_858_n165) );
  OR2X1 P2_sub_858_U162 ( .IN2(n7263), .IN1(P2_sub_858_n145), 
        .Q(P2_sub_858_n166) );
  NAND2X0 P2_sub_858_U161 ( .IN1(P2_sub_858_n165), .IN2(P2_sub_858_n166), 
        .QN(P2_sub_858_n159) );
  NAND2X0 P2_sub_858_U160 ( .IN1(n7187), .IN2(P2_sub_858_n164), 
        .QN(P2_sub_858_n160) );
  OR2X1 P2_sub_858_U159 ( .IN2(n7187), .IN1(P2_sub_858_n164), 
        .Q(P2_sub_858_n162) );
  NAND2X0 P2_sub_858_U158 ( .IN1(P2_sub_858_n162), .IN2(P2_sub_858_n163), 
        .QN(P2_sub_858_n161) );
  NAND2X0 P2_sub_858_U157 ( .IN1(P2_sub_858_n160), .IN2(P2_sub_858_n161), 
        .QN(P2_sub_858_n146) );
  NAND2X0 P2_sub_858_U156 ( .IN1(P2_sub_858_n159), .IN2(P2_sub_858_n146), 
        .QN(P2_sub_858_n157) );
  OR2X1 P2_sub_858_U155 ( .IN2(P2_sub_858_n146), .IN1(P2_sub_858_n159), 
        .Q(P2_sub_858_n158) );
  NAND2X0 P2_sub_858_U154 ( .IN1(P2_sub_858_n157), .IN2(P2_sub_858_n158), 
        .QN(P2_N1747) );
  NAND2X0 P2_sub_858_U153 ( .IN1(P2_N5072), .IN2(P2_sub_858_n156), 
        .QN(P2_sub_858_n153) );
  NAND2X0 P2_sub_858_U152 ( .IN1(P2_N1487), .IN2(n7184), .QN(P2_sub_858_n154)
         );
  NAND2X0 P2_sub_858_U151 ( .IN1(P2_sub_858_n153), .IN2(P2_sub_858_n154), 
        .QN(P2_sub_858_n151) );
  NAND2X0 P2_sub_858_U150 ( .IN1(P2_sub_858_n151), .IN2(P2_sub_858_n152), 
        .QN(P2_sub_858_n149) );
  OR2X1 P2_sub_858_U149 ( .IN2(P2_sub_858_n152), .IN1(P2_sub_858_n151), 
        .Q(P2_sub_858_n150) );
  NAND2X0 P2_sub_858_U148 ( .IN1(P2_sub_858_n149), .IN2(P2_sub_858_n150), 
        .QN(P2_N1729) );
  INVX0 P2_sub_858_U147 ( .ZN(P2_sub_858_n135), .INP(P2_N1506) );
  NAND2X0 P2_sub_858_U146 ( .IN1(n7259), .IN2(P2_sub_858_n135), 
        .QN(P2_sub_858_n147) );
  OR2X1 P2_sub_858_U145 ( .IN2(n7259), .IN1(P2_sub_858_n135), 
        .Q(P2_sub_858_n148) );
  NAND2X0 P2_sub_858_U144 ( .IN1(P2_sub_858_n147), .IN2(P2_sub_858_n148), 
        .QN(P2_sub_858_n141) );
  NAND2X0 P2_sub_858_U143 ( .IN1(n7263), .IN2(P2_sub_858_n146), 
        .QN(P2_sub_858_n142) );
  OR2X1 P2_sub_858_U142 ( .IN2(n7263), .IN1(P2_sub_858_n146), 
        .Q(P2_sub_858_n144) );
  NAND2X0 P2_sub_858_U141 ( .IN1(P2_sub_858_n144), .IN2(P2_sub_858_n145), 
        .QN(P2_sub_858_n143) );
  NAND2X0 P2_sub_858_U140 ( .IN1(P2_sub_858_n142), .IN2(P2_sub_858_n143), 
        .QN(P2_sub_858_n136) );
  NAND2X0 P2_sub_858_U139 ( .IN1(P2_sub_858_n141), .IN2(P2_sub_858_n136), 
        .QN(P2_sub_858_n139) );
  OR2X1 P2_sub_858_U138 ( .IN2(P2_sub_858_n136), .IN1(P2_sub_858_n141), 
        .Q(P2_sub_858_n140) );
  NAND2X0 P2_sub_858_U137 ( .IN1(P2_sub_858_n139), .IN2(P2_sub_858_n140), 
        .QN(P2_N1748) );
  INVX0 P2_sub_858_U136 ( .ZN(P2_sub_858_n125), .INP(P2_N1507) );
  NAND2X0 P2_sub_858_U135 ( .IN1(P2_N5092), .IN2(P2_sub_858_n125), 
        .QN(P2_sub_858_n137) );
  OR2X1 P2_sub_858_U134 ( .IN2(P2_N5092), .IN1(P2_sub_858_n125), 
        .Q(P2_sub_858_n138) );
  NAND2X0 P2_sub_858_U133 ( .IN1(P2_sub_858_n137), .IN2(P2_sub_858_n138), 
        .QN(P2_sub_858_n131) );
  NAND2X0 P2_sub_858_U132 ( .IN1(n7259), .IN2(P2_sub_858_n136), 
        .QN(P2_sub_858_n132) );
  OR2X1 P2_sub_858_U131 ( .IN2(n7259), .IN1(P2_sub_858_n136), 
        .Q(P2_sub_858_n134) );
  NAND2X0 P2_sub_858_U130 ( .IN1(P2_sub_858_n134), .IN2(P2_sub_858_n135), 
        .QN(P2_sub_858_n133) );
  NAND2X0 P2_sub_858_U129 ( .IN1(P2_sub_858_n132), .IN2(P2_sub_858_n133), 
        .QN(P2_sub_858_n126) );
  NAND2X0 P2_sub_858_U128 ( .IN1(P2_sub_858_n131), .IN2(P2_sub_858_n126), 
        .QN(P2_sub_858_n129) );
  OR2X1 P2_sub_858_U127 ( .IN2(P2_sub_858_n126), .IN1(P2_sub_858_n131), 
        .Q(P2_sub_858_n130) );
  NAND2X0 P2_sub_858_U126 ( .IN1(P2_sub_858_n129), .IN2(P2_sub_858_n130), 
        .QN(P2_N1749) );
  INVX0 P2_sub_858_U125 ( .ZN(P2_sub_858_n115), .INP(P2_N1508) );
  NAND2X0 P2_sub_858_U124 ( .IN1(n7247), .IN2(P2_sub_858_n115), 
        .QN(P2_sub_858_n127) );
  OR2X1 P2_sub_858_U123 ( .IN2(n7247), .IN1(P2_sub_858_n115), 
        .Q(P2_sub_858_n128) );
  NAND2X0 P2_sub_858_U122 ( .IN1(P2_sub_858_n127), .IN2(P2_sub_858_n128), 
        .QN(P2_sub_858_n121) );
  NAND2X0 P2_sub_858_U121 ( .IN1(P2_N5092), .IN2(P2_sub_858_n126), 
        .QN(P2_sub_858_n122) );
  OR2X1 P2_sub_858_U120 ( .IN2(P2_N5092), .IN1(P2_sub_858_n126), 
        .Q(P2_sub_858_n124) );
  NAND2X0 P2_sub_858_U119 ( .IN1(P2_sub_858_n124), .IN2(P2_sub_858_n125), 
        .QN(P2_sub_858_n123) );
  NAND2X0 P2_sub_858_U118 ( .IN1(P2_sub_858_n122), .IN2(P2_sub_858_n123), 
        .QN(P2_sub_858_n116) );
  NAND2X0 P2_sub_858_U117 ( .IN1(P2_sub_858_n121), .IN2(P2_sub_858_n116), 
        .QN(P2_sub_858_n119) );
  OR2X1 P2_sub_858_U116 ( .IN2(P2_sub_858_n116), .IN1(P2_sub_858_n121), 
        .Q(P2_sub_858_n120) );
  NAND2X0 P2_sub_858_U115 ( .IN1(P2_sub_858_n119), .IN2(P2_sub_858_n120), 
        .QN(P2_N1750) );
  INVX0 P2_sub_858_U114 ( .ZN(P2_sub_858_n105), .INP(P2_N1509) );
  NAND2X0 P2_sub_858_U113 ( .IN1(P2_N5094), .IN2(P2_sub_858_n105), 
        .QN(P2_sub_858_n117) );
  OR2X1 P2_sub_858_U112 ( .IN2(P2_N5094), .IN1(P2_sub_858_n105), 
        .Q(P2_sub_858_n118) );
  NAND2X0 P2_sub_858_U111 ( .IN1(P2_sub_858_n117), .IN2(P2_sub_858_n118), 
        .QN(P2_sub_858_n111) );
  NAND2X0 P2_sub_858_U110 ( .IN1(n7247), .IN2(P2_sub_858_n116), 
        .QN(P2_sub_858_n112) );
  OR2X1 P2_sub_858_U109 ( .IN2(n7247), .IN1(P2_sub_858_n116), 
        .Q(P2_sub_858_n114) );
  NAND2X0 P2_sub_858_U108 ( .IN1(P2_sub_858_n114), .IN2(P2_sub_858_n115), 
        .QN(P2_sub_858_n113) );
  NAND2X0 P2_sub_858_U107 ( .IN1(P2_sub_858_n112), .IN2(P2_sub_858_n113), 
        .QN(P2_sub_858_n106) );
  NAND2X0 P2_sub_858_U106 ( .IN1(P2_sub_858_n111), .IN2(P2_sub_858_n106), 
        .QN(P2_sub_858_n109) );
  OR2X1 P2_sub_858_U105 ( .IN2(P2_sub_858_n106), .IN1(P2_sub_858_n111), 
        .Q(P2_sub_858_n110) );
  NAND2X0 P2_sub_858_U104 ( .IN1(P2_sub_858_n109), .IN2(P2_sub_858_n110), 
        .QN(P2_N1751) );
  INVX0 P2_sub_858_U103 ( .ZN(P2_sub_858_n95), .INP(P2_N1510) );
  NAND2X0 P2_sub_858_U102 ( .IN1(P2_N5095), .IN2(P2_sub_858_n95), 
        .QN(P2_sub_858_n107) );
  OR2X1 P2_sub_858_U101 ( .IN2(P2_N5095), .IN1(P2_sub_858_n95), 
        .Q(P2_sub_858_n108) );
  NAND2X0 P2_sub_858_U100 ( .IN1(P2_sub_858_n107), .IN2(P2_sub_858_n108), 
        .QN(P2_sub_858_n101) );
  NAND2X0 P2_sub_858_U99 ( .IN1(P2_N5094), .IN2(P2_sub_858_n106), 
        .QN(P2_sub_858_n102) );
  OR2X1 P2_sub_858_U98 ( .IN2(P2_N5094), .IN1(P2_sub_858_n106), 
        .Q(P2_sub_858_n104) );
  NAND2X0 P2_sub_858_U97 ( .IN1(P2_sub_858_n104), .IN2(P2_sub_858_n105), 
        .QN(P2_sub_858_n103) );
  NAND2X0 P2_sub_858_U96 ( .IN1(P2_sub_858_n102), .IN2(P2_sub_858_n103), 
        .QN(P2_sub_858_n96) );
  NAND2X0 P2_sub_858_U281 ( .IN1(P2_sub_858_n265), .IN2(P2_sub_858_n266), 
        .QN(P2_sub_858_n32) );
  NAND2X0 P2_sub_858_U280 ( .IN1(n7165), .IN2(P2_sub_858_n32), 
        .QN(P2_sub_858_n262) );
  OR2X1 P2_sub_858_U279 ( .IN2(n7165), .IN1(P2_sub_858_n32), 
        .Q(P2_sub_858_n264) );
  INVX0 P2_sub_858_U278 ( .ZN(P2_sub_858_n35), .INP(P2_N1491) );
  NAND2X0 P2_sub_858_U277 ( .IN1(P2_sub_858_n264), .IN2(P2_sub_858_n35), 
        .QN(P2_sub_858_n263) );
  NAND2X0 P2_sub_858_U276 ( .IN1(P2_sub_858_n262), .IN2(P2_sub_858_n263), 
        .QN(P2_sub_858_n25) );
  NAND2X0 P2_sub_858_U275 ( .IN1(P2_N5077), .IN2(P2_sub_858_n25), 
        .QN(P2_sub_858_n259) );
  OR2X1 P2_sub_858_U274 ( .IN2(P2_N5077), .IN1(P2_sub_858_n25), 
        .Q(P2_sub_858_n261) );
  INVX0 P2_sub_858_U273 ( .ZN(P2_sub_858_n28), .INP(P2_N1492) );
  NAND2X0 P2_sub_858_U272 ( .IN1(P2_sub_858_n261), .IN2(P2_sub_858_n28), 
        .QN(P2_sub_858_n260) );
  NAND2X0 P2_sub_858_U271 ( .IN1(P2_sub_858_n259), .IN2(P2_sub_858_n260), 
        .QN(P2_sub_858_n18) );
  NAND2X0 P2_sub_858_U270 ( .IN1(n7158), .IN2(P2_sub_858_n18), 
        .QN(P2_sub_858_n256) );
  OR2X1 P2_sub_858_U269 ( .IN2(n7158), .IN1(P2_sub_858_n18), 
        .Q(P2_sub_858_n258) );
  INVX0 P2_sub_858_U268 ( .ZN(P2_sub_858_n21), .INP(P2_N1493) );
  NAND2X0 P2_sub_858_U267 ( .IN1(P2_sub_858_n258), .IN2(P2_sub_858_n21), 
        .QN(P2_sub_858_n257) );
  NAND2X0 P2_sub_858_U266 ( .IN1(P2_sub_858_n256), .IN2(P2_sub_858_n257), 
        .QN(P2_sub_858_n11) );
  NAND2X0 P2_sub_858_U265 ( .IN1(n7154), .IN2(P2_sub_858_n11), 
        .QN(P2_sub_858_n253) );
  OR2X1 P2_sub_858_U264 ( .IN2(n7154), .IN1(P2_sub_858_n11), 
        .Q(P2_sub_858_n255) );
  INVX0 P2_sub_858_U263 ( .ZN(P2_sub_858_n14), .INP(P2_N1494) );
  NAND2X0 P2_sub_858_U262 ( .IN1(P2_sub_858_n255), .IN2(P2_sub_858_n14), 
        .QN(P2_sub_858_n254) );
  NAND2X0 P2_sub_858_U261 ( .IN1(P2_sub_858_n253), .IN2(P2_sub_858_n254), 
        .QN(P2_sub_858_n4) );
  NAND2X0 P2_sub_858_U260 ( .IN1(n7151), .IN2(P2_sub_858_n4), 
        .QN(P2_sub_858_n250) );
  OR2X1 P2_sub_858_U259 ( .IN2(n7151), .IN1(P2_sub_858_n4), 
        .Q(P2_sub_858_n252) );
  INVX0 P2_sub_858_U258 ( .ZN(P2_sub_858_n7), .INP(P2_N1495) );
  NAND2X0 P2_sub_858_U257 ( .IN1(P2_sub_858_n252), .IN2(P2_sub_858_n7), 
        .QN(P2_sub_858_n251) );
  NAND2X0 P2_sub_858_U256 ( .IN1(P2_sub_858_n250), .IN2(P2_sub_858_n251), 
        .QN(P2_sub_858_n244) );
  NAND2X0 P2_sub_858_U255 ( .IN1(P2_sub_858_n249), .IN2(P2_sub_858_n244), 
        .QN(P2_sub_858_n247) );
  OR2X1 P2_sub_858_U254 ( .IN2(P2_sub_858_n244), .IN1(P2_sub_858_n249), 
        .Q(P2_sub_858_n248) );
  NAND2X0 P2_sub_858_U253 ( .IN1(P2_sub_858_n247), .IN2(P2_sub_858_n248), 
        .QN(P2_N1738) );
  INVX0 P2_sub_858_U252 ( .ZN(P2_sub_858_n233), .INP(P2_N1497) );
  NAND2X0 P2_sub_858_U251 ( .IN1(P2_N5082), .IN2(P2_sub_858_n233), 
        .QN(P2_sub_858_n245) );
  OR2X1 P2_sub_858_U250 ( .IN2(P2_N5082), .IN1(P2_sub_858_n233), 
        .Q(P2_sub_858_n246) );
  NAND2X0 P2_sub_858_U249 ( .IN1(P2_sub_858_n245), .IN2(P2_sub_858_n246), 
        .QN(P2_sub_858_n239) );
  NAND2X0 P2_sub_858_U248 ( .IN1(P2_N5081), .IN2(P2_sub_858_n244), 
        .QN(P2_sub_858_n240) );
  OR2X1 P2_sub_858_U247 ( .IN2(P2_N5081), .IN1(P2_sub_858_n244), 
        .Q(P2_sub_858_n242) );
  NAND2X0 P2_sub_858_U246 ( .IN1(P2_sub_858_n242), .IN2(P2_sub_858_n243), 
        .QN(P2_sub_858_n241) );
  NAND2X0 P2_sub_858_U245 ( .IN1(P2_sub_858_n240), .IN2(P2_sub_858_n241), 
        .QN(P2_sub_858_n234) );
  NAND2X0 P2_sub_858_U244 ( .IN1(P2_sub_858_n239), .IN2(P2_sub_858_n234), 
        .QN(P2_sub_858_n237) );
  OR2X1 P2_sub_858_U243 ( .IN2(P2_sub_858_n234), .IN1(P2_sub_858_n239), 
        .Q(P2_sub_858_n238) );
  NAND2X0 P2_sub_858_U242 ( .IN1(P2_sub_858_n237), .IN2(P2_sub_858_n238), 
        .QN(P2_N1739) );
  INVX0 P2_sub_858_U241 ( .ZN(P2_sub_858_n223), .INP(P2_N1498) );
  NAND2X0 P2_sub_858_U240 ( .IN1(n7210), .IN2(P2_sub_858_n223), 
        .QN(P2_sub_858_n235) );
  OR2X1 P2_sub_858_U239 ( .IN2(n7210), .IN1(P2_sub_858_n223), 
        .Q(P2_sub_858_n236) );
  NAND2X0 P2_sub_858_U238 ( .IN1(P2_sub_858_n235), .IN2(P2_sub_858_n236), 
        .QN(P2_sub_858_n229) );
  NAND2X0 P2_sub_858_U237 ( .IN1(P2_N5082), .IN2(P2_sub_858_n234), 
        .QN(P2_sub_858_n230) );
  OR2X1 P2_sub_858_U236 ( .IN2(P2_N5082), .IN1(P2_sub_858_n234), 
        .Q(P2_sub_858_n232) );
  NAND2X0 P2_sub_858_U235 ( .IN1(P2_sub_858_n232), .IN2(P2_sub_858_n233), 
        .QN(P2_sub_858_n231) );
  NAND2X0 P2_sub_858_U234 ( .IN1(P2_sub_858_n230), .IN2(P2_sub_858_n231), 
        .QN(P2_sub_858_n224) );
  NAND2X0 P2_sub_858_U233 ( .IN1(P2_sub_858_n229), .IN2(P2_sub_858_n224), 
        .QN(P2_sub_858_n227) );
  OR2X1 P2_sub_858_U232 ( .IN2(P2_sub_858_n224), .IN1(P2_sub_858_n229), 
        .Q(P2_sub_858_n228) );
  NAND2X0 P2_sub_858_U231 ( .IN1(P2_sub_858_n227), .IN2(P2_sub_858_n228), 
        .QN(P2_N1740) );
  INVX0 P2_sub_858_U230 ( .ZN(P2_sub_858_n213), .INP(P2_N1499) );
  NAND2X0 P2_sub_858_U229 ( .IN1(n7209), .IN2(P2_sub_858_n213), 
        .QN(P2_sub_858_n225) );
  OR2X1 P2_sub_858_U228 ( .IN2(n7209), .IN1(P2_sub_858_n213), 
        .Q(P2_sub_858_n226) );
  NAND2X0 P2_sub_858_U227 ( .IN1(P2_sub_858_n225), .IN2(P2_sub_858_n226), 
        .QN(P2_sub_858_n219) );
  NAND2X0 P2_sub_858_U226 ( .IN1(n7210), .IN2(P2_sub_858_n224), 
        .QN(P2_sub_858_n220) );
  OR2X1 P2_sub_858_U225 ( .IN2(n7210), .IN1(P2_sub_858_n224), 
        .Q(P2_sub_858_n222) );
  NAND2X0 P2_sub_858_U224 ( .IN1(P2_sub_858_n222), .IN2(P2_sub_858_n223), 
        .QN(P2_sub_858_n221) );
  NAND2X0 P2_sub_858_U223 ( .IN1(P2_sub_858_n220), .IN2(P2_sub_858_n221), 
        .QN(P2_sub_858_n214) );
  NAND2X0 P2_sub_858_U222 ( .IN1(P2_sub_858_n219), .IN2(P2_sub_858_n214), 
        .QN(P2_sub_858_n217) );
  OR2X1 P2_sub_858_U221 ( .IN2(P2_sub_858_n214), .IN1(P2_sub_858_n219), 
        .Q(P2_sub_858_n218) );
  NAND2X0 P2_sub_858_U220 ( .IN1(P2_sub_858_n217), .IN2(P2_sub_858_n218), 
        .QN(P2_N1741) );
  INVX0 P2_sub_858_U219 ( .ZN(P2_sub_858_n203), .INP(P2_N1500) );
  NAND2X0 P2_sub_858_U218 ( .IN1(n7206), .IN2(P2_sub_858_n203), 
        .QN(P2_sub_858_n215) );
  OR2X1 P2_sub_858_U217 ( .IN2(n7206), .IN1(P2_sub_858_n203), 
        .Q(P2_sub_858_n216) );
  NAND2X0 P2_sub_858_U216 ( .IN1(P2_sub_858_n215), .IN2(P2_sub_858_n216), 
        .QN(P2_sub_858_n209) );
  NAND2X0 P2_sub_858_U215 ( .IN1(n7209), .IN2(P2_sub_858_n214), 
        .QN(P2_sub_858_n210) );
  OR2X1 P2_sub_858_U214 ( .IN2(n7209), .IN1(P2_sub_858_n214), 
        .Q(P2_sub_858_n212) );
  NAND2X0 P2_sub_858_U213 ( .IN1(P2_sub_858_n212), .IN2(P2_sub_858_n213), 
        .QN(P2_sub_858_n211) );
  NAND2X0 P2_sub_858_U212 ( .IN1(P2_sub_858_n210), .IN2(P2_sub_858_n211), 
        .QN(P2_sub_858_n204) );
  NAND2X0 P2_sub_858_U211 ( .IN1(P2_sub_858_n209), .IN2(P2_sub_858_n204), 
        .QN(P2_sub_858_n207) );
  OR2X1 P2_sub_858_U210 ( .IN2(P2_sub_858_n204), .IN1(P2_sub_858_n209), 
        .Q(P2_sub_858_n208) );
  NAND2X0 P2_sub_858_U209 ( .IN1(P2_sub_858_n207), .IN2(P2_sub_858_n208), 
        .QN(P2_N1742) );
  INVX0 P2_sub_858_U208 ( .ZN(P2_sub_858_n193), .INP(P2_N1501) );
  NAND2X0 P2_sub_858_U207 ( .IN1(P2_N5086), .IN2(P2_sub_858_n193), 
        .QN(P2_sub_858_n205) );
  OR2X1 P2_sub_858_U206 ( .IN2(P2_N5086), .IN1(P2_sub_858_n193), 
        .Q(P2_sub_858_n206) );
  NAND2X0 P2_sub_858_U205 ( .IN1(P2_sub_858_n205), .IN2(P2_sub_858_n206), 
        .QN(P2_sub_858_n199) );
  NAND2X0 P2_sub_858_U204 ( .IN1(n7206), .IN2(P2_sub_858_n204), 
        .QN(P2_sub_858_n200) );
  OR2X1 P2_sub_858_U203 ( .IN2(n7206), .IN1(P2_sub_858_n204), 
        .Q(P2_sub_858_n202) );
  NAND2X0 P2_sub_858_U202 ( .IN1(P2_sub_858_n202), .IN2(P2_sub_858_n203), 
        .QN(P2_sub_858_n201) );
  NAND2X0 P2_sub_858_U201 ( .IN1(P2_sub_858_n200), .IN2(P2_sub_858_n201), 
        .QN(P2_sub_858_n194) );
  NAND2X0 P2_sub_858_U200 ( .IN1(P2_sub_858_n199), .IN2(P2_sub_858_n194), 
        .QN(P2_sub_858_n197) );
  OR2X1 P2_sub_858_U199 ( .IN2(P2_sub_858_n194), .IN1(P2_sub_858_n199), 
        .Q(P2_sub_858_n198) );
  NAND2X0 P2_sub_858_U198 ( .IN1(P2_sub_858_n197), .IN2(P2_sub_858_n198), 
        .QN(P2_N1743) );
  INVX0 P2_sub_858_U197 ( .ZN(P2_sub_858_n183), .INP(P2_N1502) );
  NAND2X0 P2_sub_858_U196 ( .IN1(P2_N5087), .IN2(P2_sub_858_n183), 
        .QN(P2_sub_858_n195) );
  OR2X1 P2_sub_858_U195 ( .IN2(P2_N5087), .IN1(P2_sub_858_n183), 
        .Q(P2_sub_858_n196) );
  NAND2X0 P2_sub_858_U194 ( .IN1(P2_sub_858_n195), .IN2(P2_sub_858_n196), 
        .QN(P2_sub_858_n189) );
  NAND2X0 P2_sub_858_U193 ( .IN1(P2_N5086), .IN2(P2_sub_858_n194), 
        .QN(P2_sub_858_n190) );
  OR2X1 P2_sub_858_U192 ( .IN2(P2_N5086), .IN1(P2_sub_858_n194), 
        .Q(P2_sub_858_n192) );
  NAND2X0 P2_sub_858_U191 ( .IN1(P2_sub_858_n192), .IN2(P2_sub_858_n193), 
        .QN(P2_sub_858_n191) );
  NAND2X0 P2_sub_858_U190 ( .IN1(P2_sub_858_n190), .IN2(P2_sub_858_n191), 
        .QN(P2_sub_858_n184) );
  NAND2X0 P2_sub_858_U189 ( .IN1(P2_sub_858_n189), .IN2(P2_sub_858_n184), 
        .QN(P2_sub_858_n187) );
  INVX0 P2_sub_858_U310 ( .ZN(P2_sub_858_n281), .INP(P2_N1486) );
  NOR2X0 P2_sub_858_U309 ( .QN(P2_sub_858_n277), .IN1(P2_sub_858_n281), 
        .IN2(n7035) );
  INVX0 P2_sub_858_U308 ( .ZN(P2_sub_858_n152), .INP(P2_sub_858_n277) );
  NAND2X0 P2_sub_858_U307 ( .IN1(n7035), .IN2(P2_sub_858_n281), 
        .QN(P2_sub_858_n280) );
  NAND2X0 P2_sub_858_U306 ( .IN1(P2_sub_858_n152), .IN2(P2_sub_858_n280), 
        .QN(P2_N1728) );
  INVX0 P2_sub_858_U305 ( .ZN(P2_sub_858_n243), .INP(P2_N1496) );
  NAND2X0 P2_sub_858_U304 ( .IN1(P2_N5081), .IN2(P2_sub_858_n243), 
        .QN(P2_sub_858_n278) );
  OR2X1 P2_sub_858_U303 ( .IN2(P2_N5081), .IN1(P2_sub_858_n243), 
        .Q(P2_sub_858_n279) );
  NAND2X0 P2_sub_858_U302 ( .IN1(P2_sub_858_n278), .IN2(P2_sub_858_n279), 
        .QN(P2_sub_858_n249) );
  NAND2X0 P2_sub_858_U301 ( .IN1(P2_N5072), .IN2(P2_sub_858_n152), 
        .QN(P2_sub_858_n274) );
  NAND2X0 P2_sub_858_U299 ( .IN1(P2_sub_858_n277), .IN2(n7184), 
        .QN(P2_sub_858_n276) );
  INVX0 P2_sub_858_U298 ( .ZN(P2_sub_858_n156), .INP(P2_N1487) );
  NAND2X0 P2_sub_858_U297 ( .IN1(P2_sub_858_n276), .IN2(P2_sub_858_n156), 
        .QN(P2_sub_858_n275) );
  NAND2X0 P2_sub_858_U296 ( .IN1(P2_sub_858_n274), .IN2(P2_sub_858_n275), 
        .QN(P2_sub_858_n53) );
  NAND2X0 P2_sub_858_U295 ( .IN1(P2_N5073), .IN2(P2_sub_858_n53), 
        .QN(P2_sub_858_n271) );
  OR2X1 P2_sub_858_U294 ( .IN2(P2_N5073), .IN1(P2_sub_858_n53), 
        .Q(P2_sub_858_n273) );
  INVX0 P2_sub_858_U293 ( .ZN(P2_sub_858_n56), .INP(P2_N1488) );
  NAND2X0 P2_sub_858_U292 ( .IN1(P2_sub_858_n273), .IN2(P2_sub_858_n56), 
        .QN(P2_sub_858_n272) );
  NAND2X0 P2_sub_858_U291 ( .IN1(P2_sub_858_n271), .IN2(P2_sub_858_n272), 
        .QN(P2_sub_858_n46) );
  NAND2X0 P2_sub_858_U290 ( .IN1(P2_N5074), .IN2(P2_sub_858_n46), 
        .QN(P2_sub_858_n268) );
  OR2X1 P2_sub_858_U289 ( .IN2(P2_N5074), .IN1(P2_sub_858_n46), 
        .Q(P2_sub_858_n270) );
  INVX0 P2_sub_858_U288 ( .ZN(P2_sub_858_n49), .INP(P2_N1489) );
  NAND2X0 P2_sub_858_U287 ( .IN1(P2_sub_858_n270), .IN2(P2_sub_858_n49), 
        .QN(P2_sub_858_n269) );
  NAND2X0 P2_sub_858_U286 ( .IN1(P2_sub_858_n268), .IN2(P2_sub_858_n269), 
        .QN(P2_sub_858_n39) );
  NAND2X0 P2_sub_858_U285 ( .IN1(n7173), .IN2(P2_sub_858_n39), 
        .QN(P2_sub_858_n265) );
  OR2X1 P2_sub_858_U284 ( .IN2(n7173), .IN1(P2_sub_858_n39), 
        .Q(P2_sub_858_n267) );
  INVX0 P2_sub_858_U283 ( .ZN(P2_sub_858_n42), .INP(P2_N1490) );
  NAND2X0 P2_sub_858_U282 ( .IN1(P2_sub_858_n267), .IN2(P2_sub_858_n42), 
        .QN(P2_sub_858_n266) );
  NAND2X0 P2_sub_878_U33 ( .IN1(P2_sub_878_n38), .IN2(P2_sub_878_n39), 
        .QN(P2_sub_878_n36) );
  OR2X1 P2_sub_878_U32 ( .IN2(P2_sub_878_n39), .IN1(P2_sub_878_n38), 
        .Q(P2_sub_878_n37) );
  NAND2X0 P2_sub_878_U31 ( .IN1(P2_sub_878_n36), .IN2(P2_sub_878_n37), 
        .QN(P2_N2105) );
  NAND2X0 P2_sub_878_U30 ( .IN1(n7165), .IN2(P2_sub_878_n35), 
        .QN(P2_sub_878_n33) );
  OR2X1 P2_sub_878_U29 ( .IN2(n7165), .IN1(P2_sub_878_n35), .Q(P2_sub_878_n34)
         );
  NAND2X0 P2_sub_878_U28 ( .IN1(P2_sub_878_n33), .IN2(P2_sub_878_n34), 
        .QN(P2_sub_878_n31) );
  NAND2X0 P2_sub_878_U27 ( .IN1(P2_sub_878_n31), .IN2(P2_sub_878_n32), 
        .QN(P2_sub_878_n29) );
  OR2X1 P2_sub_878_U26 ( .IN2(P2_sub_878_n32), .IN1(P2_sub_878_n31), 
        .Q(P2_sub_878_n30) );
  NAND2X0 P2_sub_878_U25 ( .IN1(P2_sub_878_n29), .IN2(P2_sub_878_n30), 
        .QN(P2_N2106) );
  NAND2X0 P2_sub_878_U24 ( .IN1(P2_N5077), .IN2(P2_sub_878_n28), 
        .QN(P2_sub_878_n26) );
  OR2X1 P2_sub_878_U23 ( .IN2(P2_N5077), .IN1(P2_sub_878_n28), 
        .Q(P2_sub_878_n27) );
  NAND2X0 P2_sub_878_U22 ( .IN1(P2_sub_878_n26), .IN2(P2_sub_878_n27), 
        .QN(P2_sub_878_n24) );
  NAND2X0 P2_sub_878_U21 ( .IN1(P2_sub_878_n24), .IN2(P2_sub_878_n25), 
        .QN(P2_sub_878_n22) );
  OR2X1 P2_sub_878_U20 ( .IN2(P2_sub_878_n25), .IN1(P2_sub_878_n24), 
        .Q(P2_sub_878_n23) );
  NAND2X0 P2_sub_878_U19 ( .IN1(P2_sub_878_n22), .IN2(P2_sub_878_n23), 
        .QN(P2_N2107) );
  NAND2X0 P2_sub_878_U18 ( .IN1(P2_N5078), .IN2(P2_sub_878_n21), 
        .QN(P2_sub_878_n19) );
  OR2X1 P2_sub_878_U17 ( .IN2(P2_N5078), .IN1(P2_sub_878_n21), 
        .Q(P2_sub_878_n20) );
  NAND2X0 P2_sub_878_U16 ( .IN1(P2_sub_878_n19), .IN2(P2_sub_878_n20), 
        .QN(P2_sub_878_n17) );
  NAND2X0 P2_sub_878_U15 ( .IN1(P2_sub_878_n17), .IN2(P2_sub_878_n18), 
        .QN(P2_sub_878_n15) );
  OR2X1 P2_sub_878_U14 ( .IN2(P2_sub_878_n18), .IN1(P2_sub_878_n17), 
        .Q(P2_sub_878_n16) );
  NAND2X0 P2_sub_878_U13 ( .IN1(P2_sub_878_n15), .IN2(P2_sub_878_n16), 
        .QN(P2_N2108) );
  NAND2X0 P2_sub_878_U12 ( .IN1(P2_N5079), .IN2(P2_sub_878_n14), 
        .QN(P2_sub_878_n12) );
  OR2X1 P2_sub_878_U11 ( .IN2(P2_N5079), .IN1(P2_sub_878_n14), 
        .Q(P2_sub_878_n13) );
  NAND2X0 P2_sub_878_U10 ( .IN1(P2_sub_878_n12), .IN2(P2_sub_878_n13), 
        .QN(P2_sub_878_n10) );
  NAND2X0 P2_sub_878_U9 ( .IN1(P2_sub_878_n10), .IN2(P2_sub_878_n11), 
        .QN(P2_sub_878_n8) );
  OR2X1 P2_sub_878_U8 ( .IN2(P2_sub_878_n11), .IN1(P2_sub_878_n10), 
        .Q(P2_sub_878_n9) );
  NAND2X0 P2_sub_878_U7 ( .IN1(P2_sub_878_n8), .IN2(P2_sub_878_n9), 
        .QN(P2_N2109) );
  NAND2X0 P2_sub_878_U6 ( .IN1(n7151), .IN2(P2_sub_878_n7), .QN(P2_sub_878_n5)
         );
  OR2X1 P2_sub_878_U5 ( .IN2(n7151), .IN1(P2_sub_878_n7), .Q(P2_sub_878_n6) );
  NAND2X0 P2_sub_878_U4 ( .IN1(P2_sub_878_n5), .IN2(P2_sub_878_n6), 
        .QN(P2_sub_878_n3) );
  NAND2X0 P2_sub_878_U3 ( .IN1(P2_sub_878_n3), .IN2(P2_sub_878_n4), 
        .QN(P2_sub_878_n1) );
  OR2X1 P2_sub_878_U2 ( .IN2(P2_sub_878_n4), .IN1(P2_sub_878_n3), 
        .Q(P2_sub_878_n2) );
  NAND2X0 P2_sub_878_U1 ( .IN1(P2_sub_878_n1), .IN2(P2_sub_878_n2), 
        .QN(P2_N2110) );
  NAND2X0 P2_sub_878_U126 ( .IN1(P2_sub_878_n129), .IN2(P2_sub_878_n130), 
        .QN(P2_N2122) );
  INVX0 P2_sub_878_U125 ( .ZN(P2_sub_878_n115), .INP(P2_N1881) );
  NAND2X0 P2_sub_878_U124 ( .IN1(n7247), .IN2(P2_sub_878_n115), 
        .QN(P2_sub_878_n127) );
  OR2X1 P2_sub_878_U123 ( .IN2(n7247), .IN1(P2_sub_878_n115), 
        .Q(P2_sub_878_n128) );
  NAND2X0 P2_sub_878_U122 ( .IN1(P2_sub_878_n127), .IN2(P2_sub_878_n128), 
        .QN(P2_sub_878_n121) );
  NAND2X0 P2_sub_878_U121 ( .IN1(n7252), .IN2(P2_sub_878_n126), 
        .QN(P2_sub_878_n122) );
  OR2X1 P2_sub_878_U120 ( .IN2(n7252), .IN1(P2_sub_878_n126), 
        .Q(P2_sub_878_n124) );
  NAND2X0 P2_sub_878_U119 ( .IN1(P2_sub_878_n124), .IN2(P2_sub_878_n125), 
        .QN(P2_sub_878_n123) );
  NAND2X0 P2_sub_878_U118 ( .IN1(P2_sub_878_n122), .IN2(P2_sub_878_n123), 
        .QN(P2_sub_878_n116) );
  NAND2X0 P2_sub_878_U117 ( .IN1(P2_sub_878_n121), .IN2(P2_sub_878_n116), 
        .QN(P2_sub_878_n119) );
  OR2X1 P2_sub_878_U116 ( .IN2(P2_sub_878_n116), .IN1(P2_sub_878_n121), 
        .Q(P2_sub_878_n120) );
  NAND2X0 P2_sub_878_U115 ( .IN1(P2_sub_878_n119), .IN2(P2_sub_878_n120), 
        .QN(P2_N2123) );
  INVX0 P2_sub_878_U114 ( .ZN(P2_sub_878_n105), .INP(P2_N1882) );
  NAND2X0 P2_sub_878_U113 ( .IN1(P2_N5094), .IN2(P2_sub_878_n105), 
        .QN(P2_sub_878_n117) );
  OR2X1 P2_sub_878_U112 ( .IN2(P2_N5094), .IN1(P2_sub_878_n105), 
        .Q(P2_sub_878_n118) );
  NAND2X0 P2_sub_878_U111 ( .IN1(P2_sub_878_n117), .IN2(P2_sub_878_n118), 
        .QN(P2_sub_878_n111) );
  NAND2X0 P2_sub_878_U110 ( .IN1(n7247), .IN2(P2_sub_878_n116), 
        .QN(P2_sub_878_n112) );
  OR2X1 P2_sub_878_U109 ( .IN2(n7247), .IN1(P2_sub_878_n116), 
        .Q(P2_sub_878_n114) );
  NAND2X0 P2_sub_878_U108 ( .IN1(P2_sub_878_n114), .IN2(P2_sub_878_n115), 
        .QN(P2_sub_878_n113) );
  NAND2X0 P2_sub_878_U107 ( .IN1(P2_sub_878_n112), .IN2(P2_sub_878_n113), 
        .QN(P2_sub_878_n106) );
  NAND2X0 P2_sub_878_U106 ( .IN1(P2_sub_878_n111), .IN2(P2_sub_878_n106), 
        .QN(P2_sub_878_n109) );
  OR2X1 P2_sub_878_U105 ( .IN2(P2_sub_878_n106), .IN1(P2_sub_878_n111), 
        .Q(P2_sub_878_n110) );
  NAND2X0 P2_sub_878_U104 ( .IN1(P2_sub_878_n109), .IN2(P2_sub_878_n110), 
        .QN(P2_N2124) );
  INVX0 P2_sub_878_U103 ( .ZN(P2_sub_878_n95), .INP(P2_N1883) );
  NAND2X0 P2_sub_878_U102 ( .IN1(P2_N5095), .IN2(P2_sub_878_n95), 
        .QN(P2_sub_878_n107) );
  OR2X1 P2_sub_878_U101 ( .IN2(P2_N5095), .IN1(P2_sub_878_n95), 
        .Q(P2_sub_878_n108) );
  NAND2X0 P2_sub_878_U100 ( .IN1(P2_sub_878_n107), .IN2(P2_sub_878_n108), 
        .QN(P2_sub_878_n101) );
  NAND2X0 P2_sub_878_U99 ( .IN1(P2_N5094), .IN2(P2_sub_878_n106), 
        .QN(P2_sub_878_n102) );
  OR2X1 P2_sub_878_U98 ( .IN2(P2_N5094), .IN1(P2_sub_878_n106), 
        .Q(P2_sub_878_n104) );
  NAND2X0 P2_sub_878_U97 ( .IN1(P2_sub_878_n104), .IN2(P2_sub_878_n105), 
        .QN(P2_sub_878_n103) );
  NAND2X0 P2_sub_878_U96 ( .IN1(P2_sub_878_n102), .IN2(P2_sub_878_n103), 
        .QN(P2_sub_878_n96) );
  NAND2X0 P2_sub_878_U95 ( .IN1(P2_sub_878_n101), .IN2(P2_sub_878_n96), 
        .QN(P2_sub_878_n99) );
  OR2X1 P2_sub_878_U94 ( .IN2(P2_sub_878_n96), .IN1(P2_sub_878_n101), 
        .Q(P2_sub_878_n100) );
  NAND2X0 P2_sub_878_U93 ( .IN1(P2_sub_878_n99), .IN2(P2_sub_878_n100), 
        .QN(P2_N2125) );
  INVX0 P2_sub_878_U92 ( .ZN(P2_sub_878_n85), .INP(P2_N1884) );
  NAND2X0 P2_sub_878_U91 ( .IN1(n7237), .IN2(P2_sub_878_n85), 
        .QN(P2_sub_878_n97) );
  OR2X1 P2_sub_878_U90 ( .IN2(n7237), .IN1(P2_sub_878_n85), .Q(P2_sub_878_n98)
         );
  NAND2X0 P2_sub_878_U89 ( .IN1(P2_sub_878_n97), .IN2(P2_sub_878_n98), 
        .QN(P2_sub_878_n91) );
  NAND2X0 P2_sub_878_U88 ( .IN1(P2_N5095), .IN2(P2_sub_878_n96), 
        .QN(P2_sub_878_n92) );
  OR2X1 P2_sub_878_U87 ( .IN2(P2_N5095), .IN1(P2_sub_878_n96), 
        .Q(P2_sub_878_n94) );
  NAND2X0 P2_sub_878_U86 ( .IN1(P2_sub_878_n94), .IN2(P2_sub_878_n95), 
        .QN(P2_sub_878_n93) );
  NAND2X0 P2_sub_878_U85 ( .IN1(P2_sub_878_n92), .IN2(P2_sub_878_n93), 
        .QN(P2_sub_878_n86) );
  NAND2X0 P2_sub_878_U84 ( .IN1(P2_sub_878_n91), .IN2(P2_sub_878_n86), 
        .QN(P2_sub_878_n89) );
  OR2X1 P2_sub_878_U83 ( .IN2(P2_sub_878_n86), .IN1(P2_sub_878_n91), 
        .Q(P2_sub_878_n90) );
  NAND2X0 P2_sub_878_U82 ( .IN1(P2_sub_878_n89), .IN2(P2_sub_878_n90), 
        .QN(P2_N2126) );
  INVX0 P2_sub_878_U81 ( .ZN(P2_sub_878_n75), .INP(P2_N1885) );
  NAND2X0 P2_sub_878_U80 ( .IN1(n7231), .IN2(P2_sub_878_n75), 
        .QN(P2_sub_878_n87) );
  OR2X1 P2_sub_878_U79 ( .IN2(n7231), .IN1(P2_sub_878_n75), .Q(P2_sub_878_n88)
         );
  NAND2X0 P2_sub_878_U78 ( .IN1(P2_sub_878_n87), .IN2(P2_sub_878_n88), 
        .QN(P2_sub_878_n81) );
  NAND2X0 P2_sub_878_U77 ( .IN1(n7237), .IN2(P2_sub_878_n86), 
        .QN(P2_sub_878_n82) );
  OR2X1 P2_sub_878_U76 ( .IN2(n7237), .IN1(P2_sub_878_n86), .Q(P2_sub_878_n84)
         );
  NAND2X0 P2_sub_878_U75 ( .IN1(P2_sub_878_n84), .IN2(P2_sub_878_n85), 
        .QN(P2_sub_878_n83) );
  NAND2X0 P2_sub_878_U74 ( .IN1(P2_sub_878_n82), .IN2(P2_sub_878_n83), 
        .QN(P2_sub_878_n76) );
  NAND2X0 P2_sub_878_U73 ( .IN1(P2_sub_878_n81), .IN2(P2_sub_878_n76), 
        .QN(P2_sub_878_n79) );
  OR2X1 P2_sub_878_U72 ( .IN2(P2_sub_878_n76), .IN1(P2_sub_878_n81), 
        .Q(P2_sub_878_n80) );
  NAND2X0 P2_sub_878_U71 ( .IN1(P2_sub_878_n79), .IN2(P2_sub_878_n80), 
        .QN(P2_N2127) );
  INVX0 P2_sub_878_U70 ( .ZN(P2_sub_878_n64), .INP(P2_N1886) );
  NAND2X0 P2_sub_878_U69 ( .IN1(n7227), .IN2(P2_sub_878_n64), 
        .QN(P2_sub_878_n77) );
  OR2X1 P2_sub_878_U68 ( .IN2(n7227), .IN1(P2_sub_878_n64), .Q(P2_sub_878_n78)
         );
  NAND2X0 P2_sub_878_U67 ( .IN1(P2_sub_878_n77), .IN2(P2_sub_878_n78), 
        .QN(P2_sub_878_n71) );
  NAND2X0 P2_sub_878_U66 ( .IN1(n7231), .IN2(P2_sub_878_n76), 
        .QN(P2_sub_878_n72) );
  OR2X1 P2_sub_878_U65 ( .IN2(n7231), .IN1(P2_sub_878_n76), .Q(P2_sub_878_n74)
         );
  NAND2X0 P2_sub_878_U64 ( .IN1(P2_sub_878_n74), .IN2(P2_sub_878_n75), 
        .QN(P2_sub_878_n73) );
  NAND2X0 P2_sub_878_U63 ( .IN1(P2_sub_878_n72), .IN2(P2_sub_878_n73), 
        .QN(P2_sub_878_n65) );
  NAND2X0 P2_sub_878_U62 ( .IN1(P2_sub_878_n71), .IN2(P2_sub_878_n65), 
        .QN(P2_sub_878_n69) );
  OR2X1 P2_sub_878_U61 ( .IN2(P2_sub_878_n65), .IN1(P2_sub_878_n71), 
        .Q(P2_sub_878_n70) );
  NAND2X0 P2_sub_878_U60 ( .IN1(P2_sub_878_n69), .IN2(P2_sub_878_n70), 
        .QN(P2_N2128) );
  OR2X1 P2_sub_878_U58 ( .IN2(P2_N1887), .IN1(n7222), .Q(P2_sub_878_n66) );
  NAND2X0 P2_sub_878_U57 ( .IN1(P2_N1887), .IN2(n7222), .QN(P2_sub_878_n67) );
  NAND2X0 P2_sub_878_U56 ( .IN1(P2_sub_878_n66), .IN2(P2_sub_878_n67), 
        .QN(P2_sub_878_n60) );
  NAND2X0 P2_sub_878_U55 ( .IN1(n7227), .IN2(P2_sub_878_n65), 
        .QN(P2_sub_878_n61) );
  OR2X1 P2_sub_878_U54 ( .IN2(n7227), .IN1(P2_sub_878_n65), .Q(P2_sub_878_n63)
         );
  NAND2X0 P2_sub_878_U53 ( .IN1(P2_sub_878_n63), .IN2(P2_sub_878_n64), 
        .QN(P2_sub_878_n62) );
  NAND2X0 P2_sub_878_U52 ( .IN1(P2_sub_878_n61), .IN2(P2_sub_878_n62), 
        .QN(P2_sub_878_n59) );
  NAND2X0 P2_sub_878_U51 ( .IN1(P2_sub_878_n60), .IN2(P2_sub_878_n59), 
        .QN(P2_sub_878_n57) );
  OR2X1 P2_sub_878_U50 ( .IN2(P2_sub_878_n60), .IN1(P2_sub_878_n59), 
        .Q(P2_sub_878_n58) );
  NAND2X0 P2_sub_878_U49 ( .IN1(P2_sub_878_n57), .IN2(P2_sub_878_n58), 
        .QN(P2_N2129) );
  NAND2X0 P2_sub_878_U48 ( .IN1(n7181), .IN2(P2_sub_878_n56), 
        .QN(P2_sub_878_n54) );
  OR2X1 P2_sub_878_U47 ( .IN2(n7181), .IN1(P2_sub_878_n56), .Q(P2_sub_878_n55)
         );
  NAND2X0 P2_sub_878_U46 ( .IN1(P2_sub_878_n54), .IN2(P2_sub_878_n55), 
        .QN(P2_sub_878_n52) );
  NAND2X0 P2_sub_878_U45 ( .IN1(P2_sub_878_n52), .IN2(P2_sub_878_n53), 
        .QN(P2_sub_878_n50) );
  OR2X1 P2_sub_878_U44 ( .IN2(P2_sub_878_n53), .IN1(P2_sub_878_n52), 
        .Q(P2_sub_878_n51) );
  NAND2X0 P2_sub_878_U43 ( .IN1(P2_sub_878_n50), .IN2(P2_sub_878_n51), 
        .QN(P2_N2103) );
  NAND2X0 P2_sub_878_U42 ( .IN1(n7177), .IN2(P2_sub_878_n49), 
        .QN(P2_sub_878_n47) );
  OR2X1 P2_sub_878_U41 ( .IN2(n7177), .IN1(P2_sub_878_n49), .Q(P2_sub_878_n48)
         );
  NAND2X0 P2_sub_878_U40 ( .IN1(P2_sub_878_n47), .IN2(P2_sub_878_n48), 
        .QN(P2_sub_878_n45) );
  NAND2X0 P2_sub_878_U39 ( .IN1(P2_sub_878_n45), .IN2(P2_sub_878_n46), 
        .QN(P2_sub_878_n43) );
  OR2X1 P2_sub_878_U38 ( .IN2(P2_sub_878_n46), .IN1(P2_sub_878_n45), 
        .Q(P2_sub_878_n44) );
  NAND2X0 P2_sub_878_U37 ( .IN1(P2_sub_878_n43), .IN2(P2_sub_878_n44), 
        .QN(P2_N2104) );
  NAND2X0 P2_sub_878_U36 ( .IN1(n7173), .IN2(P2_sub_878_n42), 
        .QN(P2_sub_878_n40) );
  OR2X1 P2_sub_878_U35 ( .IN2(n7173), .IN1(P2_sub_878_n42), .Q(P2_sub_878_n41)
         );
  NAND2X0 P2_sub_878_U34 ( .IN1(P2_sub_878_n40), .IN2(P2_sub_878_n41), 
        .QN(P2_sub_878_n38) );
  INVX0 P2_sub_878_U219 ( .ZN(P2_sub_878_n203), .INP(P2_N1873) );
  NAND2X0 P2_sub_878_U218 ( .IN1(P2_N5085), .IN2(P2_sub_878_n203), 
        .QN(P2_sub_878_n215) );
  OR2X1 P2_sub_878_U217 ( .IN2(P2_N5085), .IN1(P2_sub_878_n203), 
        .Q(P2_sub_878_n216) );
  NAND2X0 P2_sub_878_U216 ( .IN1(P2_sub_878_n215), .IN2(P2_sub_878_n216), 
        .QN(P2_sub_878_n209) );
  NAND2X0 P2_sub_878_U215 ( .IN1(P2_N5084), .IN2(P2_sub_878_n214), 
        .QN(P2_sub_878_n210) );
  OR2X1 P2_sub_878_U214 ( .IN2(P2_N5084), .IN1(P2_sub_878_n214), 
        .Q(P2_sub_878_n212) );
  NAND2X0 P2_sub_878_U213 ( .IN1(P2_sub_878_n212), .IN2(P2_sub_878_n213), 
        .QN(P2_sub_878_n211) );
  NAND2X0 P2_sub_878_U212 ( .IN1(P2_sub_878_n210), .IN2(P2_sub_878_n211), 
        .QN(P2_sub_878_n204) );
  NAND2X0 P2_sub_878_U211 ( .IN1(P2_sub_878_n209), .IN2(P2_sub_878_n204), 
        .QN(P2_sub_878_n207) );
  OR2X1 P2_sub_878_U210 ( .IN2(P2_sub_878_n204), .IN1(P2_sub_878_n209), 
        .Q(P2_sub_878_n208) );
  NAND2X0 P2_sub_878_U209 ( .IN1(P2_sub_878_n207), .IN2(P2_sub_878_n208), 
        .QN(P2_N2115) );
  INVX0 P2_sub_878_U208 ( .ZN(P2_sub_878_n193), .INP(P2_N1874) );
  NAND2X0 P2_sub_878_U207 ( .IN1(P2_N5086), .IN2(P2_sub_878_n193), 
        .QN(P2_sub_878_n205) );
  OR2X1 P2_sub_878_U206 ( .IN2(P2_N5086), .IN1(P2_sub_878_n193), 
        .Q(P2_sub_878_n206) );
  NAND2X0 P2_sub_878_U205 ( .IN1(P2_sub_878_n205), .IN2(P2_sub_878_n206), 
        .QN(P2_sub_878_n199) );
  NAND2X0 P2_sub_878_U204 ( .IN1(P2_N5085), .IN2(P2_sub_878_n204), 
        .QN(P2_sub_878_n200) );
  OR2X1 P2_sub_878_U203 ( .IN2(P2_N5085), .IN1(P2_sub_878_n204), 
        .Q(P2_sub_878_n202) );
  NAND2X0 P2_sub_878_U202 ( .IN1(P2_sub_878_n202), .IN2(P2_sub_878_n203), 
        .QN(P2_sub_878_n201) );
  NAND2X0 P2_sub_878_U201 ( .IN1(P2_sub_878_n200), .IN2(P2_sub_878_n201), 
        .QN(P2_sub_878_n194) );
  NAND2X0 P2_sub_878_U200 ( .IN1(P2_sub_878_n199), .IN2(P2_sub_878_n194), 
        .QN(P2_sub_878_n197) );
  OR2X1 P2_sub_878_U199 ( .IN2(P2_sub_878_n194), .IN1(P2_sub_878_n199), 
        .Q(P2_sub_878_n198) );
  NAND2X0 P2_sub_878_U198 ( .IN1(P2_sub_878_n197), .IN2(P2_sub_878_n198), 
        .QN(P2_N2116) );
  INVX0 P2_sub_878_U197 ( .ZN(P2_sub_878_n183), .INP(P2_N1875) );
  NAND2X0 P2_sub_878_U196 ( .IN1(P2_N5087), .IN2(P2_sub_878_n183), 
        .QN(P2_sub_878_n195) );
  OR2X1 P2_sub_878_U195 ( .IN2(P2_N5087), .IN1(P2_sub_878_n183), 
        .Q(P2_sub_878_n196) );
  NAND2X0 P2_sub_878_U194 ( .IN1(P2_sub_878_n195), .IN2(P2_sub_878_n196), 
        .QN(P2_sub_878_n189) );
  NAND2X0 P2_sub_878_U193 ( .IN1(P2_N5086), .IN2(P2_sub_878_n194), 
        .QN(P2_sub_878_n190) );
  OR2X1 P2_sub_878_U192 ( .IN2(P2_N5086), .IN1(P2_sub_878_n194), 
        .Q(P2_sub_878_n192) );
  NAND2X0 P2_sub_878_U191 ( .IN1(P2_sub_878_n192), .IN2(P2_sub_878_n193), 
        .QN(P2_sub_878_n191) );
  NAND2X0 P2_sub_878_U190 ( .IN1(P2_sub_878_n190), .IN2(P2_sub_878_n191), 
        .QN(P2_sub_878_n184) );
  NAND2X0 P2_sub_878_U189 ( .IN1(P2_sub_878_n189), .IN2(P2_sub_878_n184), 
        .QN(P2_sub_878_n187) );
  OR2X1 P2_sub_878_U188 ( .IN2(P2_sub_878_n184), .IN1(P2_sub_878_n189), 
        .Q(P2_sub_878_n188) );
  NAND2X0 P2_sub_878_U187 ( .IN1(P2_sub_878_n187), .IN2(P2_sub_878_n188), 
        .QN(P2_N2117) );
  INVX0 P2_sub_878_U186 ( .ZN(P2_sub_878_n173), .INP(P2_N1876) );
  NAND2X0 P2_sub_878_U185 ( .IN1(n7194), .IN2(P2_sub_878_n173), 
        .QN(P2_sub_878_n185) );
  OR2X1 P2_sub_878_U184 ( .IN2(n7194), .IN1(P2_sub_878_n173), 
        .Q(P2_sub_878_n186) );
  NAND2X0 P2_sub_878_U183 ( .IN1(P2_sub_878_n185), .IN2(P2_sub_878_n186), 
        .QN(P2_sub_878_n179) );
  NAND2X0 P2_sub_878_U182 ( .IN1(P2_N5087), .IN2(P2_sub_878_n184), 
        .QN(P2_sub_878_n180) );
  OR2X1 P2_sub_878_U181 ( .IN2(P2_N5087), .IN1(P2_sub_878_n184), 
        .Q(P2_sub_878_n182) );
  NAND2X0 P2_sub_878_U180 ( .IN1(P2_sub_878_n182), .IN2(P2_sub_878_n183), 
        .QN(P2_sub_878_n181) );
  NAND2X0 P2_sub_878_U179 ( .IN1(P2_sub_878_n180), .IN2(P2_sub_878_n181), 
        .QN(P2_sub_878_n174) );
  NAND2X0 P2_sub_878_U178 ( .IN1(P2_sub_878_n179), .IN2(P2_sub_878_n174), 
        .QN(P2_sub_878_n177) );
  OR2X1 P2_sub_878_U177 ( .IN2(P2_sub_878_n174), .IN1(P2_sub_878_n179), 
        .Q(P2_sub_878_n178) );
  NAND2X0 P2_sub_878_U176 ( .IN1(P2_sub_878_n177), .IN2(P2_sub_878_n178), 
        .QN(P2_N2118) );
  INVX0 P2_sub_878_U175 ( .ZN(P2_sub_878_n163), .INP(P2_N1877) );
  NAND2X0 P2_sub_878_U174 ( .IN1(P2_N5089), .IN2(P2_sub_878_n163), 
        .QN(P2_sub_878_n175) );
  OR2X1 P2_sub_878_U173 ( .IN2(P2_N5089), .IN1(P2_sub_878_n163), 
        .Q(P2_sub_878_n176) );
  NAND2X0 P2_sub_878_U172 ( .IN1(P2_sub_878_n175), .IN2(P2_sub_878_n176), 
        .QN(P2_sub_878_n169) );
  NAND2X0 P2_sub_878_U171 ( .IN1(n7194), .IN2(P2_sub_878_n174), 
        .QN(P2_sub_878_n170) );
  OR2X1 P2_sub_878_U170 ( .IN2(n7194), .IN1(P2_sub_878_n174), 
        .Q(P2_sub_878_n172) );
  NAND2X0 P2_sub_878_U169 ( .IN1(P2_sub_878_n172), .IN2(P2_sub_878_n173), 
        .QN(P2_sub_878_n171) );
  NAND2X0 P2_sub_878_U168 ( .IN1(P2_sub_878_n170), .IN2(P2_sub_878_n171), 
        .QN(P2_sub_878_n164) );
  NAND2X0 P2_sub_878_U167 ( .IN1(P2_sub_878_n169), .IN2(P2_sub_878_n164), 
        .QN(P2_sub_878_n167) );
  OR2X1 P2_sub_878_U166 ( .IN2(P2_sub_878_n164), .IN1(P2_sub_878_n169), 
        .Q(P2_sub_878_n168) );
  NAND2X0 P2_sub_878_U165 ( .IN1(P2_sub_878_n167), .IN2(P2_sub_878_n168), 
        .QN(P2_N2119) );
  INVX0 P2_sub_878_U164 ( .ZN(P2_sub_878_n145), .INP(P2_N1878) );
  NAND2X0 P2_sub_878_U163 ( .IN1(P2_N5090), .IN2(P2_sub_878_n145), 
        .QN(P2_sub_878_n165) );
  OR2X1 P2_sub_878_U162 ( .IN2(P2_N5090), .IN1(P2_sub_878_n145), 
        .Q(P2_sub_878_n166) );
  NAND2X0 P2_sub_878_U161 ( .IN1(P2_sub_878_n165), .IN2(P2_sub_878_n166), 
        .QN(P2_sub_878_n159) );
  NAND2X0 P2_sub_878_U160 ( .IN1(P2_N5089), .IN2(P2_sub_878_n164), 
        .QN(P2_sub_878_n160) );
  OR2X1 P2_sub_878_U159 ( .IN2(P2_N5089), .IN1(P2_sub_878_n164), 
        .Q(P2_sub_878_n162) );
  NAND2X0 P2_sub_878_U158 ( .IN1(P2_sub_878_n162), .IN2(P2_sub_878_n163), 
        .QN(P2_sub_878_n161) );
  NAND2X0 P2_sub_878_U157 ( .IN1(P2_sub_878_n160), .IN2(P2_sub_878_n161), 
        .QN(P2_sub_878_n146) );
  NAND2X0 P2_sub_878_U156 ( .IN1(P2_sub_878_n159), .IN2(P2_sub_878_n146), 
        .QN(P2_sub_878_n157) );
  OR2X1 P2_sub_878_U155 ( .IN2(P2_sub_878_n146), .IN1(P2_sub_878_n159), 
        .Q(P2_sub_878_n158) );
  NAND2X0 P2_sub_878_U154 ( .IN1(P2_sub_878_n157), .IN2(P2_sub_878_n158), 
        .QN(P2_N2120) );
  NAND2X0 P2_sub_878_U153 ( .IN1(P2_N5072), .IN2(P2_sub_878_n156), 
        .QN(P2_sub_878_n153) );
  NAND2X0 P2_sub_878_U152 ( .IN1(P2_N1860), .IN2(n7186), .QN(P2_sub_878_n154)
         );
  NAND2X0 P2_sub_878_U151 ( .IN1(P2_sub_878_n153), .IN2(P2_sub_878_n154), 
        .QN(P2_sub_878_n151) );
  NAND2X0 P2_sub_878_U150 ( .IN1(P2_sub_878_n151), .IN2(P2_sub_878_n152), 
        .QN(P2_sub_878_n149) );
  OR2X1 P2_sub_878_U149 ( .IN2(P2_sub_878_n152), .IN1(P2_sub_878_n151), 
        .Q(P2_sub_878_n150) );
  NAND2X0 P2_sub_878_U148 ( .IN1(P2_sub_878_n149), .IN2(P2_sub_878_n150), 
        .QN(P2_N2102) );
  INVX0 P2_sub_878_U147 ( .ZN(P2_sub_878_n135), .INP(P2_N1879) );
  NAND2X0 P2_sub_878_U146 ( .IN1(P2_N5091), .IN2(P2_sub_878_n135), 
        .QN(P2_sub_878_n147) );
  OR2X1 P2_sub_878_U145 ( .IN2(P2_N5091), .IN1(P2_sub_878_n135), 
        .Q(P2_sub_878_n148) );
  NAND2X0 P2_sub_878_U144 ( .IN1(P2_sub_878_n147), .IN2(P2_sub_878_n148), 
        .QN(P2_sub_878_n141) );
  NAND2X0 P2_sub_878_U143 ( .IN1(P2_N5090), .IN2(P2_sub_878_n146), 
        .QN(P2_sub_878_n142) );
  OR2X1 P2_sub_878_U142 ( .IN2(P2_N5090), .IN1(P2_sub_878_n146), 
        .Q(P2_sub_878_n144) );
  NAND2X0 P2_sub_878_U141 ( .IN1(P2_sub_878_n144), .IN2(P2_sub_878_n145), 
        .QN(P2_sub_878_n143) );
  NAND2X0 P2_sub_878_U140 ( .IN1(P2_sub_878_n142), .IN2(P2_sub_878_n143), 
        .QN(P2_sub_878_n136) );
  NAND2X0 P2_sub_878_U139 ( .IN1(P2_sub_878_n141), .IN2(P2_sub_878_n136), 
        .QN(P2_sub_878_n139) );
  OR2X1 P2_sub_878_U138 ( .IN2(P2_sub_878_n136), .IN1(P2_sub_878_n141), 
        .Q(P2_sub_878_n140) );
  NAND2X0 P2_sub_878_U137 ( .IN1(P2_sub_878_n139), .IN2(P2_sub_878_n140), 
        .QN(P2_N2121) );
  INVX0 P2_sub_878_U136 ( .ZN(P2_sub_878_n125), .INP(P2_N1880) );
  NAND2X0 P2_sub_878_U135 ( .IN1(n7252), .IN2(P2_sub_878_n125), 
        .QN(P2_sub_878_n137) );
  OR2X1 P2_sub_878_U134 ( .IN2(n7252), .IN1(P2_sub_878_n125), 
        .Q(P2_sub_878_n138) );
  NAND2X0 P2_sub_878_U133 ( .IN1(P2_sub_878_n137), .IN2(P2_sub_878_n138), 
        .QN(P2_sub_878_n131) );
  NAND2X0 P2_sub_878_U132 ( .IN1(P2_N5091), .IN2(P2_sub_878_n136), 
        .QN(P2_sub_878_n132) );
  OR2X1 P2_sub_878_U131 ( .IN2(P2_N5091), .IN1(P2_sub_878_n136), 
        .Q(P2_sub_878_n134) );
  NAND2X0 P2_sub_878_U130 ( .IN1(P2_sub_878_n134), .IN2(P2_sub_878_n135), 
        .QN(P2_sub_878_n133) );
  NAND2X0 P2_sub_878_U129 ( .IN1(P2_sub_878_n132), .IN2(P2_sub_878_n133), 
        .QN(P2_sub_878_n126) );
  NAND2X0 P2_sub_878_U128 ( .IN1(P2_sub_878_n131), .IN2(P2_sub_878_n126), 
        .QN(P2_sub_878_n129) );
  OR2X1 P2_sub_878_U127 ( .IN2(P2_sub_878_n126), .IN1(P2_sub_878_n131), 
        .Q(P2_sub_878_n130) );
  INVX0 P2_sub_878_U310 ( .ZN(P2_sub_878_n281), .INP(P2_N1859) );
  NOR2X0 P2_sub_878_U309 ( .QN(P2_sub_878_n277), .IN1(P2_sub_878_n281), 
        .IN2(n7035) );
  INVX0 P2_sub_878_U308 ( .ZN(P2_sub_878_n152), .INP(P2_sub_878_n277) );
  NAND2X0 P2_sub_878_U307 ( .IN1(n7035), .IN2(P2_sub_878_n281), 
        .QN(P2_sub_878_n280) );
  NAND2X0 P2_sub_878_U306 ( .IN1(P2_sub_878_n152), .IN2(P2_sub_878_n280), 
        .QN(P2_N2101) );
  INVX0 P2_sub_878_U305 ( .ZN(P2_sub_878_n243), .INP(P2_N1869) );
  NAND2X0 P2_sub_878_U304 ( .IN1(n7220), .IN2(P2_sub_878_n243), 
        .QN(P2_sub_878_n278) );
  OR2X1 P2_sub_878_U303 ( .IN2(n7220), .IN1(P2_sub_878_n243), 
        .Q(P2_sub_878_n279) );
  NAND2X0 P2_sub_878_U302 ( .IN1(P2_sub_878_n278), .IN2(P2_sub_878_n279), 
        .QN(P2_sub_878_n249) );
  NAND2X0 P2_sub_878_U301 ( .IN1(P2_N5072), .IN2(P2_sub_878_n152), 
        .QN(P2_sub_878_n274) );
  NAND2X0 P2_sub_878_U299 ( .IN1(P2_sub_878_n277), .IN2(n7186), 
        .QN(P2_sub_878_n276) );
  INVX0 P2_sub_878_U298 ( .ZN(P2_sub_878_n156), .INP(P2_N1860) );
  NAND2X0 P2_sub_878_U297 ( .IN1(P2_sub_878_n276), .IN2(P2_sub_878_n156), 
        .QN(P2_sub_878_n275) );
  NAND2X0 P2_sub_878_U296 ( .IN1(P2_sub_878_n274), .IN2(P2_sub_878_n275), 
        .QN(P2_sub_878_n53) );
  NAND2X0 P2_sub_878_U295 ( .IN1(n7181), .IN2(P2_sub_878_n53), 
        .QN(P2_sub_878_n271) );
  OR2X1 P2_sub_878_U294 ( .IN2(n7181), .IN1(P2_sub_878_n53), 
        .Q(P2_sub_878_n273) );
  INVX0 P2_sub_878_U293 ( .ZN(P2_sub_878_n56), .INP(P2_N1861) );
  NAND2X0 P2_sub_878_U292 ( .IN1(P2_sub_878_n273), .IN2(P2_sub_878_n56), 
        .QN(P2_sub_878_n272) );
  NAND2X0 P2_sub_878_U291 ( .IN1(P2_sub_878_n271), .IN2(P2_sub_878_n272), 
        .QN(P2_sub_878_n46) );
  NAND2X0 P2_sub_878_U290 ( .IN1(n7177), .IN2(P2_sub_878_n46), 
        .QN(P2_sub_878_n268) );
  OR2X1 P2_sub_878_U289 ( .IN2(n7177), .IN1(P2_sub_878_n46), 
        .Q(P2_sub_878_n270) );
  INVX0 P2_sub_878_U288 ( .ZN(P2_sub_878_n49), .INP(P2_N1862) );
  NAND2X0 P2_sub_878_U287 ( .IN1(P2_sub_878_n270), .IN2(P2_sub_878_n49), 
        .QN(P2_sub_878_n269) );
  NAND2X0 P2_sub_878_U286 ( .IN1(P2_sub_878_n268), .IN2(P2_sub_878_n269), 
        .QN(P2_sub_878_n39) );
  NAND2X0 P2_sub_878_U285 ( .IN1(n7173), .IN2(P2_sub_878_n39), 
        .QN(P2_sub_878_n265) );
  OR2X1 P2_sub_878_U284 ( .IN2(n7173), .IN1(P2_sub_878_n39), 
        .Q(P2_sub_878_n267) );
  INVX0 P2_sub_878_U283 ( .ZN(P2_sub_878_n42), .INP(P2_N1863) );
  NAND2X0 P2_sub_878_U282 ( .IN1(P2_sub_878_n267), .IN2(P2_sub_878_n42), 
        .QN(P2_sub_878_n266) );
  NAND2X0 P2_sub_878_U281 ( .IN1(P2_sub_878_n265), .IN2(P2_sub_878_n266), 
        .QN(P2_sub_878_n32) );
  NAND2X0 P2_sub_878_U280 ( .IN1(n7165), .IN2(P2_sub_878_n32), 
        .QN(P2_sub_878_n262) );
  OR2X1 P2_sub_878_U279 ( .IN2(n7165), .IN1(P2_sub_878_n32), 
        .Q(P2_sub_878_n264) );
  INVX0 P2_sub_878_U278 ( .ZN(P2_sub_878_n35), .INP(P2_N1864) );
  NAND2X0 P2_sub_878_U277 ( .IN1(P2_sub_878_n264), .IN2(P2_sub_878_n35), 
        .QN(P2_sub_878_n263) );
  NAND2X0 P2_sub_878_U276 ( .IN1(P2_sub_878_n262), .IN2(P2_sub_878_n263), 
        .QN(P2_sub_878_n25) );
  NAND2X0 P2_sub_878_U275 ( .IN1(P2_N5077), .IN2(P2_sub_878_n25), 
        .QN(P2_sub_878_n259) );
  OR2X1 P2_sub_878_U274 ( .IN2(P2_N5077), .IN1(P2_sub_878_n25), 
        .Q(P2_sub_878_n261) );
  INVX0 P2_sub_878_U273 ( .ZN(P2_sub_878_n28), .INP(P2_N1865) );
  NAND2X0 P2_sub_878_U272 ( .IN1(P2_sub_878_n261), .IN2(P2_sub_878_n28), 
        .QN(P2_sub_878_n260) );
  NAND2X0 P2_sub_878_U271 ( .IN1(P2_sub_878_n259), .IN2(P2_sub_878_n260), 
        .QN(P2_sub_878_n18) );
  NAND2X0 P2_sub_878_U270 ( .IN1(P2_N5078), .IN2(P2_sub_878_n18), 
        .QN(P2_sub_878_n256) );
  OR2X1 P2_sub_878_U269 ( .IN2(P2_N5078), .IN1(P2_sub_878_n18), 
        .Q(P2_sub_878_n258) );
  INVX0 P2_sub_878_U268 ( .ZN(P2_sub_878_n21), .INP(P2_N1866) );
  NAND2X0 P2_sub_878_U267 ( .IN1(P2_sub_878_n258), .IN2(P2_sub_878_n21), 
        .QN(P2_sub_878_n257) );
  NAND2X0 P2_sub_878_U266 ( .IN1(P2_sub_878_n256), .IN2(P2_sub_878_n257), 
        .QN(P2_sub_878_n11) );
  NAND2X0 P2_sub_878_U265 ( .IN1(P2_N5079), .IN2(P2_sub_878_n11), 
        .QN(P2_sub_878_n253) );
  OR2X1 P2_sub_878_U264 ( .IN2(P2_N5079), .IN1(P2_sub_878_n11), 
        .Q(P2_sub_878_n255) );
  INVX0 P2_sub_878_U263 ( .ZN(P2_sub_878_n14), .INP(P2_N1867) );
  NAND2X0 P2_sub_878_U262 ( .IN1(P2_sub_878_n255), .IN2(P2_sub_878_n14), 
        .QN(P2_sub_878_n254) );
  NAND2X0 P2_sub_878_U261 ( .IN1(P2_sub_878_n253), .IN2(P2_sub_878_n254), 
        .QN(P2_sub_878_n4) );
  NAND2X0 P2_sub_878_U260 ( .IN1(n7151), .IN2(P2_sub_878_n4), 
        .QN(P2_sub_878_n250) );
  OR2X1 P2_sub_878_U259 ( .IN2(n7151), .IN1(P2_sub_878_n4), 
        .Q(P2_sub_878_n252) );
  INVX0 P2_sub_878_U258 ( .ZN(P2_sub_878_n7), .INP(P2_N1868) );
  NAND2X0 P2_sub_878_U257 ( .IN1(P2_sub_878_n252), .IN2(P2_sub_878_n7), 
        .QN(P2_sub_878_n251) );
  NAND2X0 P2_sub_878_U256 ( .IN1(P2_sub_878_n250), .IN2(P2_sub_878_n251), 
        .QN(P2_sub_878_n244) );
  NAND2X0 P2_sub_878_U255 ( .IN1(P2_sub_878_n249), .IN2(P2_sub_878_n244), 
        .QN(P2_sub_878_n247) );
  OR2X1 P2_sub_878_U254 ( .IN2(P2_sub_878_n244), .IN1(P2_sub_878_n249), 
        .Q(P2_sub_878_n248) );
  NAND2X0 P2_sub_878_U253 ( .IN1(P2_sub_878_n247), .IN2(P2_sub_878_n248), 
        .QN(P2_N2111) );
  INVX0 P2_sub_878_U252 ( .ZN(P2_sub_878_n233), .INP(P2_N1870) );
  NAND2X0 P2_sub_878_U251 ( .IN1(P2_N5082), .IN2(P2_sub_878_n233), 
        .QN(P2_sub_878_n245) );
  OR2X1 P2_sub_878_U250 ( .IN2(P2_N5082), .IN1(P2_sub_878_n233), 
        .Q(P2_sub_878_n246) );
  NAND2X0 P2_sub_878_U249 ( .IN1(P2_sub_878_n245), .IN2(P2_sub_878_n246), 
        .QN(P2_sub_878_n239) );
  NAND2X0 P2_sub_878_U248 ( .IN1(n7220), .IN2(P2_sub_878_n244), 
        .QN(P2_sub_878_n240) );
  OR2X1 P2_sub_878_U247 ( .IN2(n7220), .IN1(P2_sub_878_n244), 
        .Q(P2_sub_878_n242) );
  NAND2X0 P2_sub_878_U246 ( .IN1(P2_sub_878_n242), .IN2(P2_sub_878_n243), 
        .QN(P2_sub_878_n241) );
  NAND2X0 P2_sub_878_U245 ( .IN1(P2_sub_878_n240), .IN2(P2_sub_878_n241), 
        .QN(P2_sub_878_n234) );
  NAND2X0 P2_sub_878_U244 ( .IN1(P2_sub_878_n239), .IN2(P2_sub_878_n234), 
        .QN(P2_sub_878_n237) );
  OR2X1 P2_sub_878_U243 ( .IN2(P2_sub_878_n234), .IN1(P2_sub_878_n239), 
        .Q(P2_sub_878_n238) );
  NAND2X0 P2_sub_878_U242 ( .IN1(P2_sub_878_n237), .IN2(P2_sub_878_n238), 
        .QN(P2_N2112) );
  INVX0 P2_sub_878_U241 ( .ZN(P2_sub_878_n223), .INP(P2_N1871) );
  NAND2X0 P2_sub_878_U240 ( .IN1(P2_N5083), .IN2(P2_sub_878_n223), 
        .QN(P2_sub_878_n235) );
  OR2X1 P2_sub_878_U239 ( .IN2(P2_N5083), .IN1(P2_sub_878_n223), 
        .Q(P2_sub_878_n236) );
  NAND2X0 P2_sub_878_U238 ( .IN1(P2_sub_878_n235), .IN2(P2_sub_878_n236), 
        .QN(P2_sub_878_n229) );
  NAND2X0 P2_sub_878_U237 ( .IN1(P2_N5082), .IN2(P2_sub_878_n234), 
        .QN(P2_sub_878_n230) );
  OR2X1 P2_sub_878_U236 ( .IN2(P2_N5082), .IN1(P2_sub_878_n234), 
        .Q(P2_sub_878_n232) );
  NAND2X0 P2_sub_878_U235 ( .IN1(P2_sub_878_n232), .IN2(P2_sub_878_n233), 
        .QN(P2_sub_878_n231) );
  NAND2X0 P2_sub_878_U234 ( .IN1(P2_sub_878_n230), .IN2(P2_sub_878_n231), 
        .QN(P2_sub_878_n224) );
  NAND2X0 P2_sub_878_U233 ( .IN1(P2_sub_878_n229), .IN2(P2_sub_878_n224), 
        .QN(P2_sub_878_n227) );
  OR2X1 P2_sub_878_U232 ( .IN2(P2_sub_878_n224), .IN1(P2_sub_878_n229), 
        .Q(P2_sub_878_n228) );
  NAND2X0 P2_sub_878_U231 ( .IN1(P2_sub_878_n227), .IN2(P2_sub_878_n228), 
        .QN(P2_N2113) );
  INVX0 P2_sub_878_U230 ( .ZN(P2_sub_878_n213), .INP(P2_N1872) );
  NAND2X0 P2_sub_878_U229 ( .IN1(P2_N5084), .IN2(P2_sub_878_n213), 
        .QN(P2_sub_878_n225) );
  OR2X1 P2_sub_878_U228 ( .IN2(P2_N5084), .IN1(P2_sub_878_n213), 
        .Q(P2_sub_878_n226) );
  NAND2X0 P2_sub_878_U227 ( .IN1(P2_sub_878_n225), .IN2(P2_sub_878_n226), 
        .QN(P2_sub_878_n219) );
  NAND2X0 P2_sub_878_U226 ( .IN1(P2_N5083), .IN2(P2_sub_878_n224), 
        .QN(P2_sub_878_n220) );
  OR2X1 P2_sub_878_U225 ( .IN2(P2_N5083), .IN1(P2_sub_878_n224), 
        .Q(P2_sub_878_n222) );
  NAND2X0 P2_sub_878_U224 ( .IN1(P2_sub_878_n222), .IN2(P2_sub_878_n223), 
        .QN(P2_sub_878_n221) );
  NAND2X0 P2_sub_878_U223 ( .IN1(P2_sub_878_n220), .IN2(P2_sub_878_n221), 
        .QN(P2_sub_878_n214) );
  NAND2X0 P2_sub_878_U222 ( .IN1(P2_sub_878_n219), .IN2(P2_sub_878_n214), 
        .QN(P2_sub_878_n217) );
  OR2X1 P2_sub_878_U221 ( .IN2(P2_sub_878_n214), .IN1(P2_sub_878_n219), 
        .Q(P2_sub_878_n218) );
  NAND2X0 P2_sub_878_U220 ( .IN1(P2_sub_878_n217), .IN2(P2_sub_878_n218), 
        .QN(P2_N2114) );
  NAND2X0 P2_add_898_U63 ( .IN1(P2_N5098), .IN2(P2_add_898_n64), 
        .QN(P2_add_898_n61) );
  OR2X1 P2_add_898_U62 ( .IN2(P2_N5098), .IN1(P2_add_898_n64), 
        .Q(P2_add_898_n63) );
  NAND2X0 P2_add_898_U61 ( .IN1(P2_N2259), .IN2(P2_add_898_n63), 
        .QN(P2_add_898_n62) );
  NAND2X0 P2_add_898_U60 ( .IN1(P2_add_898_n61), .IN2(P2_add_898_n62), 
        .QN(P2_add_898_n59) );
  NOR2X0 P2_add_898_U59 ( .QN(P2_add_898_n57), .IN1(P2_add_898_n60), 
        .IN2(P2_add_898_n59) );
  AND2X1 P2_add_898_U58 ( .IN1(P2_add_898_n59), .IN2(P2_add_898_n60), 
        .Q(P2_add_898_n58) );
  NOR2X0 P2_add_898_U57 ( .QN(P2_N2502), .IN1(P2_add_898_n57), 
        .IN2(P2_add_898_n58) );
  OR2X1 P2_add_898_U55 ( .IN2(P2_N2234), .IN1(n7182), .Q(P2_add_898_n54) );
  NAND2X0 P2_add_898_U54 ( .IN1(P2_N2234), .IN2(n7182), .QN(P2_add_898_n55) );
  NAND2X0 P2_add_898_U53 ( .IN1(P2_add_898_n54), .IN2(P2_add_898_n55), 
        .QN(P2_add_898_n53) );
  NOR2X0 P2_add_898_U52 ( .QN(P2_add_898_n50), .IN1(P2_add_898_n52), 
        .IN2(P2_add_898_n53) );
  AND2X1 P2_add_898_U51 ( .IN1(P2_add_898_n52), .IN2(P2_add_898_n53), 
        .Q(P2_add_898_n51) );
  NOR2X0 P2_add_898_U50 ( .QN(P2_N2476), .IN1(P2_add_898_n50), 
        .IN2(P2_add_898_n51) );
  OR2X1 P2_add_898_U48 ( .IN2(P2_N2235), .IN1(n7178), .Q(P2_add_898_n47) );
  NAND2X0 P2_add_898_U47 ( .IN1(P2_N2235), .IN2(n7178), .QN(P2_add_898_n48) );
  NAND2X0 P2_add_898_U46 ( .IN1(P2_add_898_n47), .IN2(P2_add_898_n48), 
        .QN(P2_add_898_n46) );
  NOR2X0 P2_add_898_U45 ( .QN(P2_add_898_n43), .IN1(P2_add_898_n45), 
        .IN2(P2_add_898_n46) );
  AND2X1 P2_add_898_U44 ( .IN1(P2_add_898_n45), .IN2(P2_add_898_n46), 
        .Q(P2_add_898_n44) );
  NOR2X0 P2_add_898_U43 ( .QN(P2_N2477), .IN1(P2_add_898_n43), 
        .IN2(P2_add_898_n44) );
  OR2X1 P2_add_898_U41 ( .IN2(P2_N2236), .IN1(n7174), .Q(P2_add_898_n40) );
  NAND2X0 P2_add_898_U40 ( .IN1(P2_N2236), .IN2(n7174), .QN(P2_add_898_n41) );
  NAND2X0 P2_add_898_U39 ( .IN1(P2_add_898_n40), .IN2(P2_add_898_n41), 
        .QN(P2_add_898_n39) );
  NOR2X0 P2_add_898_U38 ( .QN(P2_add_898_n36), .IN1(P2_add_898_n38), 
        .IN2(P2_add_898_n39) );
  AND2X1 P2_add_898_U37 ( .IN1(P2_add_898_n38), .IN2(P2_add_898_n39), 
        .Q(P2_add_898_n37) );
  NOR2X0 P2_add_898_U36 ( .QN(P2_N2478), .IN1(P2_add_898_n36), 
        .IN2(P2_add_898_n37) );
  OR2X1 P2_add_898_U34 ( .IN2(P2_N2237), .IN1(n7166), .Q(P2_add_898_n33) );
  NAND2X0 P2_add_898_U33 ( .IN1(P2_N2237), .IN2(n7166), .QN(P2_add_898_n34) );
  NAND2X0 P2_add_898_U32 ( .IN1(P2_add_898_n33), .IN2(P2_add_898_n34), 
        .QN(P2_add_898_n32) );
  NOR2X0 P2_add_898_U31 ( .QN(P2_add_898_n29), .IN1(P2_add_898_n31), 
        .IN2(P2_add_898_n32) );
  AND2X1 P2_add_898_U30 ( .IN1(P2_add_898_n31), .IN2(P2_add_898_n32), 
        .Q(P2_add_898_n30) );
  NOR2X0 P2_add_898_U29 ( .QN(P2_N2479), .IN1(P2_add_898_n29), 
        .IN2(P2_add_898_n30) );
  OR2X1 P2_add_898_U27 ( .IN2(P2_N2238), .IN1(n7164), .Q(P2_add_898_n26) );
  NAND2X0 P2_add_898_U26 ( .IN1(P2_N2238), .IN2(n7164), .QN(P2_add_898_n27) );
  NAND2X0 P2_add_898_U25 ( .IN1(P2_add_898_n26), .IN2(P2_add_898_n27), 
        .QN(P2_add_898_n25) );
  NOR2X0 P2_add_898_U24 ( .QN(P2_add_898_n22), .IN1(P2_add_898_n24), 
        .IN2(P2_add_898_n25) );
  AND2X1 P2_add_898_U23 ( .IN1(P2_add_898_n24), .IN2(P2_add_898_n25), 
        .Q(P2_add_898_n23) );
  NOR2X0 P2_add_898_U22 ( .QN(P2_N2480), .IN1(P2_add_898_n22), 
        .IN2(P2_add_898_n23) );
  OR2X1 P2_add_898_U20 ( .IN2(P2_N2239), .IN1(n7157), .Q(P2_add_898_n19) );
  NAND2X0 P2_add_898_U19 ( .IN1(P2_N2239), .IN2(n7157), .QN(P2_add_898_n20) );
  NAND2X0 P2_add_898_U18 ( .IN1(P2_add_898_n19), .IN2(P2_add_898_n20), 
        .QN(P2_add_898_n18) );
  NOR2X0 P2_add_898_U17 ( .QN(P2_add_898_n15), .IN1(P2_add_898_n17), 
        .IN2(P2_add_898_n18) );
  AND2X1 P2_add_898_U16 ( .IN1(P2_add_898_n17), .IN2(P2_add_898_n18), 
        .Q(P2_add_898_n16) );
  NOR2X0 P2_add_898_U15 ( .QN(P2_N2481), .IN1(P2_add_898_n15), 
        .IN2(P2_add_898_n16) );
  OR2X1 P2_add_898_U13 ( .IN2(P2_N2240), .IN1(n7153), .Q(P2_add_898_n12) );
  NAND2X0 P2_add_898_U12 ( .IN1(P2_N2240), .IN2(n7153), .QN(P2_add_898_n13) );
  NAND2X0 P2_add_898_U11 ( .IN1(P2_add_898_n12), .IN2(P2_add_898_n13), 
        .QN(P2_add_898_n11) );
  NOR2X0 P2_add_898_U10 ( .QN(P2_add_898_n8), .IN1(P2_add_898_n10), 
        .IN2(P2_add_898_n11) );
  AND2X1 P2_add_898_U9 ( .IN1(P2_add_898_n10), .IN2(P2_add_898_n11), 
        .Q(P2_add_898_n9) );
  NOR2X0 P2_add_898_U8 ( .QN(P2_N2482), .IN1(P2_add_898_n8), 
        .IN2(P2_add_898_n9) );
  OR2X1 P2_add_898_U6 ( .IN2(P2_N2241), .IN1(n7149), .Q(P2_add_898_n5) );
  NAND2X0 P2_add_898_U5 ( .IN1(P2_N2241), .IN2(n7149), .QN(P2_add_898_n6) );
  NAND2X0 P2_add_898_U4 ( .IN1(P2_add_898_n5), .IN2(P2_add_898_n6), 
        .QN(P2_add_898_n4) );
  NOR2X0 P2_add_898_U3 ( .QN(P2_add_898_n1), .IN1(P2_add_898_n3), 
        .IN2(P2_add_898_n4) );
  AND2X1 P2_add_898_U2 ( .IN1(P2_add_898_n3), .IN2(P2_add_898_n4), 
        .Q(P2_add_898_n2) );
  NOR2X0 P2_add_898_U1 ( .QN(P2_N2483), .IN1(P2_add_898_n1), 
        .IN2(P2_add_898_n2) );
  NAND2X0 P2_add_898_U156 ( .IN1(P2_add_898_n148), .IN2(P2_add_898_n149), 
        .QN(P2_N2475) );
  NAND2X0 P2_add_898_U155 ( .IN1(P2_N5090), .IN2(P2_add_898_n147), 
        .QN(P2_add_898_n144) );
  OR2X1 P2_add_898_U154 ( .IN2(P2_N5090), .IN1(P2_add_898_n147), 
        .Q(P2_add_898_n146) );
  NAND2X0 P2_add_898_U153 ( .IN1(P2_N2251), .IN2(P2_add_898_n146), 
        .QN(P2_add_898_n145) );
  NAND2X0 P2_add_898_U152 ( .IN1(P2_add_898_n144), .IN2(P2_add_898_n145), 
        .QN(P2_add_898_n137) );
  OR2X1 P2_add_898_U150 ( .IN2(P2_N2252), .IN1(n7260), .Q(P2_add_898_n141) );
  NAND2X0 P2_add_898_U149 ( .IN1(P2_N2252), .IN2(n7260), .QN(P2_add_898_n142)
         );
  NAND2X0 P2_add_898_U148 ( .IN1(P2_add_898_n141), .IN2(P2_add_898_n142), 
        .QN(P2_add_898_n140) );
  NOR2X0 P2_add_898_U147 ( .QN(P2_add_898_n138), .IN1(P2_add_898_n137), 
        .IN2(P2_add_898_n140) );
  AND2X1 P2_add_898_U146 ( .IN1(P2_add_898_n137), .IN2(P2_add_898_n140), 
        .Q(P2_add_898_n139) );
  NOR2X0 P2_add_898_U145 ( .QN(P2_N2494), .IN1(P2_add_898_n138), 
        .IN2(P2_add_898_n139) );
  NAND2X0 P2_add_898_U144 ( .IN1(P2_N5091), .IN2(P2_add_898_n137), 
        .QN(P2_add_898_n134) );
  OR2X1 P2_add_898_U143 ( .IN2(P2_N5091), .IN1(P2_add_898_n137), 
        .Q(P2_add_898_n136) );
  NAND2X0 P2_add_898_U142 ( .IN1(P2_N2252), .IN2(P2_add_898_n136), 
        .QN(P2_add_898_n135) );
  NAND2X0 P2_add_898_U141 ( .IN1(P2_add_898_n134), .IN2(P2_add_898_n135), 
        .QN(P2_add_898_n127) );
  OR2X1 P2_add_898_U139 ( .IN2(P2_N2253), .IN1(n7253), .Q(P2_add_898_n131) );
  NAND2X0 P2_add_898_U138 ( .IN1(P2_N2253), .IN2(n7253), .QN(P2_add_898_n132)
         );
  NAND2X0 P2_add_898_U137 ( .IN1(P2_add_898_n131), .IN2(P2_add_898_n132), 
        .QN(P2_add_898_n130) );
  NOR2X0 P2_add_898_U136 ( .QN(P2_add_898_n128), .IN1(P2_add_898_n127), 
        .IN2(P2_add_898_n130) );
  AND2X1 P2_add_898_U135 ( .IN1(P2_add_898_n127), .IN2(P2_add_898_n130), 
        .Q(P2_add_898_n129) );
  NOR2X0 P2_add_898_U134 ( .QN(P2_N2495), .IN1(P2_add_898_n128), 
        .IN2(P2_add_898_n129) );
  NAND2X0 P2_add_898_U133 ( .IN1(P2_N5092), .IN2(P2_add_898_n127), 
        .QN(P2_add_898_n124) );
  OR2X1 P2_add_898_U132 ( .IN2(P2_N5092), .IN1(P2_add_898_n127), 
        .Q(P2_add_898_n126) );
  NAND2X0 P2_add_898_U131 ( .IN1(P2_N2253), .IN2(P2_add_898_n126), 
        .QN(P2_add_898_n125) );
  NAND2X0 P2_add_898_U130 ( .IN1(P2_add_898_n124), .IN2(P2_add_898_n125), 
        .QN(P2_add_898_n117) );
  OR2X1 P2_add_898_U128 ( .IN2(P2_N2254), .IN1(n7248), .Q(P2_add_898_n121) );
  NAND2X0 P2_add_898_U127 ( .IN1(P2_N2254), .IN2(n7248), .QN(P2_add_898_n122)
         );
  NAND2X0 P2_add_898_U126 ( .IN1(P2_add_898_n121), .IN2(P2_add_898_n122), 
        .QN(P2_add_898_n120) );
  NOR2X0 P2_add_898_U125 ( .QN(P2_add_898_n118), .IN1(P2_add_898_n117), 
        .IN2(P2_add_898_n120) );
  AND2X1 P2_add_898_U124 ( .IN1(P2_add_898_n117), .IN2(P2_add_898_n120), 
        .Q(P2_add_898_n119) );
  NOR2X0 P2_add_898_U123 ( .QN(P2_N2496), .IN1(P2_add_898_n118), 
        .IN2(P2_add_898_n119) );
  NAND2X0 P2_add_898_U122 ( .IN1(n7247), .IN2(P2_add_898_n117), 
        .QN(P2_add_898_n114) );
  OR2X1 P2_add_898_U121 ( .IN2(n7247), .IN1(P2_add_898_n117), 
        .Q(P2_add_898_n116) );
  NAND2X0 P2_add_898_U120 ( .IN1(P2_N2254), .IN2(P2_add_898_n116), 
        .QN(P2_add_898_n115) );
  NAND2X0 P2_add_898_U119 ( .IN1(P2_add_898_n114), .IN2(P2_add_898_n115), 
        .QN(P2_add_898_n107) );
  OR2X1 P2_add_898_U117 ( .IN2(P2_N2255), .IN1(P2_add_898_n299), 
        .Q(P2_add_898_n111) );
  NAND2X0 P2_add_898_U116 ( .IN1(P2_N2255), .IN2(n7243), .QN(P2_add_898_n112)
         );
  NAND2X0 P2_add_898_U115 ( .IN1(P2_add_898_n111), .IN2(P2_add_898_n112), 
        .QN(P2_add_898_n110) );
  NOR2X0 P2_add_898_U114 ( .QN(P2_add_898_n108), .IN1(P2_add_898_n107), 
        .IN2(P2_add_898_n110) );
  AND2X1 P2_add_898_U113 ( .IN1(P2_add_898_n107), .IN2(P2_add_898_n110), 
        .Q(P2_add_898_n109) );
  NOR2X0 P2_add_898_U112 ( .QN(P2_N2497), .IN1(P2_add_898_n108), 
        .IN2(P2_add_898_n109) );
  NAND2X0 P2_add_898_U111 ( .IN1(P2_N5094), .IN2(P2_add_898_n107), 
        .QN(P2_add_898_n104) );
  OR2X1 P2_add_898_U110 ( .IN2(P2_N5094), .IN1(P2_add_898_n107), 
        .Q(P2_add_898_n106) );
  NAND2X0 P2_add_898_U109 ( .IN1(P2_N2255), .IN2(P2_add_898_n106), 
        .QN(P2_add_898_n105) );
  NAND2X0 P2_add_898_U108 ( .IN1(P2_add_898_n104), .IN2(P2_add_898_n105), 
        .QN(P2_add_898_n97) );
  OR2X1 P2_add_898_U106 ( .IN2(P2_N2256), .IN1(n7239), .Q(P2_add_898_n101) );
  NAND2X0 P2_add_898_U105 ( .IN1(P2_N2256), .IN2(n7239), .QN(P2_add_898_n102)
         );
  NAND2X0 P2_add_898_U104 ( .IN1(P2_add_898_n101), .IN2(P2_add_898_n102), 
        .QN(P2_add_898_n100) );
  NOR2X0 P2_add_898_U103 ( .QN(P2_add_898_n98), .IN1(P2_add_898_n97), 
        .IN2(P2_add_898_n100) );
  AND2X1 P2_add_898_U102 ( .IN1(P2_add_898_n97), .IN2(P2_add_898_n100), 
        .Q(P2_add_898_n99) );
  NOR2X0 P2_add_898_U101 ( .QN(P2_N2498), .IN1(P2_add_898_n98), 
        .IN2(P2_add_898_n99) );
  NAND2X0 P2_add_898_U100 ( .IN1(n7238), .IN2(P2_add_898_n97), 
        .QN(P2_add_898_n94) );
  OR2X1 P2_add_898_U99 ( .IN2(n7238), .IN1(P2_add_898_n97), .Q(P2_add_898_n96)
         );
  NAND2X0 P2_add_898_U98 ( .IN1(P2_N2256), .IN2(P2_add_898_n96), 
        .QN(P2_add_898_n95) );
  NAND2X0 P2_add_898_U97 ( .IN1(P2_add_898_n94), .IN2(P2_add_898_n95), 
        .QN(P2_add_898_n87) );
  OR2X1 P2_add_898_U95 ( .IN2(P2_N2257), .IN1(n7234), .Q(P2_add_898_n91) );
  NAND2X0 P2_add_898_U94 ( .IN1(P2_N2257), .IN2(n7234), .QN(P2_add_898_n92) );
  NAND2X0 P2_add_898_U93 ( .IN1(P2_add_898_n91), .IN2(P2_add_898_n92), 
        .QN(P2_add_898_n90) );
  NOR2X0 P2_add_898_U92 ( .QN(P2_add_898_n88), .IN1(P2_add_898_n87), 
        .IN2(P2_add_898_n90) );
  AND2X1 P2_add_898_U91 ( .IN1(P2_add_898_n87), .IN2(P2_add_898_n90), 
        .Q(P2_add_898_n89) );
  NOR2X0 P2_add_898_U90 ( .QN(P2_N2499), .IN1(P2_add_898_n88), 
        .IN2(P2_add_898_n89) );
  NAND2X0 P2_add_898_U89 ( .IN1(P2_N5096), .IN2(P2_add_898_n87), 
        .QN(P2_add_898_n84) );
  OR2X1 P2_add_898_U88 ( .IN2(P2_N5096), .IN1(P2_add_898_n87), 
        .Q(P2_add_898_n86) );
  NAND2X0 P2_add_898_U87 ( .IN1(P2_N2257), .IN2(P2_add_898_n86), 
        .QN(P2_add_898_n85) );
  NAND2X0 P2_add_898_U86 ( .IN1(P2_add_898_n84), .IN2(P2_add_898_n85), 
        .QN(P2_add_898_n77) );
  OR2X1 P2_add_898_U84 ( .IN2(P2_N2258), .IN1(n7229), .Q(P2_add_898_n81) );
  NAND2X0 P2_add_898_U83 ( .IN1(P2_N2258), .IN2(n7229), .QN(P2_add_898_n82) );
  NAND2X0 P2_add_898_U82 ( .IN1(P2_add_898_n81), .IN2(P2_add_898_n82), 
        .QN(P2_add_898_n80) );
  NOR2X0 P2_add_898_U81 ( .QN(P2_add_898_n78), .IN1(P2_add_898_n77), 
        .IN2(P2_add_898_n80) );
  AND2X1 P2_add_898_U80 ( .IN1(P2_add_898_n77), .IN2(P2_add_898_n80), 
        .Q(P2_add_898_n79) );
  NOR2X0 P2_add_898_U79 ( .QN(P2_N2500), .IN1(P2_add_898_n78), 
        .IN2(P2_add_898_n79) );
  NAND2X0 P2_add_898_U78 ( .IN1(P2_N5097), .IN2(P2_add_898_n77), 
        .QN(P2_add_898_n74) );
  OR2X1 P2_add_898_U77 ( .IN2(P2_N5097), .IN1(P2_add_898_n77), 
        .Q(P2_add_898_n76) );
  NAND2X0 P2_add_898_U76 ( .IN1(P2_N2258), .IN2(P2_add_898_n76), 
        .QN(P2_add_898_n75) );
  NAND2X0 P2_add_898_U75 ( .IN1(P2_add_898_n74), .IN2(P2_add_898_n75), 
        .QN(P2_add_898_n64) );
  OR2X1 P2_add_898_U73 ( .IN2(P2_N2259), .IN1(n7224), .Q(P2_add_898_n71) );
  NAND2X0 P2_add_898_U72 ( .IN1(P2_N2259), .IN2(n7224), .QN(P2_add_898_n72) );
  NAND2X0 P2_add_898_U71 ( .IN1(P2_add_898_n71), .IN2(P2_add_898_n72), 
        .QN(P2_add_898_n70) );
  NOR2X0 P2_add_898_U70 ( .QN(P2_add_898_n68), .IN1(P2_add_898_n64), 
        .IN2(P2_add_898_n70) );
  AND2X1 P2_add_898_U69 ( .IN1(P2_add_898_n64), .IN2(P2_add_898_n70), 
        .Q(P2_add_898_n69) );
  NOR2X0 P2_add_898_U68 ( .QN(P2_N2501), .IN1(P2_add_898_n68), 
        .IN2(P2_add_898_n69) );
  OR2X1 P2_add_898_U66 ( .IN2(P2_N2260), .IN1(n7222), .Q(P2_add_898_n65) );
  NAND2X0 P2_add_898_U65 ( .IN1(P2_N2260), .IN2(n7222), .QN(P2_add_898_n66) );
  NAND2X0 P2_add_898_U64 ( .IN1(P2_add_898_n65), .IN2(P2_add_898_n66), 
        .QN(P2_add_898_n60) );
  NAND2X0 P2_add_898_U249 ( .IN1(n7216), .IN2(P2_add_898_n234), 
        .QN(P2_add_898_n231) );
  OR2X1 P2_add_898_U248 ( .IN2(n7216), .IN1(P2_add_898_n234), 
        .Q(P2_add_898_n233) );
  NAND2X0 P2_add_898_U247 ( .IN1(P2_N2243), .IN2(P2_add_898_n233), 
        .QN(P2_add_898_n232) );
  NAND2X0 P2_add_898_U246 ( .IN1(P2_add_898_n231), .IN2(P2_add_898_n232), 
        .QN(P2_add_898_n224) );
  OR2X1 P2_add_898_U244 ( .IN2(P2_N2244), .IN1(n7211), .Q(P2_add_898_n228) );
  NAND2X0 P2_add_898_U243 ( .IN1(P2_N2244), .IN2(n7211), .QN(P2_add_898_n229)
         );
  NAND2X0 P2_add_898_U242 ( .IN1(P2_add_898_n228), .IN2(P2_add_898_n229), 
        .QN(P2_add_898_n227) );
  NOR2X0 P2_add_898_U241 ( .QN(P2_add_898_n225), .IN1(P2_add_898_n224), 
        .IN2(P2_add_898_n227) );
  AND2X1 P2_add_898_U240 ( .IN1(P2_add_898_n224), .IN2(P2_add_898_n227), 
        .Q(P2_add_898_n226) );
  NOR2X0 P2_add_898_U239 ( .QN(P2_N2486), .IN1(P2_add_898_n225), 
        .IN2(P2_add_898_n226) );
  NAND2X0 P2_add_898_U238 ( .IN1(n7210), .IN2(P2_add_898_n224), 
        .QN(P2_add_898_n221) );
  OR2X1 P2_add_898_U237 ( .IN2(n7210), .IN1(P2_add_898_n224), 
        .Q(P2_add_898_n223) );
  NAND2X0 P2_add_898_U236 ( .IN1(P2_N2244), .IN2(P2_add_898_n223), 
        .QN(P2_add_898_n222) );
  NAND2X0 P2_add_898_U235 ( .IN1(P2_add_898_n221), .IN2(P2_add_898_n222), 
        .QN(P2_add_898_n214) );
  OR2X1 P2_add_898_U233 ( .IN2(P2_N2245), .IN1(n7208), .Q(P2_add_898_n218) );
  NAND2X0 P2_add_898_U232 ( .IN1(P2_N2245), .IN2(n7208), .QN(P2_add_898_n219)
         );
  NAND2X0 P2_add_898_U231 ( .IN1(P2_add_898_n218), .IN2(P2_add_898_n219), 
        .QN(P2_add_898_n217) );
  NOR2X0 P2_add_898_U230 ( .QN(P2_add_898_n215), .IN1(P2_add_898_n214), 
        .IN2(P2_add_898_n217) );
  AND2X1 P2_add_898_U229 ( .IN1(P2_add_898_n214), .IN2(P2_add_898_n217), 
        .Q(P2_add_898_n216) );
  NOR2X0 P2_add_898_U228 ( .QN(P2_N2487), .IN1(P2_add_898_n215), 
        .IN2(P2_add_898_n216) );
  NAND2X0 P2_add_898_U227 ( .IN1(n7209), .IN2(P2_add_898_n214), 
        .QN(P2_add_898_n211) );
  OR2X1 P2_add_898_U226 ( .IN2(n7209), .IN1(P2_add_898_n214), 
        .Q(P2_add_898_n213) );
  NAND2X0 P2_add_898_U225 ( .IN1(P2_N2245), .IN2(P2_add_898_n213), 
        .QN(P2_add_898_n212) );
  NAND2X0 P2_add_898_U224 ( .IN1(P2_add_898_n211), .IN2(P2_add_898_n212), 
        .QN(P2_add_898_n204) );
  OR2X1 P2_add_898_U222 ( .IN2(P2_N2246), .IN1(n7205), .Q(P2_add_898_n208) );
  NAND2X0 P2_add_898_U221 ( .IN1(P2_N2246), .IN2(n7205), .QN(P2_add_898_n209)
         );
  NAND2X0 P2_add_898_U220 ( .IN1(P2_add_898_n208), .IN2(P2_add_898_n209), 
        .QN(P2_add_898_n207) );
  NOR2X0 P2_add_898_U219 ( .QN(P2_add_898_n205), .IN1(P2_add_898_n204), 
        .IN2(P2_add_898_n207) );
  AND2X1 P2_add_898_U218 ( .IN1(P2_add_898_n204), .IN2(P2_add_898_n207), 
        .Q(P2_add_898_n206) );
  NOR2X0 P2_add_898_U217 ( .QN(P2_N2488), .IN1(P2_add_898_n205), 
        .IN2(P2_add_898_n206) );
  NAND2X0 P2_add_898_U216 ( .IN1(n7206), .IN2(P2_add_898_n204), 
        .QN(P2_add_898_n201) );
  OR2X1 P2_add_898_U215 ( .IN2(n7206), .IN1(P2_add_898_n204), 
        .Q(P2_add_898_n203) );
  NAND2X0 P2_add_898_U214 ( .IN1(P2_N2246), .IN2(P2_add_898_n203), 
        .QN(P2_add_898_n202) );
  NAND2X0 P2_add_898_U213 ( .IN1(P2_add_898_n201), .IN2(P2_add_898_n202), 
        .QN(P2_add_898_n194) );
  OR2X1 P2_add_898_U211 ( .IN2(P2_N2247), .IN1(n7201), .Q(P2_add_898_n198) );
  NAND2X0 P2_add_898_U210 ( .IN1(P2_N2247), .IN2(n7201), .QN(P2_add_898_n199)
         );
  NAND2X0 P2_add_898_U209 ( .IN1(P2_add_898_n198), .IN2(P2_add_898_n199), 
        .QN(P2_add_898_n197) );
  NOR2X0 P2_add_898_U208 ( .QN(P2_add_898_n195), .IN1(P2_add_898_n194), 
        .IN2(P2_add_898_n197) );
  AND2X1 P2_add_898_U207 ( .IN1(P2_add_898_n194), .IN2(P2_add_898_n197), 
        .Q(P2_add_898_n196) );
  NOR2X0 P2_add_898_U206 ( .QN(P2_N2489), .IN1(P2_add_898_n195), 
        .IN2(P2_add_898_n196) );
  NAND2X0 P2_add_898_U205 ( .IN1(P2_N5086), .IN2(P2_add_898_n194), 
        .QN(P2_add_898_n191) );
  OR2X1 P2_add_898_U204 ( .IN2(P2_N5086), .IN1(P2_add_898_n194), 
        .Q(P2_add_898_n193) );
  NAND2X0 P2_add_898_U203 ( .IN1(P2_N2247), .IN2(P2_add_898_n193), 
        .QN(P2_add_898_n192) );
  NAND2X0 P2_add_898_U202 ( .IN1(P2_add_898_n191), .IN2(P2_add_898_n192), 
        .QN(P2_add_898_n184) );
  OR2X1 P2_add_898_U200 ( .IN2(P2_N2248), .IN1(n7197), .Q(P2_add_898_n188) );
  NAND2X0 P2_add_898_U199 ( .IN1(P2_N2248), .IN2(n7197), .QN(P2_add_898_n189)
         );
  NAND2X0 P2_add_898_U198 ( .IN1(P2_add_898_n188), .IN2(P2_add_898_n189), 
        .QN(P2_add_898_n187) );
  NOR2X0 P2_add_898_U197 ( .QN(P2_add_898_n185), .IN1(P2_add_898_n184), 
        .IN2(P2_add_898_n187) );
  AND2X1 P2_add_898_U196 ( .IN1(P2_add_898_n184), .IN2(P2_add_898_n187), 
        .Q(P2_add_898_n186) );
  NOR2X0 P2_add_898_U195 ( .QN(P2_N2490), .IN1(P2_add_898_n185), 
        .IN2(P2_add_898_n186) );
  NAND2X0 P2_add_898_U194 ( .IN1(P2_N5087), .IN2(P2_add_898_n184), 
        .QN(P2_add_898_n181) );
  OR2X1 P2_add_898_U193 ( .IN2(P2_N5087), .IN1(P2_add_898_n184), 
        .Q(P2_add_898_n183) );
  NAND2X0 P2_add_898_U192 ( .IN1(P2_N2248), .IN2(P2_add_898_n183), 
        .QN(P2_add_898_n182) );
  NAND2X0 P2_add_898_U191 ( .IN1(P2_add_898_n181), .IN2(P2_add_898_n182), 
        .QN(P2_add_898_n174) );
  OR2X1 P2_add_898_U189 ( .IN2(P2_N2249), .IN1(n7195), .Q(P2_add_898_n178) );
  NAND2X0 P2_add_898_U188 ( .IN1(P2_N2249), .IN2(n7195), .QN(P2_add_898_n179)
         );
  NAND2X0 P2_add_898_U187 ( .IN1(P2_add_898_n178), .IN2(P2_add_898_n179), 
        .QN(P2_add_898_n177) );
  NOR2X0 P2_add_898_U186 ( .QN(P2_add_898_n175), .IN1(P2_add_898_n174), 
        .IN2(P2_add_898_n177) );
  AND2X1 P2_add_898_U185 ( .IN1(P2_add_898_n174), .IN2(P2_add_898_n177), 
        .Q(P2_add_898_n176) );
  NOR2X0 P2_add_898_U184 ( .QN(P2_N2491), .IN1(P2_add_898_n175), 
        .IN2(P2_add_898_n176) );
  NAND2X0 P2_add_898_U183 ( .IN1(P2_N5088), .IN2(P2_add_898_n174), 
        .QN(P2_add_898_n171) );
  OR2X1 P2_add_898_U182 ( .IN2(P2_N5088), .IN1(P2_add_898_n174), 
        .Q(P2_add_898_n173) );
  NAND2X0 P2_add_898_U181 ( .IN1(P2_N2249), .IN2(P2_add_898_n173), 
        .QN(P2_add_898_n172) );
  NAND2X0 P2_add_898_U180 ( .IN1(P2_add_898_n171), .IN2(P2_add_898_n172), 
        .QN(P2_add_898_n164) );
  OR2X1 P2_add_898_U178 ( .IN2(P2_N2250), .IN1(n7188), .Q(P2_add_898_n168) );
  NAND2X0 P2_add_898_U177 ( .IN1(P2_N2250), .IN2(n7188), .QN(P2_add_898_n169)
         );
  NAND2X0 P2_add_898_U176 ( .IN1(P2_add_898_n168), .IN2(P2_add_898_n169), 
        .QN(P2_add_898_n167) );
  NOR2X0 P2_add_898_U175 ( .QN(P2_add_898_n165), .IN1(P2_add_898_n164), 
        .IN2(P2_add_898_n167) );
  AND2X1 P2_add_898_U174 ( .IN1(P2_add_898_n164), .IN2(P2_add_898_n167), 
        .Q(P2_add_898_n166) );
  NOR2X0 P2_add_898_U173 ( .QN(P2_N2492), .IN1(P2_add_898_n165), 
        .IN2(P2_add_898_n166) );
  NAND2X0 P2_add_898_U172 ( .IN1(P2_N5089), .IN2(P2_add_898_n164), 
        .QN(P2_add_898_n161) );
  OR2X1 P2_add_898_U171 ( .IN2(P2_N5089), .IN1(P2_add_898_n164), 
        .Q(P2_add_898_n163) );
  NAND2X0 P2_add_898_U170 ( .IN1(P2_N2250), .IN2(P2_add_898_n163), 
        .QN(P2_add_898_n162) );
  NAND2X0 P2_add_898_U169 ( .IN1(P2_add_898_n161), .IN2(P2_add_898_n162), 
        .QN(P2_add_898_n147) );
  OR2X1 P2_add_898_U167 ( .IN2(P2_N2251), .IN1(n7264), .Q(P2_add_898_n158) );
  NAND2X0 P2_add_898_U166 ( .IN1(P2_N2251), .IN2(n7264), .QN(P2_add_898_n159)
         );
  NAND2X0 P2_add_898_U165 ( .IN1(P2_add_898_n158), .IN2(P2_add_898_n159), 
        .QN(P2_add_898_n157) );
  NOR2X0 P2_add_898_U164 ( .QN(P2_add_898_n155), .IN1(P2_add_898_n147), 
        .IN2(P2_add_898_n157) );
  AND2X1 P2_add_898_U163 ( .IN1(P2_add_898_n147), .IN2(P2_add_898_n157), 
        .Q(P2_add_898_n156) );
  NOR2X0 P2_add_898_U162 ( .QN(P2_N2493), .IN1(P2_add_898_n155), 
        .IN2(P2_add_898_n156) );
  OR2X1 P2_add_898_U161 ( .IN2(P2_N2233), .IN1(n7184), .Q(P2_add_898_n152) );
  NAND2X0 P2_add_898_U160 ( .IN1(P2_N2233), .IN2(n7184), .QN(P2_add_898_n153)
         );
  NAND2X0 P2_add_898_U159 ( .IN1(P2_add_898_n152), .IN2(P2_add_898_n153), 
        .QN(P2_add_898_n150) );
  NAND2X0 P2_add_898_U158 ( .IN1(P2_add_898_n150), .IN2(P2_add_898_n151), 
        .QN(P2_add_898_n148) );
  OR2X1 P2_add_898_U157 ( .IN2(P2_add_898_n151), .IN1(P2_add_898_n150), 
        .Q(P2_add_898_n149) );
  OR2X1 P2_add_898_U308 ( .IN2(P2_N2232), .IN1(n2919), .Q(P2_add_898_n278) );
  NAND2X0 P2_add_898_U307 ( .IN1(P2_N2232), .IN2(n2919), .QN(P2_add_898_n279)
         );
  NAND2X0 P2_add_898_U306 ( .IN1(P2_add_898_n278), .IN2(P2_add_898_n279), 
        .QN(P2_N2474) );
  NAND2X0 P2_add_898_U304 ( .IN1(P2_N2232), .IN2(n7035), .QN(P2_add_898_n151)
         );
  OR2X1 P2_add_898_U303 ( .IN2(P2_add_898_n151), .IN1(n7184), 
        .Q(P2_add_898_n275) );
  NAND2X0 P2_add_898_U302 ( .IN1(n7184), .IN2(P2_add_898_n151), 
        .QN(P2_add_898_n277) );
  NAND2X0 P2_add_898_U301 ( .IN1(P2_N2233), .IN2(P2_add_898_n277), 
        .QN(P2_add_898_n276) );
  NAND2X0 P2_add_898_U300 ( .IN1(P2_add_898_n275), .IN2(P2_add_898_n276), 
        .QN(P2_add_898_n52) );
  NAND2X0 P2_add_898_U299 ( .IN1(P2_N5073), .IN2(P2_add_898_n52), 
        .QN(P2_add_898_n272) );
  OR2X1 P2_add_898_U298 ( .IN2(P2_N5073), .IN1(P2_add_898_n52), 
        .Q(P2_add_898_n274) );
  NAND2X0 P2_add_898_U297 ( .IN1(P2_N2234), .IN2(P2_add_898_n274), 
        .QN(P2_add_898_n273) );
  NAND2X0 P2_add_898_U296 ( .IN1(P2_add_898_n272), .IN2(P2_add_898_n273), 
        .QN(P2_add_898_n45) );
  NAND2X0 P2_add_898_U295 ( .IN1(P2_N5074), .IN2(P2_add_898_n45), 
        .QN(P2_add_898_n269) );
  OR2X1 P2_add_898_U294 ( .IN2(P2_N5074), .IN1(P2_add_898_n45), 
        .Q(P2_add_898_n271) );
  NAND2X0 P2_add_898_U293 ( .IN1(P2_N2235), .IN2(P2_add_898_n271), 
        .QN(P2_add_898_n270) );
  NAND2X0 P2_add_898_U292 ( .IN1(P2_add_898_n269), .IN2(P2_add_898_n270), 
        .QN(P2_add_898_n38) );
  NAND2X0 P2_add_898_U291 ( .IN1(P2_N5075), .IN2(P2_add_898_n38), 
        .QN(P2_add_898_n266) );
  OR2X1 P2_add_898_U290 ( .IN2(P2_N5075), .IN1(P2_add_898_n38), 
        .Q(P2_add_898_n268) );
  NAND2X0 P2_add_898_U289 ( .IN1(P2_N2236), .IN2(P2_add_898_n268), 
        .QN(P2_add_898_n267) );
  NAND2X0 P2_add_898_U288 ( .IN1(P2_add_898_n266), .IN2(P2_add_898_n267), 
        .QN(P2_add_898_n31) );
  NAND2X0 P2_add_898_U287 ( .IN1(P2_N5076), .IN2(P2_add_898_n31), 
        .QN(P2_add_898_n263) );
  OR2X1 P2_add_898_U286 ( .IN2(P2_N5076), .IN1(P2_add_898_n31), 
        .Q(P2_add_898_n265) );
  NAND2X0 P2_add_898_U285 ( .IN1(P2_N2237), .IN2(P2_add_898_n265), 
        .QN(P2_add_898_n264) );
  NAND2X0 P2_add_898_U284 ( .IN1(P2_add_898_n263), .IN2(P2_add_898_n264), 
        .QN(P2_add_898_n24) );
  NAND2X0 P2_add_898_U283 ( .IN1(n7162), .IN2(P2_add_898_n24), 
        .QN(P2_add_898_n260) );
  OR2X1 P2_add_898_U282 ( .IN2(n7162), .IN1(P2_add_898_n24), 
        .Q(P2_add_898_n262) );
  NAND2X0 P2_add_898_U281 ( .IN1(P2_N2238), .IN2(P2_add_898_n262), 
        .QN(P2_add_898_n261) );
  NAND2X0 P2_add_898_U280 ( .IN1(P2_add_898_n260), .IN2(P2_add_898_n261), 
        .QN(P2_add_898_n17) );
  NAND2X0 P2_add_898_U279 ( .IN1(n7158), .IN2(P2_add_898_n17), 
        .QN(P2_add_898_n257) );
  OR2X1 P2_add_898_U278 ( .IN2(n7158), .IN1(P2_add_898_n17), 
        .Q(P2_add_898_n259) );
  NAND2X0 P2_add_898_U277 ( .IN1(P2_N2239), .IN2(P2_add_898_n259), 
        .QN(P2_add_898_n258) );
  NAND2X0 P2_add_898_U276 ( .IN1(P2_add_898_n257), .IN2(P2_add_898_n258), 
        .QN(P2_add_898_n10) );
  NAND2X0 P2_add_898_U275 ( .IN1(n7154), .IN2(P2_add_898_n10), 
        .QN(P2_add_898_n254) );
  OR2X1 P2_add_898_U274 ( .IN2(n7154), .IN1(P2_add_898_n10), 
        .Q(P2_add_898_n256) );
  NAND2X0 P2_add_898_U273 ( .IN1(P2_N2240), .IN2(P2_add_898_n256), 
        .QN(P2_add_898_n255) );
  NAND2X0 P2_add_898_U272 ( .IN1(P2_add_898_n254), .IN2(P2_add_898_n255), 
        .QN(P2_add_898_n3) );
  NAND2X0 P2_add_898_U271 ( .IN1(n7151), .IN2(P2_add_898_n3), 
        .QN(P2_add_898_n251) );
  OR2X1 P2_add_898_U270 ( .IN2(n7151), .IN1(P2_add_898_n3), 
        .Q(P2_add_898_n253) );
  NAND2X0 P2_add_898_U269 ( .IN1(P2_N2241), .IN2(P2_add_898_n253), 
        .QN(P2_add_898_n252) );
  NAND2X0 P2_add_898_U268 ( .IN1(P2_add_898_n251), .IN2(P2_add_898_n252), 
        .QN(P2_add_898_n244) );
  OR2X1 P2_add_898_U266 ( .IN2(P2_N2242), .IN1(n7219), .Q(P2_add_898_n248) );
  NAND2X0 P2_add_898_U265 ( .IN1(P2_N2242), .IN2(n7219), .QN(P2_add_898_n249)
         );
  NAND2X0 P2_add_898_U264 ( .IN1(P2_add_898_n248), .IN2(P2_add_898_n249), 
        .QN(P2_add_898_n247) );
  NOR2X0 P2_add_898_U263 ( .QN(P2_add_898_n245), .IN1(P2_add_898_n244), 
        .IN2(P2_add_898_n247) );
  AND2X1 P2_add_898_U262 ( .IN1(P2_add_898_n244), .IN2(P2_add_898_n247), 
        .Q(P2_add_898_n246) );
  NOR2X0 P2_add_898_U261 ( .QN(P2_N2484), .IN1(P2_add_898_n245), 
        .IN2(P2_add_898_n246) );
  NAND2X0 P2_add_898_U260 ( .IN1(n7220), .IN2(P2_add_898_n244), 
        .QN(P2_add_898_n241) );
  OR2X1 P2_add_898_U259 ( .IN2(n7220), .IN1(P2_add_898_n244), 
        .Q(P2_add_898_n243) );
  NAND2X0 P2_add_898_U258 ( .IN1(P2_N2242), .IN2(P2_add_898_n243), 
        .QN(P2_add_898_n242) );
  NAND2X0 P2_add_898_U257 ( .IN1(P2_add_898_n241), .IN2(P2_add_898_n242), 
        .QN(P2_add_898_n234) );
  OR2X1 P2_add_898_U255 ( .IN2(P2_N2243), .IN1(n7214), .Q(P2_add_898_n238) );
  NAND2X0 P2_add_898_U254 ( .IN1(P2_N2243), .IN2(n7214), .QN(P2_add_898_n239)
         );
  NAND2X0 P2_add_898_U253 ( .IN1(P2_add_898_n238), .IN2(P2_add_898_n239), 
        .QN(P2_add_898_n237) );
  NOR2X0 P2_add_898_U252 ( .QN(P2_add_898_n235), .IN1(P2_add_898_n234), 
        .IN2(P2_add_898_n237) );
  AND2X1 P2_add_898_U251 ( .IN1(P2_add_898_n234), .IN2(P2_add_898_n237), 
        .Q(P2_add_898_n236) );
  NOR2X0 P2_add_898_U250 ( .QN(P2_N2485), .IN1(P2_add_898_n235), 
        .IN2(P2_add_898_n236) );
  INVX0 P2_add_898_U7 ( .ZN(P2_add_898_n299), .INP(P2_N5094) );
  AND2X1 P1_sub_273_U29 ( .IN1(P1_sub_273_n26), .IN2(P1_N632), 
        .Q(P1_sub_273_n24) );
  NOR2X0 P1_sub_273_U28 ( .QN(P1_sub_273_n25), .IN1(P1_N632), 
        .IN2(P1_sub_273_n26) );
  NOR2X0 P1_sub_273_U27 ( .QN(P1_N882), .IN1(P1_sub_273_n24), 
        .IN2(P1_sub_273_n25) );
  AND2X1 P1_sub_273_U26 ( .IN1(P1_sub_273_n21), .IN2(P1_N633), 
        .Q(P1_sub_273_n22) );
  NOR2X0 P1_sub_273_U25 ( .QN(P1_sub_273_n23), .IN1(P1_N633), 
        .IN2(P1_sub_273_n21) );
  NOR2X0 P1_sub_273_U24 ( .QN(P1_N883), .IN1(P1_sub_273_n22), 
        .IN2(P1_sub_273_n23) );
  OR2X1 P1_sub_273_U23 ( .IN2(P1_N633), .IN1(P1_sub_273_n21), 
        .Q(P1_sub_273_n20) );
  AND2X1 P1_sub_273_U22 ( .IN1(P1_sub_273_n20), .IN2(P1_N634), 
        .Q(P1_sub_273_n18) );
  NOR2X0 P1_sub_273_U21 ( .QN(P1_sub_273_n19), .IN1(P1_N634), 
        .IN2(P1_sub_273_n20) );
  NOR2X0 P1_sub_273_U20 ( .QN(P1_N884), .IN1(P1_sub_273_n18), 
        .IN2(P1_sub_273_n19) );
  INVX0 P1_sub_273_U19 ( .ZN(P1_sub_273_n14), .INP(P1_sub_273_n17) );
  AND2X1 P1_sub_273_U18 ( .IN1(P1_sub_273_n14), .IN2(P1_N635), 
        .Q(P1_sub_273_n15) );
  NOR2X0 P1_sub_273_U17 ( .QN(P1_sub_273_n16), .IN1(P1_N635), 
        .IN2(P1_sub_273_n14) );
  NOR2X0 P1_sub_273_U16 ( .QN(P1_N885), .IN1(P1_sub_273_n15), 
        .IN2(P1_sub_273_n16) );
  OR2X1 P1_sub_273_U15 ( .IN2(P1_N635), .IN1(P1_sub_273_n14), 
        .Q(P1_sub_273_n13) );
  AND2X1 P1_sub_273_U14 ( .IN1(P1_sub_273_n13), .IN2(P1_N636), 
        .Q(P1_sub_273_n11) );
  NOR2X0 P1_sub_273_U13 ( .QN(P1_sub_273_n12), .IN1(P1_N636), 
        .IN2(P1_sub_273_n13) );
  NOR2X0 P1_sub_273_U12 ( .QN(P1_N886), .IN1(P1_sub_273_n11), 
        .IN2(P1_sub_273_n12) );
  AND2X1 P1_sub_273_U11 ( .IN1(P1_sub_273_n8), .IN2(P1_N637), 
        .Q(P1_sub_273_n9) );
  NOR2X0 P1_sub_273_U10 ( .QN(P1_sub_273_n10), .IN1(P1_N637), 
        .IN2(P1_sub_273_n8) );
  NOR2X0 P1_sub_273_U9 ( .QN(P1_N887), .IN1(P1_sub_273_n9), 
        .IN2(P1_sub_273_n10) );
  OR2X1 P1_sub_273_U8 ( .IN2(P1_N637), .IN1(P1_sub_273_n8), .Q(P1_sub_273_n7)
         );
  AND2X1 P1_sub_273_U7 ( .IN1(P1_sub_273_n7), .IN2(P1_N638), .Q(P1_sub_273_n5)
         );
  NOR2X0 P1_sub_273_U6 ( .QN(P1_sub_273_n6), .IN1(P1_N638), 
        .IN2(P1_sub_273_n7) );
  NOR2X0 P1_sub_273_U5 ( .QN(P1_N888), .IN1(P1_sub_273_n5), 
        .IN2(P1_sub_273_n6) );
  AND2X1 P1_sub_273_U4 ( .IN1(P1_sub_273_n4), .IN2(P1_N639), .Q(P1_sub_273_n2)
         );
  NOR2X0 P1_sub_273_U3 ( .QN(P1_sub_273_n3), .IN1(P1_N639), 
        .IN2(P1_sub_273_n4) );
  NOR2X0 P1_sub_273_U2 ( .QN(P1_N889), .IN1(P1_sub_273_n2), 
        .IN2(P1_sub_273_n3) );
  OR2X1 P1_sub_273_U122 ( .IN2(P1_N639), .IN1(P1_sub_273_n4), 
        .Q(P1_sub_273_n100) );
  AND2X1 P1_sub_273_U121 ( .IN1(P1_sub_273_n100), .IN2(P1_N640), 
        .Q(P1_sub_273_n98) );
  NOR2X0 P1_sub_273_U120 ( .QN(P1_sub_273_n99), .IN1(P1_N640), 
        .IN2(P1_sub_273_n100) );
  NOR2X0 P1_sub_273_U119 ( .QN(P1_N890), .IN1(P1_sub_273_n98), 
        .IN2(P1_sub_273_n99) );
  NOR2X0 P1_sub_273_U118 ( .QN(P1_sub_273_n96), .IN1(P1_N639), .IN2(P1_N640)
         );
  NAND2X0 P1_sub_273_U117 ( .IN1(P1_sub_273_n96), .IN2(P1_sub_273_n97), 
        .QN(P1_sub_273_n90) );
  AND2X1 P1_sub_273_U116 ( .IN1(P1_sub_273_n90), .IN2(P1_N641), 
        .Q(P1_sub_273_n94) );
  NOR2X0 P1_sub_273_U115 ( .QN(P1_sub_273_n95), .IN1(P1_N641), 
        .IN2(P1_sub_273_n90) );
  NOR2X0 P1_sub_273_U114 ( .QN(P1_N891), .IN1(P1_sub_273_n94), 
        .IN2(P1_sub_273_n95) );
  OR2X1 P1_sub_273_U113 ( .IN2(P1_N641), .IN1(P1_sub_273_n90), 
        .Q(P1_sub_273_n93) );
  AND2X1 P1_sub_273_U112 ( .IN1(P1_sub_273_n93), .IN2(P1_N642), 
        .Q(P1_sub_273_n91) );
  NOR2X0 P1_sub_273_U111 ( .QN(P1_sub_273_n92), .IN1(P1_N642), 
        .IN2(P1_sub_273_n93) );
  NOR2X0 P1_sub_273_U110 ( .QN(P1_N892), .IN1(P1_sub_273_n91), 
        .IN2(P1_sub_273_n92) );
  OR2X1 P1_sub_273_U109 ( .IN2(P1_N641), .IN1(P1_N642), .Q(P1_sub_273_n89) );
  NOR2X0 P1_sub_273_U108 ( .QN(P1_sub_273_n82), .IN1(P1_sub_273_n89), 
        .IN2(P1_sub_273_n90) );
  INVX0 P1_sub_273_U107 ( .ZN(P1_sub_273_n86), .INP(P1_sub_273_n82) );
  AND2X1 P1_sub_273_U106 ( .IN1(P1_sub_273_n86), .IN2(P1_N643), 
        .Q(P1_sub_273_n87) );
  NOR2X0 P1_sub_273_U105 ( .QN(P1_sub_273_n88), .IN1(P1_N643), 
        .IN2(P1_sub_273_n86) );
  NOR2X0 P1_sub_273_U104 ( .QN(P1_N893), .IN1(P1_sub_273_n87), 
        .IN2(P1_sub_273_n88) );
  OR2X1 P1_sub_273_U103 ( .IN2(P1_N643), .IN1(P1_sub_273_n86), 
        .Q(P1_sub_273_n85) );
  AND2X1 P1_sub_273_U102 ( .IN1(P1_sub_273_n85), .IN2(P1_N644), 
        .Q(P1_sub_273_n83) );
  NOR2X0 P1_sub_273_U101 ( .QN(P1_sub_273_n84), .IN1(P1_N644), 
        .IN2(P1_sub_273_n85) );
  NOR2X0 P1_sub_273_U100 ( .QN(P1_N894), .IN1(P1_sub_273_n83), 
        .IN2(P1_sub_273_n84) );
  NOR2X0 P1_sub_273_U99 ( .QN(P1_sub_273_n81), .IN1(P1_N644), .IN2(P1_N643) );
  NAND2X0 P1_sub_273_U98 ( .IN1(P1_sub_273_n81), .IN2(P1_sub_273_n82), 
        .QN(P1_sub_273_n75) );
  AND2X1 P1_sub_273_U97 ( .IN1(P1_sub_273_n75), .IN2(P1_N645), 
        .Q(P1_sub_273_n79) );
  NOR2X0 P1_sub_273_U96 ( .QN(P1_sub_273_n80), .IN1(P1_N645), 
        .IN2(P1_sub_273_n75) );
  NOR2X0 P1_sub_273_U95 ( .QN(P1_N895), .IN1(P1_sub_273_n79), 
        .IN2(P1_sub_273_n80) );
  OR2X1 P1_sub_273_U94 ( .IN2(P1_N645), .IN1(P1_sub_273_n75), 
        .Q(P1_sub_273_n78) );
  AND2X1 P1_sub_273_U93 ( .IN1(P1_sub_273_n78), .IN2(P1_N646), 
        .Q(P1_sub_273_n76) );
  NOR2X0 P1_sub_273_U92 ( .QN(P1_sub_273_n77), .IN1(P1_N646), 
        .IN2(P1_sub_273_n78) );
  NOR2X0 P1_sub_273_U91 ( .QN(P1_N896), .IN1(P1_sub_273_n76), 
        .IN2(P1_sub_273_n77) );
  OR2X1 P1_sub_273_U90 ( .IN2(P1_N645), .IN1(P1_N646), .Q(P1_sub_273_n74) );
  NOR2X0 P1_sub_273_U89 ( .QN(P1_sub_273_n67), .IN1(P1_sub_273_n74), 
        .IN2(P1_sub_273_n75) );
  INVX0 P1_sub_273_U88 ( .ZN(P1_sub_273_n71), .INP(P1_sub_273_n67) );
  AND2X1 P1_sub_273_U87 ( .IN1(P1_sub_273_n71), .IN2(P1_N647), 
        .Q(P1_sub_273_n72) );
  NOR2X0 P1_sub_273_U86 ( .QN(P1_sub_273_n73), .IN1(P1_N647), 
        .IN2(P1_sub_273_n71) );
  NOR2X0 P1_sub_273_U85 ( .QN(P1_N897), .IN1(P1_sub_273_n72), 
        .IN2(P1_sub_273_n73) );
  OR2X1 P1_sub_273_U84 ( .IN2(P1_N647), .IN1(P1_sub_273_n71), 
        .Q(P1_sub_273_n70) );
  AND2X1 P1_sub_273_U83 ( .IN1(P1_sub_273_n70), .IN2(P1_N648), 
        .Q(P1_sub_273_n68) );
  NOR2X0 P1_sub_273_U82 ( .QN(P1_sub_273_n69), .IN1(P1_N648), 
        .IN2(P1_sub_273_n70) );
  NOR2X0 P1_sub_273_U81 ( .QN(P1_N898), .IN1(P1_sub_273_n68), 
        .IN2(P1_sub_273_n69) );
  NOR2X0 P1_sub_273_U80 ( .QN(P1_sub_273_n66), .IN1(P1_N648), .IN2(P1_N647) );
  NAND2X0 P1_sub_273_U79 ( .IN1(P1_sub_273_n66), .IN2(P1_sub_273_n67), 
        .QN(P1_sub_273_n57) );
  AND2X1 P1_sub_273_U78 ( .IN1(P1_sub_273_n57), .IN2(P1_N649), 
        .Q(P1_sub_273_n64) );
  NOR2X0 P1_sub_273_U77 ( .QN(P1_sub_273_n65), .IN1(P1_N649), 
        .IN2(P1_sub_273_n57) );
  NOR2X0 P1_sub_273_U76 ( .QN(P1_N899), .IN1(P1_sub_273_n64), 
        .IN2(P1_sub_273_n65) );
  OR2X1 P1_sub_273_U75 ( .IN2(P1_N631), .IN1(n7274), .Q(P1_sub_273_n61) );
  NAND2X0 P1_sub_273_U74 ( .IN1(P1_N631), .IN2(n7274), .QN(P1_sub_273_n62) );
  NAND2X0 P1_sub_273_U73 ( .IN1(P1_sub_273_n61), .IN2(P1_sub_273_n62), 
        .QN(P1_N881) );
  OR2X1 P1_sub_273_U72 ( .IN2(P1_N649), .IN1(P1_sub_273_n57), 
        .Q(P1_sub_273_n60) );
  AND2X1 P1_sub_273_U71 ( .IN1(P1_sub_273_n60), .IN2(P1_N650), 
        .Q(P1_sub_273_n58) );
  NOR2X0 P1_sub_273_U70 ( .QN(P1_sub_273_n59), .IN1(P1_N650), 
        .IN2(P1_sub_273_n60) );
  NOR2X0 P1_sub_273_U69 ( .QN(P1_N900), .IN1(P1_sub_273_n58), 
        .IN2(P1_sub_273_n59) );
  OR2X1 P1_sub_273_U68 ( .IN2(P1_N649), .IN1(P1_N650), .Q(P1_sub_273_n56) );
  NOR2X0 P1_sub_273_U67 ( .QN(P1_sub_273_n49), .IN1(P1_sub_273_n56), 
        .IN2(P1_sub_273_n57) );
  INVX0 P1_sub_273_U66 ( .ZN(P1_sub_273_n53), .INP(P1_sub_273_n49) );
  AND2X1 P1_sub_273_U65 ( .IN1(P1_sub_273_n53), .IN2(P1_N651), 
        .Q(P1_sub_273_n54) );
  NOR2X0 P1_sub_273_U64 ( .QN(P1_sub_273_n55), .IN1(P1_N651), 
        .IN2(P1_sub_273_n53) );
  NOR2X0 P1_sub_273_U63 ( .QN(P1_N901), .IN1(P1_sub_273_n54), 
        .IN2(P1_sub_273_n55) );
  OR2X1 P1_sub_273_U62 ( .IN2(P1_N651), .IN1(P1_sub_273_n53), 
        .Q(P1_sub_273_n52) );
  AND2X1 P1_sub_273_U61 ( .IN1(P1_sub_273_n52), .IN2(P1_N652), 
        .Q(P1_sub_273_n50) );
  NOR2X0 P1_sub_273_U60 ( .QN(P1_sub_273_n51), .IN1(P1_N652), 
        .IN2(P1_sub_273_n52) );
  NOR2X0 P1_sub_273_U59 ( .QN(P1_N902), .IN1(P1_sub_273_n50), 
        .IN2(P1_sub_273_n51) );
  NOR2X0 P1_sub_273_U58 ( .QN(P1_sub_273_n48), .IN1(P1_N652), .IN2(P1_N651) );
  NAND2X0 P1_sub_273_U57 ( .IN1(P1_sub_273_n48), .IN2(P1_sub_273_n49), 
        .QN(P1_sub_273_n42) );
  AND2X1 P1_sub_273_U56 ( .IN1(P1_sub_273_n42), .IN2(P1_N653), 
        .Q(P1_sub_273_n46) );
  NOR2X0 P1_sub_273_U55 ( .QN(P1_sub_273_n47), .IN1(P1_N653), 
        .IN2(P1_sub_273_n42) );
  NOR2X0 P1_sub_273_U54 ( .QN(P1_N903), .IN1(P1_sub_273_n46), 
        .IN2(P1_sub_273_n47) );
  OR2X1 P1_sub_273_U53 ( .IN2(P1_N653), .IN1(P1_sub_273_n42), 
        .Q(P1_sub_273_n45) );
  AND2X1 P1_sub_273_U52 ( .IN1(P1_sub_273_n45), .IN2(P1_N654), 
        .Q(P1_sub_273_n43) );
  NOR2X0 P1_sub_273_U51 ( .QN(P1_sub_273_n44), .IN1(P1_N654), 
        .IN2(P1_sub_273_n45) );
  NOR2X0 P1_sub_273_U50 ( .QN(P1_N904), .IN1(P1_sub_273_n43), 
        .IN2(P1_sub_273_n44) );
  OR2X1 P1_sub_273_U49 ( .IN2(P1_N653), .IN1(P1_N654), .Q(P1_sub_273_n41) );
  NOR2X0 P1_sub_273_U48 ( .QN(P1_sub_273_n34), .IN1(P1_sub_273_n41), 
        .IN2(P1_sub_273_n42) );
  INVX0 P1_sub_273_U47 ( .ZN(P1_sub_273_n38), .INP(P1_sub_273_n34) );
  AND2X1 P1_sub_273_U46 ( .IN1(P1_sub_273_n38), .IN2(P1_N655), 
        .Q(P1_sub_273_n39) );
  NOR2X0 P1_sub_273_U45 ( .QN(P1_sub_273_n40), .IN1(P1_N655), 
        .IN2(P1_sub_273_n38) );
  NOR2X0 P1_sub_273_U44 ( .QN(P1_N905), .IN1(P1_sub_273_n39), 
        .IN2(P1_sub_273_n40) );
  OR2X1 P1_sub_273_U43 ( .IN2(P1_N655), .IN1(P1_sub_273_n38), 
        .Q(P1_sub_273_n37) );
  AND2X1 P1_sub_273_U42 ( .IN1(P1_sub_273_n37), .IN2(P1_N656), 
        .Q(P1_sub_273_n35) );
  NOR2X0 P1_sub_273_U41 ( .QN(P1_sub_273_n36), .IN1(P1_N656), 
        .IN2(P1_sub_273_n37) );
  NOR2X0 P1_sub_273_U40 ( .QN(P1_N906), .IN1(P1_sub_273_n35), 
        .IN2(P1_sub_273_n36) );
  NOR2X0 P1_sub_273_U39 ( .QN(P1_sub_273_n33), .IN1(P1_N656), .IN2(P1_N655) );
  NAND2X0 P1_sub_273_U38 ( .IN1(P1_sub_273_n33), .IN2(P1_sub_273_n34), 
        .QN(P1_sub_273_n30) );
  AND2X1 P1_sub_273_U37 ( .IN1(P1_sub_273_n30), .IN2(P1_N657), 
        .Q(P1_sub_273_n31) );
  NOR2X0 P1_sub_273_U36 ( .QN(P1_sub_273_n32), .IN1(P1_N657), 
        .IN2(P1_sub_273_n30) );
  NOR2X0 P1_sub_273_U35 ( .QN(P1_N907), .IN1(P1_sub_273_n31), 
        .IN2(P1_sub_273_n32) );
  OR2X1 P1_sub_273_U34 ( .IN2(P1_N657), .IN1(P1_sub_273_n30), 
        .Q(P1_sub_273_n29) );
  AND2X1 P1_sub_273_U33 ( .IN1(P1_sub_273_n29), .IN2(P1_N658), 
        .Q(P1_sub_273_n27) );
  NOR2X0 P1_sub_273_U32 ( .QN(P1_sub_273_n28), .IN1(P1_N658), 
        .IN2(P1_sub_273_n29) );
  NOR2X0 P1_sub_273_U31 ( .QN(P1_N908), .IN1(P1_sub_273_n27), 
        .IN2(P1_sub_273_n28) );
  OR2X1 P1_sub_273_U30 ( .IN2(P1_N630), .IN1(P1_N631), .Q(P1_sub_273_n26) );
  OR2X1 P1_sub_273_U132 ( .IN2(P1_N637), .IN1(P1_N638), .Q(P1_sub_273_n101) );
  NOR2X0 P1_sub_273_U131 ( .QN(P1_sub_273_n102), .IN1(P1_N636), .IN2(P1_N635)
         );
  OR2X1 P1_sub_273_U130 ( .IN2(P1_N633), .IN1(P1_N634), .Q(P1_sub_273_n103) );
  NOR2X0 P1_sub_273_U129 ( .QN(P1_sub_273_n104), .IN1(P1_N632), .IN2(P1_N631)
         );
  NAND2X0 P1_sub_273_U127 ( .IN1(P1_sub_273_n104), .IN2(n7274), 
        .QN(P1_sub_273_n21) );
  NOR2X0 P1_sub_273_U126 ( .QN(P1_sub_273_n17), .IN1(P1_sub_273_n103), 
        .IN2(P1_sub_273_n21) );
  NAND2X0 P1_sub_273_U125 ( .IN1(P1_sub_273_n102), .IN2(P1_sub_273_n17), 
        .QN(P1_sub_273_n8) );
  NOR2X0 P1_sub_273_U124 ( .QN(P1_sub_273_n97), .IN1(P1_sub_273_n101), 
        .IN2(P1_sub_273_n8) );
  INVX0 P1_sub_273_U123 ( .ZN(P1_sub_273_n4), .INP(P1_sub_273_n97) );
  NOR2X0 P1_add_348_U59 ( .QN(P1_add_348_n57), .IN1(P1_add_348_n60), 
        .IN2(P1_add_348_n59) );
  AND2X1 P1_add_348_U58 ( .IN1(P1_add_348_n59), .IN2(P1_add_348_n60), 
        .Q(P1_add_348_n58) );
  NOR2X0 P1_add_348_U57 ( .QN(P1_N1882), .IN1(P1_add_348_n57), 
        .IN2(P1_add_348_n58) );
  OR2X1 P1_add_348_U55 ( .IN2(P1_N1614), .IN1(n7045), .Q(P1_add_348_n54) );
  NAND2X0 P1_add_348_U54 ( .IN1(P1_N1614), .IN2(n7045), .QN(P1_add_348_n55) );
  NAND2X0 P1_add_348_U53 ( .IN1(P1_add_348_n54), .IN2(P1_add_348_n55), 
        .QN(P1_add_348_n53) );
  NOR2X0 P1_add_348_U52 ( .QN(P1_add_348_n50), .IN1(P1_add_348_n52), 
        .IN2(P1_add_348_n53) );
  AND2X1 P1_add_348_U51 ( .IN1(P1_add_348_n52), .IN2(P1_add_348_n53), 
        .Q(P1_add_348_n51) );
  NOR2X0 P1_add_348_U50 ( .QN(P1_N1856), .IN1(P1_add_348_n50), 
        .IN2(P1_add_348_n51) );
  OR2X1 P1_add_348_U48 ( .IN2(P1_N1615), .IN1(n7043), .Q(P1_add_348_n47) );
  NAND2X0 P1_add_348_U47 ( .IN1(P1_N1615), .IN2(n7043), .QN(P1_add_348_n48) );
  NAND2X0 P1_add_348_U46 ( .IN1(P1_add_348_n47), .IN2(P1_add_348_n48), 
        .QN(P1_add_348_n46) );
  NOR2X0 P1_add_348_U45 ( .QN(P1_add_348_n43), .IN1(P1_add_348_n45), 
        .IN2(P1_add_348_n46) );
  AND2X1 P1_add_348_U44 ( .IN1(P1_add_348_n45), .IN2(P1_add_348_n46), 
        .Q(P1_add_348_n44) );
  NOR2X0 P1_add_348_U43 ( .QN(P1_N1857), .IN1(P1_add_348_n43), 
        .IN2(P1_add_348_n44) );
  OR2X1 P1_add_348_U41 ( .IN2(P1_N1616), .IN1(n7037), .Q(P1_add_348_n40) );
  NAND2X0 P1_add_348_U40 ( .IN1(P1_N1616), .IN2(n7037), .QN(P1_add_348_n41) );
  NAND2X0 P1_add_348_U39 ( .IN1(P1_add_348_n40), .IN2(P1_add_348_n41), 
        .QN(P1_add_348_n39) );
  NOR2X0 P1_add_348_U38 ( .QN(P1_add_348_n36), .IN1(P1_add_348_n38), 
        .IN2(P1_add_348_n39) );
  AND2X1 P1_add_348_U37 ( .IN1(P1_add_348_n38), .IN2(P1_add_348_n39), 
        .Q(P1_add_348_n37) );
  NOR2X0 P1_add_348_U36 ( .QN(P1_N1858), .IN1(P1_add_348_n36), 
        .IN2(P1_add_348_n37) );
  OR2X1 P1_add_348_U34 ( .IN2(P1_N1617), .IN1(n7082), .Q(P1_add_348_n33) );
  NAND2X0 P1_add_348_U33 ( .IN1(P1_N1617), .IN2(n7082), .QN(P1_add_348_n34) );
  NAND2X0 P1_add_348_U32 ( .IN1(P1_add_348_n33), .IN2(P1_add_348_n34), 
        .QN(P1_add_348_n32) );
  NOR2X0 P1_add_348_U31 ( .QN(P1_add_348_n29), .IN1(P1_add_348_n31), 
        .IN2(P1_add_348_n32) );
  AND2X1 P1_add_348_U30 ( .IN1(P1_add_348_n31), .IN2(P1_add_348_n32), 
        .Q(P1_add_348_n30) );
  NOR2X0 P1_add_348_U29 ( .QN(P1_N1859), .IN1(P1_add_348_n29), 
        .IN2(P1_add_348_n30) );
  OR2X1 P1_add_348_U27 ( .IN2(P1_N1618), .IN1(n7079), .Q(P1_add_348_n26) );
  NAND2X0 P1_add_348_U26 ( .IN1(P1_N1618), .IN2(n7079), .QN(P1_add_348_n27) );
  NAND2X0 P1_add_348_U25 ( .IN1(P1_add_348_n26), .IN2(P1_add_348_n27), 
        .QN(P1_add_348_n25) );
  NOR2X0 P1_add_348_U24 ( .QN(P1_add_348_n22), .IN1(P1_add_348_n24), 
        .IN2(P1_add_348_n25) );
  AND2X1 P1_add_348_U23 ( .IN1(P1_add_348_n24), .IN2(P1_add_348_n25), 
        .Q(P1_add_348_n23) );
  NOR2X0 P1_add_348_U22 ( .QN(P1_N1860), .IN1(P1_add_348_n22), 
        .IN2(P1_add_348_n23) );
  OR2X1 P1_add_348_U20 ( .IN2(P1_N1619), .IN1(n7076), .Q(P1_add_348_n19) );
  NAND2X0 P1_add_348_U19 ( .IN1(P1_N1619), .IN2(n7076), .QN(P1_add_348_n20) );
  NAND2X0 P1_add_348_U18 ( .IN1(P1_add_348_n19), .IN2(P1_add_348_n20), 
        .QN(P1_add_348_n18) );
  NOR2X0 P1_add_348_U17 ( .QN(P1_add_348_n15), .IN1(P1_add_348_n17), 
        .IN2(P1_add_348_n18) );
  AND2X1 P1_add_348_U16 ( .IN1(P1_add_348_n17), .IN2(P1_add_348_n18), 
        .Q(P1_add_348_n16) );
  NOR2X0 P1_add_348_U15 ( .QN(P1_N1861), .IN1(P1_add_348_n15), 
        .IN2(P1_add_348_n16) );
  OR2X1 P1_add_348_U13 ( .IN2(P1_N1620), .IN1(P1_add_348_n180), 
        .Q(P1_add_348_n12) );
  NAND2X0 P1_add_348_U12 ( .IN1(P1_N1620), .IN2(P1_add_348_n180), 
        .QN(P1_add_348_n13) );
  NAND2X0 P1_add_348_U11 ( .IN1(P1_add_348_n12), .IN2(P1_add_348_n13), 
        .QN(P1_add_348_n11) );
  NOR2X0 P1_add_348_U10 ( .QN(P1_add_348_n8), .IN1(P1_add_348_n10), 
        .IN2(P1_add_348_n11) );
  AND2X1 P1_add_348_U9 ( .IN1(P1_add_348_n10), .IN2(P1_add_348_n11), 
        .Q(P1_add_348_n9) );
  NOR2X0 P1_add_348_U8 ( .QN(P1_N1862), .IN1(P1_add_348_n8), 
        .IN2(P1_add_348_n9) );
  OR2X1 P1_add_348_U6 ( .IN2(P1_N1621), .IN1(n7071), .Q(P1_add_348_n5) );
  NAND2X0 P1_add_348_U5 ( .IN1(P1_N1621), .IN2(n7071), .QN(P1_add_348_n6) );
  NAND2X0 P1_add_348_U4 ( .IN1(P1_add_348_n5), .IN2(P1_add_348_n6), 
        .QN(P1_add_348_n4) );
  NOR2X0 P1_add_348_U3 ( .QN(P1_add_348_n1), .IN1(P1_add_348_n3), 
        .IN2(P1_add_348_n4) );
  AND2X1 P1_add_348_U2 ( .IN1(P1_add_348_n3), .IN2(P1_add_348_n4), 
        .Q(P1_add_348_n2) );
  NOR2X0 P1_add_348_U1 ( .QN(P1_N1863), .IN1(P1_add_348_n1), 
        .IN2(P1_add_348_n2) );
  NAND2X0 P1_add_348_U152 ( .IN1(P1_add_348_n144), .IN2(P1_add_348_n145), 
        .QN(P1_add_348_n137) );
  OR2X1 P1_add_348_U150 ( .IN2(P1_N1632), .IN1(n7095), .Q(P1_add_348_n141) );
  NAND2X0 P1_add_348_U149 ( .IN1(P1_N1632), .IN2(n7095), .QN(P1_add_348_n142)
         );
  NAND2X0 P1_add_348_U148 ( .IN1(P1_add_348_n141), .IN2(P1_add_348_n142), 
        .QN(P1_add_348_n140) );
  NOR2X0 P1_add_348_U147 ( .QN(P1_add_348_n138), .IN1(P1_add_348_n137), 
        .IN2(P1_add_348_n140) );
  AND2X1 P1_add_348_U146 ( .IN1(P1_add_348_n137), .IN2(P1_add_348_n140), 
        .Q(P1_add_348_n139) );
  NOR2X0 P1_add_348_U145 ( .QN(P1_N1874), .IN1(P1_add_348_n138), 
        .IN2(P1_add_348_n139) );
  NAND2X0 P1_add_348_U144 ( .IN1(P1_N5169), .IN2(P1_add_348_n137), 
        .QN(P1_add_348_n134) );
  OR2X1 P1_add_348_U143 ( .IN2(P1_N5169), .IN1(P1_add_348_n137), 
        .Q(P1_add_348_n136) );
  NAND2X0 P1_add_348_U142 ( .IN1(P1_N1632), .IN2(P1_add_348_n136), 
        .QN(P1_add_348_n135) );
  NAND2X0 P1_add_348_U141 ( .IN1(P1_add_348_n134), .IN2(P1_add_348_n135), 
        .QN(P1_add_348_n127) );
  OR2X1 P1_add_348_U139 ( .IN2(P1_N1633), .IN1(n7092), .Q(P1_add_348_n131) );
  NAND2X0 P1_add_348_U138 ( .IN1(P1_N1633), .IN2(n7092), .QN(P1_add_348_n132)
         );
  NAND2X0 P1_add_348_U137 ( .IN1(P1_add_348_n131), .IN2(P1_add_348_n132), 
        .QN(P1_add_348_n130) );
  NOR2X0 P1_add_348_U136 ( .QN(P1_add_348_n128), .IN1(P1_add_348_n127), 
        .IN2(P1_add_348_n130) );
  AND2X1 P1_add_348_U135 ( .IN1(P1_add_348_n127), .IN2(P1_add_348_n130), 
        .Q(P1_add_348_n129) );
  NOR2X0 P1_add_348_U134 ( .QN(P1_N1875), .IN1(P1_add_348_n128), 
        .IN2(P1_add_348_n129) );
  NAND2X0 P1_add_348_U133 ( .IN1(P1_N5170), .IN2(P1_add_348_n127), 
        .QN(P1_add_348_n124) );
  OR2X1 P1_add_348_U132 ( .IN2(P1_N5170), .IN1(P1_add_348_n127), 
        .Q(P1_add_348_n126) );
  NAND2X0 P1_add_348_U131 ( .IN1(P1_N1633), .IN2(P1_add_348_n126), 
        .QN(P1_add_348_n125) );
  NAND2X0 P1_add_348_U130 ( .IN1(P1_add_348_n124), .IN2(P1_add_348_n125), 
        .QN(P1_add_348_n117) );
  OR2X1 P1_add_348_U128 ( .IN2(P1_N1634), .IN1(n7090), .Q(P1_add_348_n121) );
  NAND2X0 P1_add_348_U127 ( .IN1(P1_N1634), .IN2(n7090), .QN(P1_add_348_n122)
         );
  NAND2X0 P1_add_348_U126 ( .IN1(P1_add_348_n121), .IN2(P1_add_348_n122), 
        .QN(P1_add_348_n120) );
  NOR2X0 P1_add_348_U125 ( .QN(P1_add_348_n118), .IN1(P1_add_348_n117), 
        .IN2(P1_add_348_n120) );
  AND2X1 P1_add_348_U124 ( .IN1(P1_add_348_n117), .IN2(P1_add_348_n120), 
        .Q(P1_add_348_n119) );
  NOR2X0 P1_add_348_U123 ( .QN(P1_N1876), .IN1(P1_add_348_n118), 
        .IN2(P1_add_348_n119) );
  NAND2X0 P1_add_348_U122 ( .IN1(P1_N5171), .IN2(P1_add_348_n117), 
        .QN(P1_add_348_n114) );
  OR2X1 P1_add_348_U121 ( .IN2(P1_N5171), .IN1(P1_add_348_n117), 
        .Q(P1_add_348_n116) );
  NAND2X0 P1_add_348_U120 ( .IN1(P1_N1634), .IN2(P1_add_348_n116), 
        .QN(P1_add_348_n115) );
  NAND2X0 P1_add_348_U119 ( .IN1(P1_add_348_n114), .IN2(P1_add_348_n115), 
        .QN(P1_add_348_n107) );
  OR2X1 P1_add_348_U117 ( .IN2(P1_N1635), .IN1(n7144), .Q(P1_add_348_n111) );
  NAND2X0 P1_add_348_U116 ( .IN1(P1_N1635), .IN2(n7144), .QN(P1_add_348_n112)
         );
  NAND2X0 P1_add_348_U115 ( .IN1(P1_add_348_n111), .IN2(P1_add_348_n112), 
        .QN(P1_add_348_n110) );
  NOR2X0 P1_add_348_U114 ( .QN(P1_add_348_n108), .IN1(P1_add_348_n107), 
        .IN2(P1_add_348_n110) );
  AND2X1 P1_add_348_U113 ( .IN1(P1_add_348_n107), .IN2(P1_add_348_n110), 
        .Q(P1_add_348_n109) );
  NOR2X0 P1_add_348_U112 ( .QN(P1_N1877), .IN1(P1_add_348_n108), 
        .IN2(P1_add_348_n109) );
  NAND2X0 P1_add_348_U111 ( .IN1(P1_N5172), .IN2(P1_add_348_n107), 
        .QN(P1_add_348_n104) );
  OR2X1 P1_add_348_U110 ( .IN2(P1_N5172), .IN1(P1_add_348_n107), 
        .Q(P1_add_348_n106) );
  NAND2X0 P1_add_348_U109 ( .IN1(P1_N1635), .IN2(P1_add_348_n106), 
        .QN(P1_add_348_n105) );
  NAND2X0 P1_add_348_U108 ( .IN1(P1_add_348_n104), .IN2(P1_add_348_n105), 
        .QN(P1_add_348_n97) );
  OR2X1 P1_add_348_U106 ( .IN2(P1_N1636), .IN1(n7136), .Q(P1_add_348_n101) );
  NAND2X0 P1_add_348_U105 ( .IN1(P1_N1636), .IN2(n7136), .QN(P1_add_348_n102)
         );
  NAND2X0 P1_add_348_U104 ( .IN1(P1_add_348_n101), .IN2(P1_add_348_n102), 
        .QN(P1_add_348_n100) );
  NOR2X0 P1_add_348_U103 ( .QN(P1_add_348_n98), .IN1(P1_add_348_n97), 
        .IN2(P1_add_348_n100) );
  AND2X1 P1_add_348_U102 ( .IN1(P1_add_348_n97), .IN2(P1_add_348_n100), 
        .Q(P1_add_348_n99) );
  NOR2X0 P1_add_348_U101 ( .QN(P1_N1878), .IN1(P1_add_348_n98), 
        .IN2(P1_add_348_n99) );
  NAND2X0 P1_add_348_U100 ( .IN1(n7138), .IN2(P1_add_348_n97), 
        .QN(P1_add_348_n94) );
  OR2X1 P1_add_348_U99 ( .IN2(n7138), .IN1(P1_add_348_n97), .Q(P1_add_348_n96)
         );
  NAND2X0 P1_add_348_U98 ( .IN1(P1_N1636), .IN2(P1_add_348_n96), 
        .QN(P1_add_348_n95) );
  NAND2X0 P1_add_348_U97 ( .IN1(P1_add_348_n94), .IN2(P1_add_348_n95), 
        .QN(P1_add_348_n87) );
  OR2X1 P1_add_348_U95 ( .IN2(P1_N1637), .IN1(n7130), .Q(P1_add_348_n91) );
  NAND2X0 P1_add_348_U94 ( .IN1(P1_N1637), .IN2(n7130), .QN(P1_add_348_n92) );
  NAND2X0 P1_add_348_U93 ( .IN1(P1_add_348_n91), .IN2(P1_add_348_n92), 
        .QN(P1_add_348_n90) );
  NOR2X0 P1_add_348_U92 ( .QN(P1_add_348_n88), .IN1(P1_add_348_n87), 
        .IN2(P1_add_348_n90) );
  AND2X1 P1_add_348_U91 ( .IN1(P1_add_348_n87), .IN2(P1_add_348_n90), 
        .Q(P1_add_348_n89) );
  NOR2X0 P1_add_348_U90 ( .QN(P1_N1879), .IN1(P1_add_348_n88), 
        .IN2(P1_add_348_n89) );
  NAND2X0 P1_add_348_U89 ( .IN1(n7129), .IN2(P1_add_348_n87), 
        .QN(P1_add_348_n84) );
  OR2X1 P1_add_348_U88 ( .IN2(n7129), .IN1(P1_add_348_n87), .Q(P1_add_348_n86)
         );
  NAND2X0 P1_add_348_U87 ( .IN1(P1_N1637), .IN2(P1_add_348_n86), 
        .QN(P1_add_348_n85) );
  NAND2X0 P1_add_348_U86 ( .IN1(P1_add_348_n84), .IN2(P1_add_348_n85), 
        .QN(P1_add_348_n77) );
  OR2X1 P1_add_348_U84 ( .IN2(P1_N1638), .IN1(n7125), .Q(P1_add_348_n81) );
  NAND2X0 P1_add_348_U83 ( .IN1(P1_N1638), .IN2(n7125), .QN(P1_add_348_n82) );
  NAND2X0 P1_add_348_U82 ( .IN1(P1_add_348_n81), .IN2(P1_add_348_n82), 
        .QN(P1_add_348_n80) );
  NOR2X0 P1_add_348_U81 ( .QN(P1_add_348_n78), .IN1(P1_add_348_n77), 
        .IN2(P1_add_348_n80) );
  AND2X1 P1_add_348_U80 ( .IN1(P1_add_348_n77), .IN2(P1_add_348_n80), 
        .Q(P1_add_348_n79) );
  NOR2X0 P1_add_348_U79 ( .QN(P1_N1880), .IN1(P1_add_348_n78), 
        .IN2(P1_add_348_n79) );
  NAND2X0 P1_add_348_U78 ( .IN1(n7124), .IN2(P1_add_348_n77), 
        .QN(P1_add_348_n74) );
  OR2X1 P1_add_348_U77 ( .IN2(n7124), .IN1(P1_add_348_n77), .Q(P1_add_348_n76)
         );
  NAND2X0 P1_add_348_U76 ( .IN1(P1_N1638), .IN2(P1_add_348_n76), 
        .QN(P1_add_348_n75) );
  NAND2X0 P1_add_348_U75 ( .IN1(P1_add_348_n74), .IN2(P1_add_348_n75), 
        .QN(P1_add_348_n64) );
  OR2X1 P1_add_348_U73 ( .IN2(P1_N1639), .IN1(n7119), .Q(P1_add_348_n71) );
  NAND2X0 P1_add_348_U72 ( .IN1(P1_N1639), .IN2(n7119), .QN(P1_add_348_n72) );
  NAND2X0 P1_add_348_U71 ( .IN1(P1_add_348_n71), .IN2(P1_add_348_n72), 
        .QN(P1_add_348_n70) );
  NOR2X0 P1_add_348_U70 ( .QN(P1_add_348_n68), .IN1(P1_add_348_n64), 
        .IN2(P1_add_348_n70) );
  AND2X1 P1_add_348_U69 ( .IN1(P1_add_348_n64), .IN2(P1_add_348_n70), 
        .Q(P1_add_348_n69) );
  NOR2X0 P1_add_348_U68 ( .QN(P1_N1881), .IN1(P1_add_348_n68), 
        .IN2(P1_add_348_n69) );
  OR2X1 P1_add_348_U66 ( .IN2(P1_N1640), .IN1(n7117), .Q(P1_add_348_n65) );
  NAND2X0 P1_add_348_U65 ( .IN1(P1_N1640), .IN2(n7117), .QN(P1_add_348_n66) );
  NAND2X0 P1_add_348_U64 ( .IN1(P1_add_348_n65), .IN2(P1_add_348_n66), 
        .QN(P1_add_348_n60) );
  NAND2X0 P1_add_348_U63 ( .IN1(P1_N5176), .IN2(P1_add_348_n64), 
        .QN(P1_add_348_n61) );
  OR2X1 P1_add_348_U62 ( .IN2(P1_N5176), .IN1(P1_add_348_n64), 
        .Q(P1_add_348_n63) );
  NAND2X0 P1_add_348_U61 ( .IN1(P1_N1639), .IN2(P1_add_348_n63), 
        .QN(P1_add_348_n62) );
  NAND2X0 P1_add_348_U60 ( .IN1(P1_add_348_n61), .IN2(P1_add_348_n62), 
        .QN(P1_add_348_n59) );
  OR2X1 P1_add_348_U244 ( .IN2(P1_N1624), .IN1(P1_add_348_n93), 
        .Q(P1_add_348_n228) );
  NAND2X0 P1_add_348_U243 ( .IN1(P1_N1624), .IN2(P1_add_348_n93), 
        .QN(P1_add_348_n229) );
  NAND2X0 P1_add_348_U242 ( .IN1(P1_add_348_n228), .IN2(P1_add_348_n229), 
        .QN(P1_add_348_n227) );
  NOR2X0 P1_add_348_U241 ( .QN(P1_add_348_n225), .IN1(P1_add_348_n224), 
        .IN2(P1_add_348_n227) );
  AND2X1 P1_add_348_U240 ( .IN1(P1_add_348_n224), .IN2(P1_add_348_n227), 
        .Q(P1_add_348_n226) );
  NOR2X0 P1_add_348_U239 ( .QN(P1_N1866), .IN1(P1_add_348_n225), 
        .IN2(P1_add_348_n226) );
  NAND2X0 P1_add_348_U238 ( .IN1(n7059), .IN2(P1_add_348_n224), 
        .QN(P1_add_348_n221) );
  OR2X1 P1_add_348_U237 ( .IN2(n7059), .IN1(P1_add_348_n224), 
        .Q(P1_add_348_n223) );
  NAND2X0 P1_add_348_U236 ( .IN1(P1_N1624), .IN2(P1_add_348_n223), 
        .QN(P1_add_348_n222) );
  NAND2X0 P1_add_348_U235 ( .IN1(P1_add_348_n221), .IN2(P1_add_348_n222), 
        .QN(P1_add_348_n214) );
  OR2X1 P1_add_348_U233 ( .IN2(P1_N1625), .IN1(n7056), .Q(P1_add_348_n218) );
  NAND2X0 P1_add_348_U232 ( .IN1(P1_N1625), .IN2(n7056), .QN(P1_add_348_n219)
         );
  NAND2X0 P1_add_348_U231 ( .IN1(P1_add_348_n218), .IN2(P1_add_348_n219), 
        .QN(P1_add_348_n217) );
  NOR2X0 P1_add_348_U230 ( .QN(P1_add_348_n215), .IN1(P1_add_348_n214), 
        .IN2(P1_add_348_n217) );
  AND2X1 P1_add_348_U229 ( .IN1(P1_add_348_n214), .IN2(P1_add_348_n217), 
        .Q(P1_add_348_n216) );
  NOR2X0 P1_add_348_U228 ( .QN(P1_N1867), .IN1(P1_add_348_n215), 
        .IN2(P1_add_348_n216) );
  NAND2X0 P1_add_348_U227 ( .IN1(n7055), .IN2(P1_add_348_n214), 
        .QN(P1_add_348_n211) );
  OR2X1 P1_add_348_U226 ( .IN2(n7055), .IN1(P1_add_348_n214), 
        .Q(P1_add_348_n213) );
  NAND2X0 P1_add_348_U225 ( .IN1(P1_N1625), .IN2(P1_add_348_n213), 
        .QN(P1_add_348_n212) );
  NAND2X0 P1_add_348_U224 ( .IN1(P1_add_348_n211), .IN2(P1_add_348_n212), 
        .QN(P1_add_348_n204) );
  OR2X1 P1_add_348_U222 ( .IN2(P1_N1626), .IN1(n7115), .Q(P1_add_348_n208) );
  NAND2X0 P1_add_348_U221 ( .IN1(P1_N1626), .IN2(n7115), .QN(P1_add_348_n209)
         );
  NAND2X0 P1_add_348_U220 ( .IN1(P1_add_348_n208), .IN2(P1_add_348_n209), 
        .QN(P1_add_348_n207) );
  NOR2X0 P1_add_348_U219 ( .QN(P1_add_348_n205), .IN1(P1_add_348_n204), 
        .IN2(P1_add_348_n207) );
  AND2X1 P1_add_348_U218 ( .IN1(P1_add_348_n204), .IN2(P1_add_348_n207), 
        .Q(P1_add_348_n206) );
  NOR2X0 P1_add_348_U217 ( .QN(P1_N1868), .IN1(P1_add_348_n205), 
        .IN2(P1_add_348_n206) );
  NAND2X0 P1_add_348_U216 ( .IN1(n7116), .IN2(P1_add_348_n204), 
        .QN(P1_add_348_n201) );
  OR2X1 P1_add_348_U215 ( .IN2(n7116), .IN1(P1_add_348_n204), 
        .Q(P1_add_348_n203) );
  NAND2X0 P1_add_348_U214 ( .IN1(P1_N1626), .IN2(P1_add_348_n203), 
        .QN(P1_add_348_n202) );
  NAND2X0 P1_add_348_U213 ( .IN1(P1_add_348_n201), .IN2(P1_add_348_n202), 
        .QN(P1_add_348_n194) );
  OR2X1 P1_add_348_U211 ( .IN2(P1_N1627), .IN1(n7112), .Q(P1_add_348_n198) );
  NAND2X0 P1_add_348_U210 ( .IN1(P1_N1627), .IN2(n7112), .QN(P1_add_348_n199)
         );
  NAND2X0 P1_add_348_U209 ( .IN1(P1_add_348_n198), .IN2(P1_add_348_n199), 
        .QN(P1_add_348_n197) );
  NOR2X0 P1_add_348_U208 ( .QN(P1_add_348_n195), .IN1(P1_add_348_n194), 
        .IN2(P1_add_348_n197) );
  AND2X1 P1_add_348_U207 ( .IN1(P1_add_348_n194), .IN2(P1_add_348_n197), 
        .Q(P1_add_348_n196) );
  NOR2X0 P1_add_348_U206 ( .QN(P1_N1869), .IN1(P1_add_348_n195), 
        .IN2(P1_add_348_n196) );
  NAND2X0 P1_add_348_U205 ( .IN1(P1_N5164), .IN2(P1_add_348_n194), 
        .QN(P1_add_348_n191) );
  OR2X1 P1_add_348_U204 ( .IN2(P1_N5164), .IN1(P1_add_348_n194), 
        .Q(P1_add_348_n193) );
  NAND2X0 P1_add_348_U203 ( .IN1(P1_N1627), .IN2(P1_add_348_n193), 
        .QN(P1_add_348_n192) );
  NAND2X0 P1_add_348_U202 ( .IN1(P1_add_348_n191), .IN2(P1_add_348_n192), 
        .QN(P1_add_348_n184) );
  OR2X1 P1_add_348_U200 ( .IN2(P1_N1628), .IN1(n7109), .Q(P1_add_348_n188) );
  NAND2X0 P1_add_348_U199 ( .IN1(P1_N1628), .IN2(n7109), .QN(P1_add_348_n189)
         );
  NAND2X0 P1_add_348_U198 ( .IN1(P1_add_348_n188), .IN2(P1_add_348_n189), 
        .QN(P1_add_348_n187) );
  NOR2X0 P1_add_348_U197 ( .QN(P1_add_348_n185), .IN1(P1_add_348_n184), 
        .IN2(P1_add_348_n187) );
  AND2X1 P1_add_348_U196 ( .IN1(P1_add_348_n184), .IN2(P1_add_348_n187), 
        .Q(P1_add_348_n186) );
  NOR2X0 P1_add_348_U195 ( .QN(P1_N1870), .IN1(P1_add_348_n185), 
        .IN2(P1_add_348_n186) );
  NAND2X0 P1_add_348_U194 ( .IN1(P1_N5165), .IN2(P1_add_348_n184), 
        .QN(P1_add_348_n181) );
  OR2X1 P1_add_348_U193 ( .IN2(P1_N5165), .IN1(P1_add_348_n184), 
        .Q(P1_add_348_n183) );
  NAND2X0 P1_add_348_U192 ( .IN1(P1_N1628), .IN2(P1_add_348_n183), 
        .QN(P1_add_348_n182) );
  NAND2X0 P1_add_348_U191 ( .IN1(P1_add_348_n181), .IN2(P1_add_348_n182), 
        .QN(P1_add_348_n174) );
  OR2X1 P1_add_348_U189 ( .IN2(P1_N1629), .IN1(n7105), .Q(P1_add_348_n178) );
  NAND2X0 P1_add_348_U188 ( .IN1(P1_N1629), .IN2(n7105), .QN(P1_add_348_n179)
         );
  NAND2X0 P1_add_348_U187 ( .IN1(P1_add_348_n178), .IN2(P1_add_348_n179), 
        .QN(P1_add_348_n177) );
  NOR2X0 P1_add_348_U186 ( .QN(P1_add_348_n175), .IN1(P1_add_348_n174), 
        .IN2(P1_add_348_n177) );
  AND2X1 P1_add_348_U185 ( .IN1(P1_add_348_n174), .IN2(P1_add_348_n177), 
        .Q(P1_add_348_n176) );
  NOR2X0 P1_add_348_U184 ( .QN(P1_N1871), .IN1(P1_add_348_n175), 
        .IN2(P1_add_348_n176) );
  NAND2X0 P1_add_348_U183 ( .IN1(n7106), .IN2(P1_add_348_n174), 
        .QN(P1_add_348_n171) );
  OR2X1 P1_add_348_U182 ( .IN2(n7106), .IN1(P1_add_348_n174), 
        .Q(P1_add_348_n173) );
  NAND2X0 P1_add_348_U181 ( .IN1(P1_N1629), .IN2(P1_add_348_n173), 
        .QN(P1_add_348_n172) );
  NAND2X0 P1_add_348_U180 ( .IN1(P1_add_348_n171), .IN2(P1_add_348_n172), 
        .QN(P1_add_348_n164) );
  OR2X1 P1_add_348_U178 ( .IN2(P1_N1630), .IN1(n7102), .Q(P1_add_348_n168) );
  NAND2X0 P1_add_348_U177 ( .IN1(P1_N1630), .IN2(n7102), .QN(P1_add_348_n169)
         );
  NAND2X0 P1_add_348_U176 ( .IN1(P1_add_348_n168), .IN2(P1_add_348_n169), 
        .QN(P1_add_348_n167) );
  NOR2X0 P1_add_348_U175 ( .QN(P1_add_348_n165), .IN1(P1_add_348_n164), 
        .IN2(P1_add_348_n167) );
  AND2X1 P1_add_348_U174 ( .IN1(P1_add_348_n164), .IN2(P1_add_348_n167), 
        .Q(P1_add_348_n166) );
  NOR2X0 P1_add_348_U173 ( .QN(P1_N1872), .IN1(P1_add_348_n165), 
        .IN2(P1_add_348_n166) );
  NAND2X0 P1_add_348_U172 ( .IN1(P1_N5167), .IN2(P1_add_348_n164), 
        .QN(P1_add_348_n161) );
  OR2X1 P1_add_348_U171 ( .IN2(P1_N5167), .IN1(P1_add_348_n164), 
        .Q(P1_add_348_n163) );
  NAND2X0 P1_add_348_U170 ( .IN1(P1_N1630), .IN2(P1_add_348_n163), 
        .QN(P1_add_348_n162) );
  NAND2X0 P1_add_348_U169 ( .IN1(P1_add_348_n161), .IN2(P1_add_348_n162), 
        .QN(P1_add_348_n147) );
  OR2X1 P1_add_348_U167 ( .IN2(P1_N1631), .IN1(n7098), .Q(P1_add_348_n158) );
  NAND2X0 P1_add_348_U166 ( .IN1(P1_N1631), .IN2(n7098), .QN(P1_add_348_n159)
         );
  NAND2X0 P1_add_348_U165 ( .IN1(P1_add_348_n158), .IN2(P1_add_348_n159), 
        .QN(P1_add_348_n157) );
  NOR2X0 P1_add_348_U164 ( .QN(P1_add_348_n155), .IN1(P1_add_348_n147), 
        .IN2(P1_add_348_n157) );
  AND2X1 P1_add_348_U163 ( .IN1(P1_add_348_n147), .IN2(P1_add_348_n157), 
        .Q(P1_add_348_n156) );
  NOR2X0 P1_add_348_U162 ( .QN(P1_N1873), .IN1(P1_add_348_n155), 
        .IN2(P1_add_348_n156) );
  OR2X1 P1_add_348_U161 ( .IN2(P1_N1613), .IN1(n7051), .Q(P1_add_348_n152) );
  NAND2X0 P1_add_348_U160 ( .IN1(P1_N1613), .IN2(n7051), .QN(P1_add_348_n153)
         );
  NAND2X0 P1_add_348_U159 ( .IN1(P1_add_348_n152), .IN2(P1_add_348_n153), 
        .QN(P1_add_348_n150) );
  NAND2X0 P1_add_348_U158 ( .IN1(P1_add_348_n150), .IN2(P1_add_348_n151), 
        .QN(P1_add_348_n148) );
  OR2X1 P1_add_348_U157 ( .IN2(P1_add_348_n151), .IN1(P1_add_348_n150), 
        .Q(P1_add_348_n149) );
  NAND2X0 P1_add_348_U156 ( .IN1(P1_add_348_n148), .IN2(P1_add_348_n149), 
        .QN(P1_N1855) );
  NAND2X0 P1_add_348_U155 ( .IN1(n7099), .IN2(P1_add_348_n147), 
        .QN(P1_add_348_n144) );
  OR2X1 P1_add_348_U154 ( .IN2(n7099), .IN1(P1_add_348_n147), 
        .Q(P1_add_348_n146) );
  NAND2X0 P1_add_348_U153 ( .IN1(P1_N1631), .IN2(P1_add_348_n146), 
        .QN(P1_add_348_n145) );
  OR2X1 P1_add_348_U308 ( .IN2(P1_N1612), .IN1(n4803), .Q(P1_add_348_n278) );
  NAND2X0 P1_add_348_U307 ( .IN1(P1_N1612), .IN2(n4803), .QN(P1_add_348_n279)
         );
  NAND2X0 P1_add_348_U306 ( .IN1(P1_add_348_n278), .IN2(P1_add_348_n279), 
        .QN(P1_N1854) );
  NAND2X0 P1_add_348_U304 ( .IN1(P1_N1612), .IN2(n7034), .QN(P1_add_348_n151)
         );
  OR2X1 P1_add_348_U303 ( .IN2(P1_add_348_n151), .IN1(n7051), 
        .Q(P1_add_348_n275) );
  NAND2X0 P1_add_348_U302 ( .IN1(n7051), .IN2(P1_add_348_n151), 
        .QN(P1_add_348_n277) );
  NAND2X0 P1_add_348_U301 ( .IN1(P1_N1613), .IN2(P1_add_348_n277), 
        .QN(P1_add_348_n276) );
  NAND2X0 P1_add_348_U300 ( .IN1(P1_add_348_n275), .IN2(P1_add_348_n276), 
        .QN(P1_add_348_n52) );
  NAND2X0 P1_add_348_U299 ( .IN1(n7046), .IN2(P1_add_348_n52), 
        .QN(P1_add_348_n272) );
  OR2X1 P1_add_348_U298 ( .IN2(n7046), .IN1(P1_add_348_n52), 
        .Q(P1_add_348_n274) );
  NAND2X0 P1_add_348_U297 ( .IN1(P1_N1614), .IN2(P1_add_348_n274), 
        .QN(P1_add_348_n273) );
  NAND2X0 P1_add_348_U296 ( .IN1(P1_add_348_n272), .IN2(P1_add_348_n273), 
        .QN(P1_add_348_n45) );
  NAND2X0 P1_add_348_U295 ( .IN1(n7041), .IN2(P1_add_348_n45), 
        .QN(P1_add_348_n269) );
  OR2X1 P1_add_348_U294 ( .IN2(n7041), .IN1(P1_add_348_n45), 
        .Q(P1_add_348_n271) );
  NAND2X0 P1_add_348_U293 ( .IN1(P1_N1615), .IN2(P1_add_348_n271), 
        .QN(P1_add_348_n270) );
  NAND2X0 P1_add_348_U292 ( .IN1(P1_add_348_n269), .IN2(P1_add_348_n270), 
        .QN(P1_add_348_n38) );
  NAND2X0 P1_add_348_U291 ( .IN1(n7036), .IN2(P1_add_348_n38), 
        .QN(P1_add_348_n266) );
  OR2X1 P1_add_348_U290 ( .IN2(n7036), .IN1(P1_add_348_n38), 
        .Q(P1_add_348_n268) );
  NAND2X0 P1_add_348_U289 ( .IN1(P1_N1616), .IN2(P1_add_348_n268), 
        .QN(P1_add_348_n267) );
  NAND2X0 P1_add_348_U288 ( .IN1(P1_add_348_n266), .IN2(P1_add_348_n267), 
        .QN(P1_add_348_n31) );
  NAND2X0 P1_add_348_U287 ( .IN1(n7081), .IN2(P1_add_348_n31), 
        .QN(P1_add_348_n263) );
  OR2X1 P1_add_348_U286 ( .IN2(n7081), .IN1(P1_add_348_n31), 
        .Q(P1_add_348_n265) );
  NAND2X0 P1_add_348_U285 ( .IN1(P1_N1617), .IN2(P1_add_348_n265), 
        .QN(P1_add_348_n264) );
  NAND2X0 P1_add_348_U284 ( .IN1(P1_add_348_n263), .IN2(P1_add_348_n264), 
        .QN(P1_add_348_n24) );
  NAND2X0 P1_add_348_U283 ( .IN1(P1_N5155), .IN2(P1_add_348_n24), 
        .QN(P1_add_348_n260) );
  OR2X1 P1_add_348_U282 ( .IN2(P1_N5155), .IN1(P1_add_348_n24), 
        .Q(P1_add_348_n262) );
  NAND2X0 P1_add_348_U281 ( .IN1(P1_N1618), .IN2(P1_add_348_n262), 
        .QN(P1_add_348_n261) );
  NAND2X0 P1_add_348_U280 ( .IN1(P1_add_348_n260), .IN2(P1_add_348_n261), 
        .QN(P1_add_348_n17) );
  NAND2X0 P1_add_348_U279 ( .IN1(n7075), .IN2(P1_add_348_n17), 
        .QN(P1_add_348_n257) );
  OR2X1 P1_add_348_U278 ( .IN2(n7075), .IN1(P1_add_348_n17), 
        .Q(P1_add_348_n259) );
  NAND2X0 P1_add_348_U277 ( .IN1(P1_N1619), .IN2(P1_add_348_n259), 
        .QN(P1_add_348_n258) );
  NAND2X0 P1_add_348_U276 ( .IN1(P1_add_348_n257), .IN2(P1_add_348_n258), 
        .QN(P1_add_348_n10) );
  NAND2X0 P1_add_348_U275 ( .IN1(n7072), .IN2(P1_add_348_n10), 
        .QN(P1_add_348_n254) );
  OR2X1 P1_add_348_U274 ( .IN2(n7072), .IN1(P1_add_348_n10), 
        .Q(P1_add_348_n256) );
  NAND2X0 P1_add_348_U273 ( .IN1(P1_N1620), .IN2(P1_add_348_n256), 
        .QN(P1_add_348_n255) );
  NAND2X0 P1_add_348_U272 ( .IN1(P1_add_348_n254), .IN2(P1_add_348_n255), 
        .QN(P1_add_348_n3) );
  NAND2X0 P1_add_348_U271 ( .IN1(n7070), .IN2(P1_add_348_n3), 
        .QN(P1_add_348_n251) );
  OR2X1 P1_add_348_U270 ( .IN2(P1_N5158), .IN1(P1_add_348_n3), 
        .Q(P1_add_348_n253) );
  NAND2X0 P1_add_348_U269 ( .IN1(P1_N1621), .IN2(P1_add_348_n253), 
        .QN(P1_add_348_n252) );
  NAND2X0 P1_add_348_U268 ( .IN1(P1_add_348_n251), .IN2(P1_add_348_n252), 
        .QN(P1_add_348_n244) );
  OR2X1 P1_add_348_U266 ( .IN2(P1_N1622), .IN1(n7067), .Q(P1_add_348_n248) );
  NAND2X0 P1_add_348_U265 ( .IN1(P1_N1622), .IN2(n7067), .QN(P1_add_348_n249)
         );
  NAND2X0 P1_add_348_U264 ( .IN1(P1_add_348_n248), .IN2(P1_add_348_n249), 
        .QN(P1_add_348_n247) );
  NOR2X0 P1_add_348_U263 ( .QN(P1_add_348_n245), .IN1(P1_add_348_n244), 
        .IN2(P1_add_348_n247) );
  AND2X1 P1_add_348_U262 ( .IN1(P1_add_348_n244), .IN2(P1_add_348_n247), 
        .Q(P1_add_348_n246) );
  NOR2X0 P1_add_348_U261 ( .QN(P1_N1864), .IN1(P1_add_348_n245), 
        .IN2(P1_add_348_n246) );
  NAND2X0 P1_add_348_U260 ( .IN1(n7066), .IN2(P1_add_348_n244), 
        .QN(P1_add_348_n241) );
  OR2X1 P1_add_348_U259 ( .IN2(n7066), .IN1(P1_add_348_n244), 
        .Q(P1_add_348_n243) );
  NAND2X0 P1_add_348_U258 ( .IN1(P1_N1622), .IN2(P1_add_348_n243), 
        .QN(P1_add_348_n242) );
  NAND2X0 P1_add_348_U257 ( .IN1(P1_add_348_n241), .IN2(P1_add_348_n242), 
        .QN(P1_add_348_n234) );
  OR2X1 P1_add_348_U255 ( .IN2(P1_N1623), .IN1(n7063), .Q(P1_add_348_n238) );
  NAND2X0 P1_add_348_U254 ( .IN1(P1_N1623), .IN2(n7063), .QN(P1_add_348_n239)
         );
  NAND2X0 P1_add_348_U253 ( .IN1(P1_add_348_n238), .IN2(P1_add_348_n239), 
        .QN(P1_add_348_n237) );
  NOR2X0 P1_add_348_U252 ( .QN(P1_add_348_n235), .IN1(P1_add_348_n234), 
        .IN2(P1_add_348_n237) );
  AND2X1 P1_add_348_U251 ( .IN1(P1_add_348_n234), .IN2(P1_add_348_n237), 
        .Q(P1_add_348_n236) );
  NOR2X0 P1_add_348_U250 ( .QN(P1_N1865), .IN1(P1_add_348_n235), 
        .IN2(P1_add_348_n236) );
  NAND2X0 P1_add_348_U249 ( .IN1(n7062), .IN2(P1_add_348_n234), 
        .QN(P1_add_348_n231) );
  OR2X1 P1_add_348_U248 ( .IN2(n7062), .IN1(P1_add_348_n234), 
        .Q(P1_add_348_n233) );
  NAND2X0 P1_add_348_U247 ( .IN1(P1_N1623), .IN2(P1_add_348_n233), 
        .QN(P1_add_348_n232) );
  NAND2X0 P1_add_348_U246 ( .IN1(P1_add_348_n231), .IN2(P1_add_348_n232), 
        .QN(P1_add_348_n224) );
  INVX0 P1_add_348_U7 ( .ZN(P1_add_348_n93), .INP(n7059) );
  INVX0 P1_add_348_U14 ( .ZN(P1_add_348_n180), .INP(n7072) );
  NAND2X0 P1_add_368_U89 ( .IN1(n7129), .IN2(P1_add_368_n87), 
        .QN(P1_add_368_n84) );
  OR2X1 P1_add_368_U88 ( .IN2(n7129), .IN1(P1_add_368_n87), .Q(P1_add_368_n86)
         );
  NAND2X0 P1_add_368_U87 ( .IN1(P1_N2010), .IN2(P1_add_368_n86), 
        .QN(P1_add_368_n85) );
  NAND2X0 P1_add_368_U86 ( .IN1(P1_add_368_n84), .IN2(P1_add_368_n85), 
        .QN(P1_add_368_n77) );
  OR2X1 P1_add_368_U84 ( .IN2(P1_N2011), .IN1(n7125), .Q(P1_add_368_n81) );
  NAND2X0 P1_add_368_U83 ( .IN1(P1_N2011), .IN2(n7125), .QN(P1_add_368_n82) );
  NAND2X0 P1_add_368_U82 ( .IN1(P1_add_368_n81), .IN2(P1_add_368_n82), 
        .QN(P1_add_368_n80) );
  NOR2X0 P1_add_368_U81 ( .QN(P1_add_368_n78), .IN1(P1_add_368_n77), 
        .IN2(P1_add_368_n80) );
  AND2X1 P1_add_368_U80 ( .IN1(P1_add_368_n77), .IN2(P1_add_368_n80), 
        .Q(P1_add_368_n79) );
  NOR2X0 P1_add_368_U79 ( .QN(P1_N2253), .IN1(P1_add_368_n78), 
        .IN2(P1_add_368_n79) );
  NAND2X0 P1_add_368_U78 ( .IN1(n7124), .IN2(P1_add_368_n77), 
        .QN(P1_add_368_n74) );
  OR2X1 P1_add_368_U77 ( .IN2(n7124), .IN1(P1_add_368_n77), .Q(P1_add_368_n76)
         );
  NAND2X0 P1_add_368_U76 ( .IN1(P1_N2011), .IN2(P1_add_368_n76), 
        .QN(P1_add_368_n75) );
  NAND2X0 P1_add_368_U75 ( .IN1(P1_add_368_n74), .IN2(P1_add_368_n75), 
        .QN(P1_add_368_n64) );
  OR2X1 P1_add_368_U73 ( .IN2(P1_N2012), .IN1(n7119), .Q(P1_add_368_n71) );
  NAND2X0 P1_add_368_U72 ( .IN1(P1_N2012), .IN2(n7119), .QN(P1_add_368_n72) );
  NAND2X0 P1_add_368_U71 ( .IN1(P1_add_368_n71), .IN2(P1_add_368_n72), 
        .QN(P1_add_368_n70) );
  NOR2X0 P1_add_368_U70 ( .QN(P1_add_368_n68), .IN1(P1_add_368_n64), 
        .IN2(P1_add_368_n70) );
  AND2X1 P1_add_368_U69 ( .IN1(P1_add_368_n64), .IN2(P1_add_368_n70), 
        .Q(P1_add_368_n69) );
  NOR2X0 P1_add_368_U68 ( .QN(P1_N2254), .IN1(P1_add_368_n68), 
        .IN2(P1_add_368_n69) );
  OR2X1 P1_add_368_U66 ( .IN2(P1_N2013), .IN1(n7117), .Q(P1_add_368_n65) );
  NAND2X0 P1_add_368_U65 ( .IN1(P1_N2013), .IN2(n7117), .QN(P1_add_368_n66) );
  NAND2X0 P1_add_368_U64 ( .IN1(P1_add_368_n65), .IN2(P1_add_368_n66), 
        .QN(P1_add_368_n60) );
  NAND2X0 P1_add_368_U63 ( .IN1(P1_N5176), .IN2(P1_add_368_n64), 
        .QN(P1_add_368_n61) );
  OR2X1 P1_add_368_U62 ( .IN2(P1_N5176), .IN1(P1_add_368_n64), 
        .Q(P1_add_368_n63) );
  NAND2X0 P1_add_368_U61 ( .IN1(P1_N2012), .IN2(P1_add_368_n63), 
        .QN(P1_add_368_n62) );
  NAND2X0 P1_add_368_U60 ( .IN1(P1_add_368_n61), .IN2(P1_add_368_n62), 
        .QN(P1_add_368_n59) );
  NOR2X0 P1_add_368_U59 ( .QN(P1_add_368_n57), .IN1(P1_add_368_n60), 
        .IN2(P1_add_368_n59) );
  AND2X1 P1_add_368_U58 ( .IN1(P1_add_368_n59), .IN2(P1_add_368_n60), 
        .Q(P1_add_368_n58) );
  NOR2X0 P1_add_368_U57 ( .QN(P1_N2255), .IN1(P1_add_368_n57), 
        .IN2(P1_add_368_n58) );
  OR2X1 P1_add_368_U55 ( .IN2(P1_N1987), .IN1(n7045), .Q(P1_add_368_n54) );
  NAND2X0 P1_add_368_U54 ( .IN1(P1_N1987), .IN2(n7045), .QN(P1_add_368_n55) );
  NAND2X0 P1_add_368_U53 ( .IN1(P1_add_368_n54), .IN2(P1_add_368_n55), 
        .QN(P1_add_368_n53) );
  NOR2X0 P1_add_368_U52 ( .QN(P1_add_368_n50), .IN1(P1_add_368_n52), 
        .IN2(P1_add_368_n53) );
  AND2X1 P1_add_368_U51 ( .IN1(P1_add_368_n52), .IN2(P1_add_368_n53), 
        .Q(P1_add_368_n51) );
  NOR2X0 P1_add_368_U50 ( .QN(P1_N2229), .IN1(P1_add_368_n50), 
        .IN2(P1_add_368_n51) );
  OR2X1 P1_add_368_U48 ( .IN2(P1_N1988), .IN1(n7043), .Q(P1_add_368_n47) );
  NAND2X0 P1_add_368_U47 ( .IN1(P1_N1988), .IN2(n7043), .QN(P1_add_368_n48) );
  NAND2X0 P1_add_368_U46 ( .IN1(P1_add_368_n47), .IN2(P1_add_368_n48), 
        .QN(P1_add_368_n46) );
  NOR2X0 P1_add_368_U45 ( .QN(P1_add_368_n43), .IN1(P1_add_368_n45), 
        .IN2(P1_add_368_n46) );
  AND2X1 P1_add_368_U44 ( .IN1(P1_add_368_n45), .IN2(P1_add_368_n46), 
        .Q(P1_add_368_n44) );
  NOR2X0 P1_add_368_U43 ( .QN(P1_N2230), .IN1(P1_add_368_n43), 
        .IN2(P1_add_368_n44) );
  OR2X1 P1_add_368_U41 ( .IN2(P1_N1989), .IN1(n7037), .Q(P1_add_368_n40) );
  NAND2X0 P1_add_368_U40 ( .IN1(P1_N1989), .IN2(n7037), .QN(P1_add_368_n41) );
  NAND2X0 P1_add_368_U39 ( .IN1(P1_add_368_n40), .IN2(P1_add_368_n41), 
        .QN(P1_add_368_n39) );
  NOR2X0 P1_add_368_U38 ( .QN(P1_add_368_n36), .IN1(P1_add_368_n38), 
        .IN2(P1_add_368_n39) );
  AND2X1 P1_add_368_U37 ( .IN1(P1_add_368_n38), .IN2(P1_add_368_n39), 
        .Q(P1_add_368_n37) );
  NOR2X0 P1_add_368_U36 ( .QN(P1_N2231), .IN1(P1_add_368_n36), 
        .IN2(P1_add_368_n37) );
  OR2X1 P1_add_368_U34 ( .IN2(P1_N1990), .IN1(n7082), .Q(P1_add_368_n33) );
  NAND2X0 P1_add_368_U33 ( .IN1(P1_N1990), .IN2(n7082), .QN(P1_add_368_n34) );
  NAND2X0 P1_add_368_U32 ( .IN1(P1_add_368_n33), .IN2(P1_add_368_n34), 
        .QN(P1_add_368_n32) );
  NOR2X0 P1_add_368_U31 ( .QN(P1_add_368_n29), .IN1(P1_add_368_n31), 
        .IN2(P1_add_368_n32) );
  AND2X1 P1_add_368_U30 ( .IN1(P1_add_368_n31), .IN2(P1_add_368_n32), 
        .Q(P1_add_368_n30) );
  NOR2X0 P1_add_368_U29 ( .QN(P1_N2232), .IN1(P1_add_368_n29), 
        .IN2(P1_add_368_n30) );
  OR2X1 P1_add_368_U27 ( .IN2(P1_N1991), .IN1(n7079), .Q(P1_add_368_n26) );
  NAND2X0 P1_add_368_U26 ( .IN1(P1_N1991), .IN2(n7079), .QN(P1_add_368_n27) );
  NAND2X0 P1_add_368_U25 ( .IN1(P1_add_368_n26), .IN2(P1_add_368_n27), 
        .QN(P1_add_368_n25) );
  NOR2X0 P1_add_368_U24 ( .QN(P1_add_368_n22), .IN1(P1_add_368_n24), 
        .IN2(P1_add_368_n25) );
  AND2X1 P1_add_368_U23 ( .IN1(P1_add_368_n24), .IN2(P1_add_368_n25), 
        .Q(P1_add_368_n23) );
  NOR2X0 P1_add_368_U22 ( .QN(P1_N2233), .IN1(P1_add_368_n22), 
        .IN2(P1_add_368_n23) );
  OR2X1 P1_add_368_U20 ( .IN2(P1_N1992), .IN1(n7076), .Q(P1_add_368_n19) );
  NAND2X0 P1_add_368_U19 ( .IN1(P1_N1992), .IN2(n7076), .QN(P1_add_368_n20) );
  NAND2X0 P1_add_368_U18 ( .IN1(P1_add_368_n19), .IN2(P1_add_368_n20), 
        .QN(P1_add_368_n18) );
  NOR2X0 P1_add_368_U17 ( .QN(P1_add_368_n15), .IN1(P1_add_368_n17), 
        .IN2(P1_add_368_n18) );
  AND2X1 P1_add_368_U16 ( .IN1(P1_add_368_n17), .IN2(P1_add_368_n18), 
        .Q(P1_add_368_n16) );
  NOR2X0 P1_add_368_U15 ( .QN(P1_N2234), .IN1(P1_add_368_n15), 
        .IN2(P1_add_368_n16) );
  OR2X1 P1_add_368_U13 ( .IN2(P1_N1993), .IN1(n7073), .Q(P1_add_368_n12) );
  NAND2X0 P1_add_368_U12 ( .IN1(P1_N1993), .IN2(n7073), .QN(P1_add_368_n13) );
  NAND2X0 P1_add_368_U11 ( .IN1(P1_add_368_n12), .IN2(P1_add_368_n13), 
        .QN(P1_add_368_n11) );
  NOR2X0 P1_add_368_U10 ( .QN(P1_add_368_n8), .IN1(P1_add_368_n10), 
        .IN2(P1_add_368_n11) );
  AND2X1 P1_add_368_U9 ( .IN1(P1_add_368_n10), .IN2(P1_add_368_n11), 
        .Q(P1_add_368_n9) );
  NOR2X0 P1_add_368_U8 ( .QN(P1_N2235), .IN1(P1_add_368_n8), 
        .IN2(P1_add_368_n9) );
  OR2X1 P1_add_368_U6 ( .IN2(P1_N1994), .IN1(n7071), .Q(P1_add_368_n5) );
  NAND2X0 P1_add_368_U5 ( .IN1(P1_N1994), .IN2(n7071), .QN(P1_add_368_n6) );
  NAND2X0 P1_add_368_U4 ( .IN1(P1_add_368_n5), .IN2(P1_add_368_n6), 
        .QN(P1_add_368_n4) );
  NOR2X0 P1_add_368_U3 ( .QN(P1_add_368_n1), .IN1(P1_add_368_n3), 
        .IN2(P1_add_368_n4) );
  AND2X1 P1_add_368_U2 ( .IN1(P1_add_368_n3), .IN2(P1_add_368_n4), 
        .Q(P1_add_368_n2) );
  NOR2X0 P1_add_368_U1 ( .QN(P1_N2236), .IN1(P1_add_368_n1), 
        .IN2(P1_add_368_n2) );
  OR2X1 P1_add_368_U182 ( .IN2(n7106), .IN1(P1_add_368_n174), 
        .Q(P1_add_368_n173) );
  NAND2X0 P1_add_368_U181 ( .IN1(P1_N2002), .IN2(P1_add_368_n173), 
        .QN(P1_add_368_n172) );
  NAND2X0 P1_add_368_U180 ( .IN1(P1_add_368_n171), .IN2(P1_add_368_n172), 
        .QN(P1_add_368_n164) );
  OR2X1 P1_add_368_U178 ( .IN2(P1_N2003), .IN1(n7102), .Q(P1_add_368_n168) );
  NAND2X0 P1_add_368_U177 ( .IN1(P1_N2003), .IN2(n7102), .QN(P1_add_368_n169)
         );
  NAND2X0 P1_add_368_U176 ( .IN1(P1_add_368_n168), .IN2(P1_add_368_n169), 
        .QN(P1_add_368_n167) );
  NOR2X0 P1_add_368_U175 ( .QN(P1_add_368_n165), .IN1(P1_add_368_n164), 
        .IN2(P1_add_368_n167) );
  AND2X1 P1_add_368_U174 ( .IN1(P1_add_368_n164), .IN2(P1_add_368_n167), 
        .Q(P1_add_368_n166) );
  NOR2X0 P1_add_368_U173 ( .QN(P1_N2245), .IN1(P1_add_368_n165), 
        .IN2(P1_add_368_n166) );
  NAND2X0 P1_add_368_U172 ( .IN1(P1_N5167), .IN2(P1_add_368_n164), 
        .QN(P1_add_368_n161) );
  OR2X1 P1_add_368_U171 ( .IN2(P1_N5167), .IN1(P1_add_368_n164), 
        .Q(P1_add_368_n163) );
  NAND2X0 P1_add_368_U170 ( .IN1(P1_N2003), .IN2(P1_add_368_n163), 
        .QN(P1_add_368_n162) );
  NAND2X0 P1_add_368_U169 ( .IN1(P1_add_368_n161), .IN2(P1_add_368_n162), 
        .QN(P1_add_368_n147) );
  OR2X1 P1_add_368_U167 ( .IN2(P1_N2004), .IN1(n7098), .Q(P1_add_368_n158) );
  NAND2X0 P1_add_368_U166 ( .IN1(P1_N2004), .IN2(n7098), .QN(P1_add_368_n159)
         );
  NAND2X0 P1_add_368_U165 ( .IN1(P1_add_368_n158), .IN2(P1_add_368_n159), 
        .QN(P1_add_368_n157) );
  NOR2X0 P1_add_368_U164 ( .QN(P1_add_368_n155), .IN1(P1_add_368_n147), 
        .IN2(P1_add_368_n157) );
  AND2X1 P1_add_368_U163 ( .IN1(P1_add_368_n147), .IN2(P1_add_368_n157), 
        .Q(P1_add_368_n156) );
  NOR2X0 P1_add_368_U162 ( .QN(P1_N2246), .IN1(P1_add_368_n155), 
        .IN2(P1_add_368_n156) );
  OR2X1 P1_add_368_U161 ( .IN2(P1_N1986), .IN1(n7048), .Q(P1_add_368_n152) );
  NAND2X0 P1_add_368_U160 ( .IN1(P1_N1986), .IN2(n7048), .QN(P1_add_368_n153)
         );
  NAND2X0 P1_add_368_U159 ( .IN1(P1_add_368_n152), .IN2(P1_add_368_n153), 
        .QN(P1_add_368_n150) );
  NAND2X0 P1_add_368_U158 ( .IN1(P1_add_368_n150), .IN2(P1_add_368_n151), 
        .QN(P1_add_368_n148) );
  OR2X1 P1_add_368_U157 ( .IN2(P1_add_368_n151), .IN1(P1_add_368_n150), 
        .Q(P1_add_368_n149) );
  NAND2X0 P1_add_368_U156 ( .IN1(P1_add_368_n148), .IN2(P1_add_368_n149), 
        .QN(P1_N2228) );
  NAND2X0 P1_add_368_U155 ( .IN1(P1_N5168), .IN2(P1_add_368_n147), 
        .QN(P1_add_368_n144) );
  OR2X1 P1_add_368_U154 ( .IN2(P1_N5168), .IN1(P1_add_368_n147), 
        .Q(P1_add_368_n146) );
  NAND2X0 P1_add_368_U153 ( .IN1(P1_N2004), .IN2(P1_add_368_n146), 
        .QN(P1_add_368_n145) );
  NAND2X0 P1_add_368_U152 ( .IN1(P1_add_368_n144), .IN2(P1_add_368_n145), 
        .QN(P1_add_368_n137) );
  OR2X1 P1_add_368_U150 ( .IN2(P1_N2005), .IN1(n7095), .Q(P1_add_368_n141) );
  NAND2X0 P1_add_368_U149 ( .IN1(P1_N2005), .IN2(n7095), .QN(P1_add_368_n142)
         );
  NAND2X0 P1_add_368_U148 ( .IN1(P1_add_368_n141), .IN2(P1_add_368_n142), 
        .QN(P1_add_368_n140) );
  NOR2X0 P1_add_368_U147 ( .QN(P1_add_368_n138), .IN1(P1_add_368_n137), 
        .IN2(P1_add_368_n140) );
  AND2X1 P1_add_368_U146 ( .IN1(P1_add_368_n137), .IN2(P1_add_368_n140), 
        .Q(P1_add_368_n139) );
  NOR2X0 P1_add_368_U145 ( .QN(P1_N2247), .IN1(P1_add_368_n138), 
        .IN2(P1_add_368_n139) );
  NAND2X0 P1_add_368_U144 ( .IN1(n7096), .IN2(P1_add_368_n137), 
        .QN(P1_add_368_n134) );
  OR2X1 P1_add_368_U143 ( .IN2(n7096), .IN1(P1_add_368_n137), 
        .Q(P1_add_368_n136) );
  NAND2X0 P1_add_368_U142 ( .IN1(P1_N2005), .IN2(P1_add_368_n136), 
        .QN(P1_add_368_n135) );
  NAND2X0 P1_add_368_U141 ( .IN1(P1_add_368_n134), .IN2(P1_add_368_n135), 
        .QN(P1_add_368_n127) );
  OR2X1 P1_add_368_U139 ( .IN2(P1_N2006), .IN1(n7092), .Q(P1_add_368_n131) );
  NAND2X0 P1_add_368_U138 ( .IN1(P1_N2006), .IN2(n7092), .QN(P1_add_368_n132)
         );
  NAND2X0 P1_add_368_U137 ( .IN1(P1_add_368_n131), .IN2(P1_add_368_n132), 
        .QN(P1_add_368_n130) );
  NOR2X0 P1_add_368_U136 ( .QN(P1_add_368_n128), .IN1(P1_add_368_n127), 
        .IN2(P1_add_368_n130) );
  AND2X1 P1_add_368_U135 ( .IN1(P1_add_368_n127), .IN2(P1_add_368_n130), 
        .Q(P1_add_368_n129) );
  NOR2X0 P1_add_368_U134 ( .QN(P1_N2248), .IN1(P1_add_368_n128), 
        .IN2(P1_add_368_n129) );
  NAND2X0 P1_add_368_U133 ( .IN1(n7093), .IN2(P1_add_368_n127), 
        .QN(P1_add_368_n124) );
  OR2X1 P1_add_368_U132 ( .IN2(P1_N5170), .IN1(P1_add_368_n127), 
        .Q(P1_add_368_n126) );
  NAND2X0 P1_add_368_U131 ( .IN1(P1_N2006), .IN2(P1_add_368_n126), 
        .QN(P1_add_368_n125) );
  NAND2X0 P1_add_368_U130 ( .IN1(P1_add_368_n124), .IN2(P1_add_368_n125), 
        .QN(P1_add_368_n117) );
  OR2X1 P1_add_368_U128 ( .IN2(P1_N2007), .IN1(n7090), .Q(P1_add_368_n121) );
  NAND2X0 P1_add_368_U127 ( .IN1(P1_N2007), .IN2(n7090), .QN(P1_add_368_n122)
         );
  NAND2X0 P1_add_368_U126 ( .IN1(P1_add_368_n121), .IN2(P1_add_368_n122), 
        .QN(P1_add_368_n120) );
  NOR2X0 P1_add_368_U125 ( .QN(P1_add_368_n118), .IN1(P1_add_368_n117), 
        .IN2(P1_add_368_n120) );
  AND2X1 P1_add_368_U124 ( .IN1(P1_add_368_n117), .IN2(P1_add_368_n120), 
        .Q(P1_add_368_n119) );
  NOR2X0 P1_add_368_U123 ( .QN(P1_N2249), .IN1(P1_add_368_n118), 
        .IN2(P1_add_368_n119) );
  NAND2X0 P1_add_368_U122 ( .IN1(n7089), .IN2(P1_add_368_n117), 
        .QN(P1_add_368_n114) );
  OR2X1 P1_add_368_U121 ( .IN2(n7089), .IN1(P1_add_368_n117), 
        .Q(P1_add_368_n116) );
  NAND2X0 P1_add_368_U120 ( .IN1(P1_N2007), .IN2(P1_add_368_n116), 
        .QN(P1_add_368_n115) );
  NAND2X0 P1_add_368_U119 ( .IN1(P1_add_368_n114), .IN2(P1_add_368_n115), 
        .QN(P1_add_368_n107) );
  OR2X1 P1_add_368_U117 ( .IN2(P1_N2008), .IN1(n7144), .Q(P1_add_368_n111) );
  NAND2X0 P1_add_368_U116 ( .IN1(P1_N2008), .IN2(n7144), .QN(P1_add_368_n112)
         );
  NAND2X0 P1_add_368_U115 ( .IN1(P1_add_368_n111), .IN2(P1_add_368_n112), 
        .QN(P1_add_368_n110) );
  NOR2X0 P1_add_368_U114 ( .QN(P1_add_368_n108), .IN1(P1_add_368_n107), 
        .IN2(P1_add_368_n110) );
  AND2X1 P1_add_368_U113 ( .IN1(P1_add_368_n107), .IN2(P1_add_368_n110), 
        .Q(P1_add_368_n109) );
  NOR2X0 P1_add_368_U112 ( .QN(P1_N2250), .IN1(P1_add_368_n108), 
        .IN2(P1_add_368_n109) );
  NAND2X0 P1_add_368_U111 ( .IN1(n7141), .IN2(P1_add_368_n107), 
        .QN(P1_add_368_n104) );
  OR2X1 P1_add_368_U110 ( .IN2(n7141), .IN1(P1_add_368_n107), 
        .Q(P1_add_368_n106) );
  NAND2X0 P1_add_368_U109 ( .IN1(P1_N2008), .IN2(P1_add_368_n106), 
        .QN(P1_add_368_n105) );
  NAND2X0 P1_add_368_U108 ( .IN1(P1_add_368_n104), .IN2(P1_add_368_n105), 
        .QN(P1_add_368_n97) );
  OR2X1 P1_add_368_U106 ( .IN2(P1_N2009), .IN1(n7136), .Q(P1_add_368_n101) );
  NAND2X0 P1_add_368_U105 ( .IN1(P1_N2009), .IN2(n7136), .QN(P1_add_368_n102)
         );
  NAND2X0 P1_add_368_U104 ( .IN1(P1_add_368_n101), .IN2(P1_add_368_n102), 
        .QN(P1_add_368_n100) );
  NOR2X0 P1_add_368_U103 ( .QN(P1_add_368_n98), .IN1(P1_add_368_n97), 
        .IN2(P1_add_368_n100) );
  AND2X1 P1_add_368_U102 ( .IN1(P1_add_368_n97), .IN2(P1_add_368_n100), 
        .Q(P1_add_368_n99) );
  NOR2X0 P1_add_368_U101 ( .QN(P1_N2251), .IN1(P1_add_368_n98), 
        .IN2(P1_add_368_n99) );
  NAND2X0 P1_add_368_U100 ( .IN1(n7138), .IN2(P1_add_368_n97), 
        .QN(P1_add_368_n94) );
  OR2X1 P1_add_368_U99 ( .IN2(n7138), .IN1(P1_add_368_n97), .Q(P1_add_368_n96)
         );
  NAND2X0 P1_add_368_U98 ( .IN1(P1_N2009), .IN2(P1_add_368_n96), 
        .QN(P1_add_368_n95) );
  NAND2X0 P1_add_368_U97 ( .IN1(P1_add_368_n94), .IN2(P1_add_368_n95), 
        .QN(P1_add_368_n87) );
  OR2X1 P1_add_368_U95 ( .IN2(P1_N2010), .IN1(n7130), .Q(P1_add_368_n91) );
  NAND2X0 P1_add_368_U94 ( .IN1(P1_N2010), .IN2(n7130), .QN(P1_add_368_n92) );
  NAND2X0 P1_add_368_U93 ( .IN1(P1_add_368_n91), .IN2(P1_add_368_n92), 
        .QN(P1_add_368_n90) );
  NOR2X0 P1_add_368_U92 ( .QN(P1_add_368_n88), .IN1(P1_add_368_n87), 
        .IN2(P1_add_368_n90) );
  AND2X1 P1_add_368_U91 ( .IN1(P1_add_368_n87), .IN2(P1_add_368_n90), 
        .Q(P1_add_368_n89) );
  NOR2X0 P1_add_368_U90 ( .QN(P1_N2252), .IN1(P1_add_368_n88), 
        .IN2(P1_add_368_n89) );
  NAND2X0 P1_add_368_U275 ( .IN1(n7072), .IN2(P1_add_368_n10), 
        .QN(P1_add_368_n254) );
  OR2X1 P1_add_368_U274 ( .IN2(n7072), .IN1(P1_add_368_n10), 
        .Q(P1_add_368_n256) );
  NAND2X0 P1_add_368_U273 ( .IN1(P1_N1993), .IN2(P1_add_368_n256), 
        .QN(P1_add_368_n255) );
  NAND2X0 P1_add_368_U272 ( .IN1(P1_add_368_n254), .IN2(P1_add_368_n255), 
        .QN(P1_add_368_n3) );
  NAND2X0 P1_add_368_U271 ( .IN1(n7070), .IN2(P1_add_368_n3), 
        .QN(P1_add_368_n251) );
  OR2X1 P1_add_368_U270 ( .IN2(n7070), .IN1(P1_add_368_n3), 
        .Q(P1_add_368_n253) );
  NAND2X0 P1_add_368_U269 ( .IN1(P1_N1994), .IN2(P1_add_368_n253), 
        .QN(P1_add_368_n252) );
  NAND2X0 P1_add_368_U268 ( .IN1(P1_add_368_n251), .IN2(P1_add_368_n252), 
        .QN(P1_add_368_n244) );
  OR2X1 P1_add_368_U266 ( .IN2(P1_N1995), .IN1(n7067), .Q(P1_add_368_n248) );
  NAND2X0 P1_add_368_U265 ( .IN1(P1_N1995), .IN2(n7067), .QN(P1_add_368_n249)
         );
  NAND2X0 P1_add_368_U264 ( .IN1(P1_add_368_n248), .IN2(P1_add_368_n249), 
        .QN(P1_add_368_n247) );
  NOR2X0 P1_add_368_U263 ( .QN(P1_add_368_n245), .IN1(P1_add_368_n244), 
        .IN2(P1_add_368_n247) );
  AND2X1 P1_add_368_U262 ( .IN1(P1_add_368_n244), .IN2(P1_add_368_n247), 
        .Q(P1_add_368_n246) );
  NOR2X0 P1_add_368_U261 ( .QN(P1_N2237), .IN1(P1_add_368_n245), 
        .IN2(P1_add_368_n246) );
  NAND2X0 P1_add_368_U260 ( .IN1(n7066), .IN2(P1_add_368_n244), 
        .QN(P1_add_368_n241) );
  OR2X1 P1_add_368_U259 ( .IN2(n7066), .IN1(P1_add_368_n244), 
        .Q(P1_add_368_n243) );
  NAND2X0 P1_add_368_U258 ( .IN1(P1_N1995), .IN2(P1_add_368_n243), 
        .QN(P1_add_368_n242) );
  NAND2X0 P1_add_368_U257 ( .IN1(P1_add_368_n241), .IN2(P1_add_368_n242), 
        .QN(P1_add_368_n234) );
  OR2X1 P1_add_368_U255 ( .IN2(P1_N1996), .IN1(n7063), .Q(P1_add_368_n238) );
  NAND2X0 P1_add_368_U254 ( .IN1(P1_N1996), .IN2(n7063), .QN(P1_add_368_n239)
         );
  NAND2X0 P1_add_368_U253 ( .IN1(P1_add_368_n238), .IN2(P1_add_368_n239), 
        .QN(P1_add_368_n237) );
  NOR2X0 P1_add_368_U252 ( .QN(P1_add_368_n235), .IN1(P1_add_368_n234), 
        .IN2(P1_add_368_n237) );
  AND2X1 P1_add_368_U251 ( .IN1(P1_add_368_n234), .IN2(P1_add_368_n237), 
        .Q(P1_add_368_n236) );
  NOR2X0 P1_add_368_U250 ( .QN(P1_N2238), .IN1(P1_add_368_n235), 
        .IN2(P1_add_368_n236) );
  NAND2X0 P1_add_368_U249 ( .IN1(n7062), .IN2(P1_add_368_n234), 
        .QN(P1_add_368_n231) );
  OR2X1 P1_add_368_U248 ( .IN2(n7062), .IN1(P1_add_368_n234), 
        .Q(P1_add_368_n233) );
  NAND2X0 P1_add_368_U247 ( .IN1(P1_N1996), .IN2(P1_add_368_n233), 
        .QN(P1_add_368_n232) );
  NAND2X0 P1_add_368_U246 ( .IN1(P1_add_368_n231), .IN2(P1_add_368_n232), 
        .QN(P1_add_368_n224) );
  OR2X1 P1_add_368_U244 ( .IN2(P1_N1997), .IN1(n7058), .Q(P1_add_368_n228) );
  NAND2X0 P1_add_368_U243 ( .IN1(P1_N1997), .IN2(n7058), .QN(P1_add_368_n229)
         );
  NAND2X0 P1_add_368_U242 ( .IN1(P1_add_368_n228), .IN2(P1_add_368_n229), 
        .QN(P1_add_368_n227) );
  NOR2X0 P1_add_368_U241 ( .QN(P1_add_368_n225), .IN1(P1_add_368_n224), 
        .IN2(P1_add_368_n227) );
  AND2X1 P1_add_368_U240 ( .IN1(P1_add_368_n224), .IN2(P1_add_368_n227), 
        .Q(P1_add_368_n226) );
  NOR2X0 P1_add_368_U239 ( .QN(P1_N2239), .IN1(P1_add_368_n225), 
        .IN2(P1_add_368_n226) );
  NAND2X0 P1_add_368_U238 ( .IN1(n7059), .IN2(P1_add_368_n224), 
        .QN(P1_add_368_n221) );
  OR2X1 P1_add_368_U237 ( .IN2(n7059), .IN1(P1_add_368_n224), 
        .Q(P1_add_368_n223) );
  NAND2X0 P1_add_368_U236 ( .IN1(P1_N1997), .IN2(P1_add_368_n223), 
        .QN(P1_add_368_n222) );
  NAND2X0 P1_add_368_U235 ( .IN1(P1_add_368_n221), .IN2(P1_add_368_n222), 
        .QN(P1_add_368_n214) );
  OR2X1 P1_add_368_U233 ( .IN2(P1_N1998), .IN1(n7056), .Q(P1_add_368_n218) );
  NAND2X0 P1_add_368_U232 ( .IN1(P1_N1998), .IN2(n7056), .QN(P1_add_368_n219)
         );
  NAND2X0 P1_add_368_U231 ( .IN1(P1_add_368_n218), .IN2(P1_add_368_n219), 
        .QN(P1_add_368_n217) );
  NOR2X0 P1_add_368_U230 ( .QN(P1_add_368_n215), .IN1(P1_add_368_n214), 
        .IN2(P1_add_368_n217) );
  AND2X1 P1_add_368_U229 ( .IN1(P1_add_368_n214), .IN2(P1_add_368_n217), 
        .Q(P1_add_368_n216) );
  NOR2X0 P1_add_368_U228 ( .QN(P1_N2240), .IN1(P1_add_368_n215), 
        .IN2(P1_add_368_n216) );
  NAND2X0 P1_add_368_U227 ( .IN1(n7055), .IN2(P1_add_368_n214), 
        .QN(P1_add_368_n211) );
  OR2X1 P1_add_368_U226 ( .IN2(n7055), .IN1(P1_add_368_n214), 
        .Q(P1_add_368_n213) );
  NAND2X0 P1_add_368_U225 ( .IN1(P1_N1998), .IN2(P1_add_368_n213), 
        .QN(P1_add_368_n212) );
  NAND2X0 P1_add_368_U224 ( .IN1(P1_add_368_n211), .IN2(P1_add_368_n212), 
        .QN(P1_add_368_n204) );
  OR2X1 P1_add_368_U222 ( .IN2(P1_N1999), .IN1(n7115), .Q(P1_add_368_n208) );
  NAND2X0 P1_add_368_U221 ( .IN1(P1_N1999), .IN2(n7115), .QN(P1_add_368_n209)
         );
  NAND2X0 P1_add_368_U220 ( .IN1(P1_add_368_n208), .IN2(P1_add_368_n209), 
        .QN(P1_add_368_n207) );
  NOR2X0 P1_add_368_U219 ( .QN(P1_add_368_n205), .IN1(P1_add_368_n204), 
        .IN2(P1_add_368_n207) );
  AND2X1 P1_add_368_U218 ( .IN1(P1_add_368_n204), .IN2(P1_add_368_n207), 
        .Q(P1_add_368_n206) );
  NOR2X0 P1_add_368_U217 ( .QN(P1_N2241), .IN1(P1_add_368_n205), 
        .IN2(P1_add_368_n206) );
  NAND2X0 P1_add_368_U216 ( .IN1(P1_N5163), .IN2(P1_add_368_n204), 
        .QN(P1_add_368_n201) );
  OR2X1 P1_add_368_U215 ( .IN2(P1_N5163), .IN1(P1_add_368_n204), 
        .Q(P1_add_368_n203) );
  NAND2X0 P1_add_368_U214 ( .IN1(P1_N1999), .IN2(P1_add_368_n203), 
        .QN(P1_add_368_n202) );
  NAND2X0 P1_add_368_U213 ( .IN1(P1_add_368_n201), .IN2(P1_add_368_n202), 
        .QN(P1_add_368_n194) );
  OR2X1 P1_add_368_U211 ( .IN2(P1_N2000), .IN1(n7112), .Q(P1_add_368_n198) );
  NAND2X0 P1_add_368_U210 ( .IN1(P1_N2000), .IN2(n7112), .QN(P1_add_368_n199)
         );
  NAND2X0 P1_add_368_U209 ( .IN1(P1_add_368_n198), .IN2(P1_add_368_n199), 
        .QN(P1_add_368_n197) );
  NOR2X0 P1_add_368_U208 ( .QN(P1_add_368_n195), .IN1(P1_add_368_n194), 
        .IN2(P1_add_368_n197) );
  AND2X1 P1_add_368_U207 ( .IN1(P1_add_368_n194), .IN2(P1_add_368_n197), 
        .Q(P1_add_368_n196) );
  NOR2X0 P1_add_368_U206 ( .QN(P1_N2242), .IN1(P1_add_368_n195), 
        .IN2(P1_add_368_n196) );
  NAND2X0 P1_add_368_U205 ( .IN1(n7113), .IN2(P1_add_368_n194), 
        .QN(P1_add_368_n191) );
  OR2X1 P1_add_368_U204 ( .IN2(n7113), .IN1(P1_add_368_n194), 
        .Q(P1_add_368_n193) );
  NAND2X0 P1_add_368_U203 ( .IN1(P1_N2000), .IN2(P1_add_368_n193), 
        .QN(P1_add_368_n192) );
  NAND2X0 P1_add_368_U202 ( .IN1(P1_add_368_n191), .IN2(P1_add_368_n192), 
        .QN(P1_add_368_n184) );
  OR2X1 P1_add_368_U200 ( .IN2(P1_N2001), .IN1(n7109), .Q(P1_add_368_n188) );
  NAND2X0 P1_add_368_U199 ( .IN1(P1_N2001), .IN2(n7109), .QN(P1_add_368_n189)
         );
  NAND2X0 P1_add_368_U198 ( .IN1(P1_add_368_n188), .IN2(P1_add_368_n189), 
        .QN(P1_add_368_n187) );
  NOR2X0 P1_add_368_U197 ( .QN(P1_add_368_n185), .IN1(P1_add_368_n184), 
        .IN2(P1_add_368_n187) );
  AND2X1 P1_add_368_U196 ( .IN1(P1_add_368_n184), .IN2(P1_add_368_n187), 
        .Q(P1_add_368_n186) );
  NOR2X0 P1_add_368_U195 ( .QN(P1_N2243), .IN1(P1_add_368_n185), 
        .IN2(P1_add_368_n186) );
  NAND2X0 P1_add_368_U194 ( .IN1(P1_N5165), .IN2(P1_add_368_n184), 
        .QN(P1_add_368_n181) );
  OR2X1 P1_add_368_U193 ( .IN2(P1_N5165), .IN1(P1_add_368_n184), 
        .Q(P1_add_368_n183) );
  NAND2X0 P1_add_368_U192 ( .IN1(P1_N2001), .IN2(P1_add_368_n183), 
        .QN(P1_add_368_n182) );
  NAND2X0 P1_add_368_U191 ( .IN1(P1_add_368_n181), .IN2(P1_add_368_n182), 
        .QN(P1_add_368_n174) );
  OR2X1 P1_add_368_U189 ( .IN2(P1_N2002), .IN1(n7105), .Q(P1_add_368_n178) );
  NAND2X0 P1_add_368_U188 ( .IN1(P1_N2002), .IN2(n7105), .QN(P1_add_368_n179)
         );
  NAND2X0 P1_add_368_U187 ( .IN1(P1_add_368_n178), .IN2(P1_add_368_n179), 
        .QN(P1_add_368_n177) );
  NOR2X0 P1_add_368_U186 ( .QN(P1_add_368_n175), .IN1(P1_add_368_n174), 
        .IN2(P1_add_368_n177) );
  AND2X1 P1_add_368_U185 ( .IN1(P1_add_368_n174), .IN2(P1_add_368_n177), 
        .Q(P1_add_368_n176) );
  NOR2X0 P1_add_368_U184 ( .QN(P1_N2244), .IN1(P1_add_368_n175), 
        .IN2(P1_add_368_n176) );
  NAND2X0 P1_add_368_U183 ( .IN1(n7106), .IN2(P1_add_368_n174), 
        .QN(P1_add_368_n171) );
  OR2X1 P1_add_368_U308 ( .IN2(P1_N1985), .IN1(n4803), .Q(P1_add_368_n278) );
  NAND2X0 P1_add_368_U307 ( .IN1(P1_N1985), .IN2(n4803), .QN(P1_add_368_n279)
         );
  NAND2X0 P1_add_368_U306 ( .IN1(P1_add_368_n278), .IN2(P1_add_368_n279), 
        .QN(P1_N2227) );
  NAND2X0 P1_add_368_U304 ( .IN1(P1_N1985), .IN2(n7034), .QN(P1_add_368_n151)
         );
  OR2X1 P1_add_368_U303 ( .IN2(P1_add_368_n151), .IN1(n7048), 
        .Q(P1_add_368_n275) );
  NAND2X0 P1_add_368_U302 ( .IN1(n7048), .IN2(P1_add_368_n151), 
        .QN(P1_add_368_n277) );
  NAND2X0 P1_add_368_U301 ( .IN1(P1_N1986), .IN2(P1_add_368_n277), 
        .QN(P1_add_368_n276) );
  NAND2X0 P1_add_368_U300 ( .IN1(P1_add_368_n275), .IN2(P1_add_368_n276), 
        .QN(P1_add_368_n52) );
  NAND2X0 P1_add_368_U299 ( .IN1(n7046), .IN2(P1_add_368_n52), 
        .QN(P1_add_368_n272) );
  OR2X1 P1_add_368_U298 ( .IN2(n7046), .IN1(P1_add_368_n52), 
        .Q(P1_add_368_n274) );
  NAND2X0 P1_add_368_U297 ( .IN1(P1_N1987), .IN2(P1_add_368_n274), 
        .QN(P1_add_368_n273) );
  NAND2X0 P1_add_368_U296 ( .IN1(P1_add_368_n272), .IN2(P1_add_368_n273), 
        .QN(P1_add_368_n45) );
  NAND2X0 P1_add_368_U295 ( .IN1(n7041), .IN2(P1_add_368_n45), 
        .QN(P1_add_368_n269) );
  OR2X1 P1_add_368_U294 ( .IN2(n7041), .IN1(P1_add_368_n45), 
        .Q(P1_add_368_n271) );
  NAND2X0 P1_add_368_U293 ( .IN1(P1_N1988), .IN2(P1_add_368_n271), 
        .QN(P1_add_368_n270) );
  NAND2X0 P1_add_368_U292 ( .IN1(P1_add_368_n269), .IN2(P1_add_368_n270), 
        .QN(P1_add_368_n38) );
  NAND2X0 P1_add_368_U291 ( .IN1(n7036), .IN2(P1_add_368_n38), 
        .QN(P1_add_368_n266) );
  OR2X1 P1_add_368_U290 ( .IN2(n7036), .IN1(P1_add_368_n38), 
        .Q(P1_add_368_n268) );
  NAND2X0 P1_add_368_U289 ( .IN1(P1_N1989), .IN2(P1_add_368_n268), 
        .QN(P1_add_368_n267) );
  NAND2X0 P1_add_368_U288 ( .IN1(P1_add_368_n266), .IN2(P1_add_368_n267), 
        .QN(P1_add_368_n31) );
  NAND2X0 P1_add_368_U287 ( .IN1(n7081), .IN2(P1_add_368_n31), 
        .QN(P1_add_368_n263) );
  OR2X1 P1_add_368_U286 ( .IN2(n7081), .IN1(P1_add_368_n31), 
        .Q(P1_add_368_n265) );
  NAND2X0 P1_add_368_U285 ( .IN1(P1_N1990), .IN2(P1_add_368_n265), 
        .QN(P1_add_368_n264) );
  NAND2X0 P1_add_368_U284 ( .IN1(P1_add_368_n263), .IN2(P1_add_368_n264), 
        .QN(P1_add_368_n24) );
  NAND2X0 P1_add_368_U283 ( .IN1(n7080), .IN2(P1_add_368_n24), 
        .QN(P1_add_368_n260) );
  OR2X1 P1_add_368_U282 ( .IN2(n7080), .IN1(P1_add_368_n24), 
        .Q(P1_add_368_n262) );
  NAND2X0 P1_add_368_U281 ( .IN1(P1_N1991), .IN2(P1_add_368_n262), 
        .QN(P1_add_368_n261) );
  NAND2X0 P1_add_368_U280 ( .IN1(P1_add_368_n260), .IN2(P1_add_368_n261), 
        .QN(P1_add_368_n17) );
  NAND2X0 P1_add_368_U279 ( .IN1(n7075), .IN2(P1_add_368_n17), 
        .QN(P1_add_368_n257) );
  OR2X1 P1_add_368_U278 ( .IN2(n7075), .IN1(P1_add_368_n17), 
        .Q(P1_add_368_n259) );
  NAND2X0 P1_add_368_U277 ( .IN1(P1_N1992), .IN2(P1_add_368_n259), 
        .QN(P1_add_368_n258) );
  NAND2X0 P1_add_368_U276 ( .IN1(P1_add_368_n257), .IN2(P1_add_368_n258), 
        .QN(P1_add_368_n10) );
  NAND2X0 P1_sub_388_U27 ( .IN1(P1_sub_388_n31), .IN2(P1_sub_388_n32), 
        .QN(P1_sub_388_n29) );
  OR2X1 P1_sub_388_U26 ( .IN2(P1_sub_388_n32), .IN1(P1_sub_388_n31), 
        .Q(P1_sub_388_n30) );
  NAND2X0 P1_sub_388_U25 ( .IN1(P1_sub_388_n29), .IN2(P1_sub_388_n30), 
        .QN(P1_N2605) );
  NAND2X0 P1_sub_388_U24 ( .IN1(n7080), .IN2(P1_sub_388_n28), 
        .QN(P1_sub_388_n26) );
  OR2X1 P1_sub_388_U23 ( .IN2(n7080), .IN1(P1_sub_388_n28), .Q(P1_sub_388_n27)
         );
  NAND2X0 P1_sub_388_U22 ( .IN1(P1_sub_388_n26), .IN2(P1_sub_388_n27), 
        .QN(P1_sub_388_n24) );
  NAND2X0 P1_sub_388_U21 ( .IN1(P1_sub_388_n24), .IN2(P1_sub_388_n25), 
        .QN(P1_sub_388_n22) );
  OR2X1 P1_sub_388_U20 ( .IN2(P1_sub_388_n25), .IN1(P1_sub_388_n24), 
        .Q(P1_sub_388_n23) );
  NAND2X0 P1_sub_388_U19 ( .IN1(P1_sub_388_n22), .IN2(P1_sub_388_n23), 
        .QN(P1_N2606) );
  NAND2X0 P1_sub_388_U18 ( .IN1(P1_N5156), .IN2(P1_sub_388_n21), 
        .QN(P1_sub_388_n19) );
  OR2X1 P1_sub_388_U17 ( .IN2(P1_N5156), .IN1(P1_sub_388_n21), 
        .Q(P1_sub_388_n20) );
  NAND2X0 P1_sub_388_U16 ( .IN1(P1_sub_388_n19), .IN2(P1_sub_388_n20), 
        .QN(P1_sub_388_n17) );
  NAND2X0 P1_sub_388_U15 ( .IN1(P1_sub_388_n17), .IN2(P1_sub_388_n18), 
        .QN(P1_sub_388_n15) );
  OR2X1 P1_sub_388_U14 ( .IN2(P1_sub_388_n18), .IN1(P1_sub_388_n17), 
        .Q(P1_sub_388_n16) );
  NAND2X0 P1_sub_388_U13 ( .IN1(P1_sub_388_n15), .IN2(P1_sub_388_n16), 
        .QN(P1_N2607) );
  NAND2X0 P1_sub_388_U12 ( .IN1(n7072), .IN2(P1_sub_388_n14), 
        .QN(P1_sub_388_n12) );
  OR2X1 P1_sub_388_U11 ( .IN2(n7072), .IN1(P1_sub_388_n14), .Q(P1_sub_388_n13)
         );
  NAND2X0 P1_sub_388_U10 ( .IN1(P1_sub_388_n12), .IN2(P1_sub_388_n13), 
        .QN(P1_sub_388_n10) );
  NAND2X0 P1_sub_388_U9 ( .IN1(P1_sub_388_n10), .IN2(P1_sub_388_n11), 
        .QN(P1_sub_388_n8) );
  OR2X1 P1_sub_388_U8 ( .IN2(P1_sub_388_n11), .IN1(P1_sub_388_n10), 
        .Q(P1_sub_388_n9) );
  NAND2X0 P1_sub_388_U7 ( .IN1(P1_sub_388_n8), .IN2(P1_sub_388_n9), 
        .QN(P1_N2608) );
  NAND2X0 P1_sub_388_U6 ( .IN1(n7070), .IN2(P1_sub_388_n7), .QN(P1_sub_388_n5)
         );
  OR2X1 P1_sub_388_U5 ( .IN2(n7070), .IN1(P1_sub_388_n7), .Q(P1_sub_388_n6) );
  NAND2X0 P1_sub_388_U4 ( .IN1(P1_sub_388_n5), .IN2(P1_sub_388_n6), 
        .QN(P1_sub_388_n3) );
  NAND2X0 P1_sub_388_U3 ( .IN1(P1_sub_388_n3), .IN2(P1_sub_388_n4), 
        .QN(P1_sub_388_n1) );
  OR2X1 P1_sub_388_U2 ( .IN2(P1_sub_388_n4), .IN1(P1_sub_388_n3), 
        .Q(P1_sub_388_n2) );
  NAND2X0 P1_sub_388_U1 ( .IN1(P1_sub_388_n1), .IN2(P1_sub_388_n2), 
        .QN(P1_N2609) );
  OR2X1 P1_sub_388_U120 ( .IN2(P1_N5170), .IN1(P1_sub_388_n126), 
        .Q(P1_sub_388_n124) );
  NAND2X0 P1_sub_388_U119 ( .IN1(P1_sub_388_n124), .IN2(P1_sub_388_n125), 
        .QN(P1_sub_388_n123) );
  NAND2X0 P1_sub_388_U118 ( .IN1(P1_sub_388_n122), .IN2(P1_sub_388_n123), 
        .QN(P1_sub_388_n116) );
  NAND2X0 P1_sub_388_U117 ( .IN1(P1_sub_388_n121), .IN2(P1_sub_388_n116), 
        .QN(P1_sub_388_n119) );
  OR2X1 P1_sub_388_U116 ( .IN2(P1_sub_388_n116), .IN1(P1_sub_388_n121), 
        .Q(P1_sub_388_n120) );
  NAND2X0 P1_sub_388_U115 ( .IN1(P1_sub_388_n119), .IN2(P1_sub_388_n120), 
        .QN(P1_N2622) );
  INVX0 P1_sub_388_U114 ( .ZN(P1_sub_388_n105), .INP(P1_N2381) );
  NAND2X0 P1_sub_388_U113 ( .IN1(n7141), .IN2(P1_sub_388_n105), 
        .QN(P1_sub_388_n117) );
  OR2X1 P1_sub_388_U112 ( .IN2(n7141), .IN1(P1_sub_388_n105), 
        .Q(P1_sub_388_n118) );
  NAND2X0 P1_sub_388_U111 ( .IN1(P1_sub_388_n117), .IN2(P1_sub_388_n118), 
        .QN(P1_sub_388_n111) );
  NAND2X0 P1_sub_388_U110 ( .IN1(P1_N5171), .IN2(P1_sub_388_n116), 
        .QN(P1_sub_388_n112) );
  OR2X1 P1_sub_388_U109 ( .IN2(P1_N5171), .IN1(P1_sub_388_n116), 
        .Q(P1_sub_388_n114) );
  NAND2X0 P1_sub_388_U108 ( .IN1(P1_sub_388_n114), .IN2(P1_sub_388_n115), 
        .QN(P1_sub_388_n113) );
  NAND2X0 P1_sub_388_U107 ( .IN1(P1_sub_388_n112), .IN2(P1_sub_388_n113), 
        .QN(P1_sub_388_n106) );
  NAND2X0 P1_sub_388_U106 ( .IN1(P1_sub_388_n111), .IN2(P1_sub_388_n106), 
        .QN(P1_sub_388_n109) );
  OR2X1 P1_sub_388_U105 ( .IN2(P1_sub_388_n106), .IN1(P1_sub_388_n111), 
        .Q(P1_sub_388_n110) );
  NAND2X0 P1_sub_388_U104 ( .IN1(P1_sub_388_n109), .IN2(P1_sub_388_n110), 
        .QN(P1_N2623) );
  INVX0 P1_sub_388_U103 ( .ZN(P1_sub_388_n95), .INP(P1_N2382) );
  NAND2X0 P1_sub_388_U102 ( .IN1(P1_N5173), .IN2(P1_sub_388_n95), 
        .QN(P1_sub_388_n107) );
  OR2X1 P1_sub_388_U101 ( .IN2(P1_N5173), .IN1(P1_sub_388_n95), 
        .Q(P1_sub_388_n108) );
  NAND2X0 P1_sub_388_U100 ( .IN1(P1_sub_388_n107), .IN2(P1_sub_388_n108), 
        .QN(P1_sub_388_n101) );
  NAND2X0 P1_sub_388_U99 ( .IN1(n7141), .IN2(P1_sub_388_n106), 
        .QN(P1_sub_388_n102) );
  OR2X1 P1_sub_388_U98 ( .IN2(n7141), .IN1(P1_sub_388_n106), 
        .Q(P1_sub_388_n104) );
  NAND2X0 P1_sub_388_U97 ( .IN1(P1_sub_388_n104), .IN2(P1_sub_388_n105), 
        .QN(P1_sub_388_n103) );
  NAND2X0 P1_sub_388_U96 ( .IN1(P1_sub_388_n102), .IN2(P1_sub_388_n103), 
        .QN(P1_sub_388_n96) );
  NAND2X0 P1_sub_388_U95 ( .IN1(P1_sub_388_n101), .IN2(P1_sub_388_n96), 
        .QN(P1_sub_388_n99) );
  OR2X1 P1_sub_388_U94 ( .IN2(P1_sub_388_n96), .IN1(P1_sub_388_n101), 
        .Q(P1_sub_388_n100) );
  NAND2X0 P1_sub_388_U93 ( .IN1(P1_sub_388_n99), .IN2(P1_sub_388_n100), 
        .QN(P1_N2624) );
  INVX0 P1_sub_388_U92 ( .ZN(P1_sub_388_n85), .INP(P1_N2383) );
  NAND2X0 P1_sub_388_U91 ( .IN1(n7129), .IN2(P1_sub_388_n85), 
        .QN(P1_sub_388_n97) );
  OR2X1 P1_sub_388_U90 ( .IN2(n7129), .IN1(P1_sub_388_n85), .Q(P1_sub_388_n98)
         );
  NAND2X0 P1_sub_388_U89 ( .IN1(P1_sub_388_n97), .IN2(P1_sub_388_n98), 
        .QN(P1_sub_388_n91) );
  NAND2X0 P1_sub_388_U88 ( .IN1(P1_N5173), .IN2(P1_sub_388_n96), 
        .QN(P1_sub_388_n92) );
  OR2X1 P1_sub_388_U87 ( .IN2(P1_N5173), .IN1(P1_sub_388_n96), 
        .Q(P1_sub_388_n94) );
  NAND2X0 P1_sub_388_U86 ( .IN1(P1_sub_388_n94), .IN2(P1_sub_388_n95), 
        .QN(P1_sub_388_n93) );
  NAND2X0 P1_sub_388_U85 ( .IN1(P1_sub_388_n92), .IN2(P1_sub_388_n93), 
        .QN(P1_sub_388_n86) );
  NAND2X0 P1_sub_388_U84 ( .IN1(P1_sub_388_n91), .IN2(P1_sub_388_n86), 
        .QN(P1_sub_388_n89) );
  OR2X1 P1_sub_388_U83 ( .IN2(P1_sub_388_n86), .IN1(P1_sub_388_n91), 
        .Q(P1_sub_388_n90) );
  NAND2X0 P1_sub_388_U82 ( .IN1(P1_sub_388_n89), .IN2(P1_sub_388_n90), 
        .QN(P1_N2625) );
  INVX0 P1_sub_388_U81 ( .ZN(P1_sub_388_n75), .INP(P1_N2384) );
  NAND2X0 P1_sub_388_U80 ( .IN1(P1_N5175), .IN2(P1_sub_388_n75), 
        .QN(P1_sub_388_n87) );
  OR2X1 P1_sub_388_U79 ( .IN2(P1_N5175), .IN1(P1_sub_388_n75), 
        .Q(P1_sub_388_n88) );
  NAND2X0 P1_sub_388_U78 ( .IN1(P1_sub_388_n87), .IN2(P1_sub_388_n88), 
        .QN(P1_sub_388_n81) );
  NAND2X0 P1_sub_388_U77 ( .IN1(n7129), .IN2(P1_sub_388_n86), 
        .QN(P1_sub_388_n82) );
  OR2X1 P1_sub_388_U76 ( .IN2(n7129), .IN1(P1_sub_388_n86), .Q(P1_sub_388_n84)
         );
  NAND2X0 P1_sub_388_U75 ( .IN1(P1_sub_388_n84), .IN2(P1_sub_388_n85), 
        .QN(P1_sub_388_n83) );
  NAND2X0 P1_sub_388_U74 ( .IN1(P1_sub_388_n82), .IN2(P1_sub_388_n83), 
        .QN(P1_sub_388_n76) );
  NAND2X0 P1_sub_388_U73 ( .IN1(P1_sub_388_n81), .IN2(P1_sub_388_n76), 
        .QN(P1_sub_388_n79) );
  OR2X1 P1_sub_388_U72 ( .IN2(P1_sub_388_n76), .IN1(P1_sub_388_n81), 
        .Q(P1_sub_388_n80) );
  NAND2X0 P1_sub_388_U71 ( .IN1(P1_sub_388_n79), .IN2(P1_sub_388_n80), 
        .QN(P1_N2626) );
  INVX0 P1_sub_388_U70 ( .ZN(P1_sub_388_n64), .INP(P1_N2385) );
  NAND2X0 P1_sub_388_U69 ( .IN1(P1_N5176), .IN2(P1_sub_388_n64), 
        .QN(P1_sub_388_n77) );
  OR2X1 P1_sub_388_U68 ( .IN2(P1_N5176), .IN1(P1_sub_388_n64), 
        .Q(P1_sub_388_n78) );
  NAND2X0 P1_sub_388_U67 ( .IN1(P1_sub_388_n77), .IN2(P1_sub_388_n78), 
        .QN(P1_sub_388_n71) );
  NAND2X0 P1_sub_388_U66 ( .IN1(P1_N5175), .IN2(P1_sub_388_n76), 
        .QN(P1_sub_388_n72) );
  OR2X1 P1_sub_388_U65 ( .IN2(P1_N5175), .IN1(P1_sub_388_n76), 
        .Q(P1_sub_388_n74) );
  NAND2X0 P1_sub_388_U64 ( .IN1(P1_sub_388_n74), .IN2(P1_sub_388_n75), 
        .QN(P1_sub_388_n73) );
  NAND2X0 P1_sub_388_U63 ( .IN1(P1_sub_388_n72), .IN2(P1_sub_388_n73), 
        .QN(P1_sub_388_n65) );
  NAND2X0 P1_sub_388_U62 ( .IN1(P1_sub_388_n71), .IN2(P1_sub_388_n65), 
        .QN(P1_sub_388_n69) );
  OR2X1 P1_sub_388_U61 ( .IN2(P1_sub_388_n65), .IN1(P1_sub_388_n71), 
        .Q(P1_sub_388_n70) );
  NAND2X0 P1_sub_388_U60 ( .IN1(P1_sub_388_n69), .IN2(P1_sub_388_n70), 
        .QN(P1_N2627) );
  OR2X1 P1_sub_388_U58 ( .IN2(P1_N2386), .IN1(n7117), .Q(P1_sub_388_n66) );
  NAND2X0 P1_sub_388_U57 ( .IN1(P1_N2386), .IN2(n7117), .QN(P1_sub_388_n67) );
  NAND2X0 P1_sub_388_U56 ( .IN1(P1_sub_388_n66), .IN2(P1_sub_388_n67), 
        .QN(P1_sub_388_n60) );
  NAND2X0 P1_sub_388_U55 ( .IN1(P1_N5176), .IN2(P1_sub_388_n65), 
        .QN(P1_sub_388_n61) );
  OR2X1 P1_sub_388_U54 ( .IN2(P1_N5176), .IN1(P1_sub_388_n65), 
        .Q(P1_sub_388_n63) );
  NAND2X0 P1_sub_388_U53 ( .IN1(P1_sub_388_n63), .IN2(P1_sub_388_n64), 
        .QN(P1_sub_388_n62) );
  NAND2X0 P1_sub_388_U52 ( .IN1(P1_sub_388_n61), .IN2(P1_sub_388_n62), 
        .QN(P1_sub_388_n59) );
  NAND2X0 P1_sub_388_U51 ( .IN1(P1_sub_388_n60), .IN2(P1_sub_388_n59), 
        .QN(P1_sub_388_n57) );
  OR2X1 P1_sub_388_U50 ( .IN2(P1_sub_388_n60), .IN1(P1_sub_388_n59), 
        .Q(P1_sub_388_n58) );
  NAND2X0 P1_sub_388_U49 ( .IN1(P1_sub_388_n57), .IN2(P1_sub_388_n58), 
        .QN(P1_N2628) );
  NAND2X0 P1_sub_388_U48 ( .IN1(n7046), .IN2(P1_sub_388_n56), 
        .QN(P1_sub_388_n54) );
  OR2X1 P1_sub_388_U47 ( .IN2(n7046), .IN1(P1_sub_388_n56), .Q(P1_sub_388_n55)
         );
  NAND2X0 P1_sub_388_U46 ( .IN1(P1_sub_388_n54), .IN2(P1_sub_388_n55), 
        .QN(P1_sub_388_n52) );
  NAND2X0 P1_sub_388_U45 ( .IN1(P1_sub_388_n52), .IN2(P1_sub_388_n53), 
        .QN(P1_sub_388_n50) );
  OR2X1 P1_sub_388_U44 ( .IN2(P1_sub_388_n53), .IN1(P1_sub_388_n52), 
        .Q(P1_sub_388_n51) );
  NAND2X0 P1_sub_388_U43 ( .IN1(P1_sub_388_n50), .IN2(P1_sub_388_n51), 
        .QN(P1_N2602) );
  NAND2X0 P1_sub_388_U42 ( .IN1(P1_N5152), .IN2(P1_sub_388_n49), 
        .QN(P1_sub_388_n47) );
  OR2X1 P1_sub_388_U41 ( .IN2(P1_N5152), .IN1(P1_sub_388_n49), 
        .Q(P1_sub_388_n48) );
  NAND2X0 P1_sub_388_U40 ( .IN1(P1_sub_388_n47), .IN2(P1_sub_388_n48), 
        .QN(P1_sub_388_n45) );
  NAND2X0 P1_sub_388_U39 ( .IN1(P1_sub_388_n45), .IN2(P1_sub_388_n46), 
        .QN(P1_sub_388_n43) );
  OR2X1 P1_sub_388_U38 ( .IN2(P1_sub_388_n46), .IN1(P1_sub_388_n45), 
        .Q(P1_sub_388_n44) );
  NAND2X0 P1_sub_388_U37 ( .IN1(P1_sub_388_n43), .IN2(P1_sub_388_n44), 
        .QN(P1_N2603) );
  NAND2X0 P1_sub_388_U36 ( .IN1(n7036), .IN2(P1_sub_388_n42), 
        .QN(P1_sub_388_n40) );
  OR2X1 P1_sub_388_U35 ( .IN2(n7036), .IN1(P1_sub_388_n42), .Q(P1_sub_388_n41)
         );
  NAND2X0 P1_sub_388_U34 ( .IN1(P1_sub_388_n40), .IN2(P1_sub_388_n41), 
        .QN(P1_sub_388_n38) );
  NAND2X0 P1_sub_388_U33 ( .IN1(P1_sub_388_n38), .IN2(P1_sub_388_n39), 
        .QN(P1_sub_388_n36) );
  OR2X1 P1_sub_388_U32 ( .IN2(P1_sub_388_n39), .IN1(P1_sub_388_n38), 
        .Q(P1_sub_388_n37) );
  NAND2X0 P1_sub_388_U31 ( .IN1(P1_sub_388_n36), .IN2(P1_sub_388_n37), 
        .QN(P1_N2604) );
  NAND2X0 P1_sub_388_U30 ( .IN1(n7081), .IN2(P1_sub_388_n35), 
        .QN(P1_sub_388_n33) );
  OR2X1 P1_sub_388_U29 ( .IN2(n7081), .IN1(P1_sub_388_n35), .Q(P1_sub_388_n34)
         );
  NAND2X0 P1_sub_388_U28 ( .IN1(P1_sub_388_n33), .IN2(P1_sub_388_n34), 
        .QN(P1_sub_388_n31) );
  NAND2X0 P1_sub_388_U213 ( .IN1(P1_sub_388_n212), .IN2(P1_sub_388_n213), 
        .QN(P1_sub_388_n211) );
  NAND2X0 P1_sub_388_U212 ( .IN1(P1_sub_388_n210), .IN2(P1_sub_388_n211), 
        .QN(P1_sub_388_n204) );
  NAND2X0 P1_sub_388_U211 ( .IN1(P1_sub_388_n209), .IN2(P1_sub_388_n204), 
        .QN(P1_sub_388_n207) );
  OR2X1 P1_sub_388_U210 ( .IN2(P1_sub_388_n204), .IN1(P1_sub_388_n209), 
        .Q(P1_sub_388_n208) );
  NAND2X0 P1_sub_388_U209 ( .IN1(P1_sub_388_n207), .IN2(P1_sub_388_n208), 
        .QN(P1_N2614) );
  INVX0 P1_sub_388_U208 ( .ZN(P1_sub_388_n193), .INP(P1_N2373) );
  NAND2X0 P1_sub_388_U207 ( .IN1(P1_N5164), .IN2(P1_sub_388_n193), 
        .QN(P1_sub_388_n205) );
  OR2X1 P1_sub_388_U206 ( .IN2(P1_N5164), .IN1(P1_sub_388_n193), 
        .Q(P1_sub_388_n206) );
  NAND2X0 P1_sub_388_U205 ( .IN1(P1_sub_388_n205), .IN2(P1_sub_388_n206), 
        .QN(P1_sub_388_n199) );
  NAND2X0 P1_sub_388_U204 ( .IN1(n7116), .IN2(P1_sub_388_n204), 
        .QN(P1_sub_388_n200) );
  OR2X1 P1_sub_388_U203 ( .IN2(n7116), .IN1(P1_sub_388_n204), 
        .Q(P1_sub_388_n202) );
  NAND2X0 P1_sub_388_U202 ( .IN1(P1_sub_388_n202), .IN2(P1_sub_388_n203), 
        .QN(P1_sub_388_n201) );
  NAND2X0 P1_sub_388_U201 ( .IN1(P1_sub_388_n200), .IN2(P1_sub_388_n201), 
        .QN(P1_sub_388_n194) );
  NAND2X0 P1_sub_388_U200 ( .IN1(P1_sub_388_n199), .IN2(P1_sub_388_n194), 
        .QN(P1_sub_388_n197) );
  OR2X1 P1_sub_388_U199 ( .IN2(P1_sub_388_n194), .IN1(P1_sub_388_n199), 
        .Q(P1_sub_388_n198) );
  NAND2X0 P1_sub_388_U198 ( .IN1(P1_sub_388_n197), .IN2(P1_sub_388_n198), 
        .QN(P1_N2615) );
  INVX0 P1_sub_388_U197 ( .ZN(P1_sub_388_n183), .INP(P1_N2374) );
  NAND2X0 P1_sub_388_U196 ( .IN1(P1_N5165), .IN2(P1_sub_388_n183), 
        .QN(P1_sub_388_n195) );
  OR2X1 P1_sub_388_U195 ( .IN2(P1_N5165), .IN1(P1_sub_388_n183), 
        .Q(P1_sub_388_n196) );
  NAND2X0 P1_sub_388_U194 ( .IN1(P1_sub_388_n195), .IN2(P1_sub_388_n196), 
        .QN(P1_sub_388_n189) );
  NAND2X0 P1_sub_388_U193 ( .IN1(n7113), .IN2(P1_sub_388_n194), 
        .QN(P1_sub_388_n190) );
  OR2X1 P1_sub_388_U192 ( .IN2(n7113), .IN1(P1_sub_388_n194), 
        .Q(P1_sub_388_n192) );
  NAND2X0 P1_sub_388_U191 ( .IN1(P1_sub_388_n192), .IN2(P1_sub_388_n193), 
        .QN(P1_sub_388_n191) );
  NAND2X0 P1_sub_388_U190 ( .IN1(P1_sub_388_n190), .IN2(P1_sub_388_n191), 
        .QN(P1_sub_388_n184) );
  NAND2X0 P1_sub_388_U189 ( .IN1(P1_sub_388_n189), .IN2(P1_sub_388_n184), 
        .QN(P1_sub_388_n187) );
  OR2X1 P1_sub_388_U188 ( .IN2(P1_sub_388_n184), .IN1(P1_sub_388_n189), 
        .Q(P1_sub_388_n188) );
  NAND2X0 P1_sub_388_U187 ( .IN1(P1_sub_388_n187), .IN2(P1_sub_388_n188), 
        .QN(P1_N2616) );
  INVX0 P1_sub_388_U186 ( .ZN(P1_sub_388_n173), .INP(P1_N2375) );
  NAND2X0 P1_sub_388_U185 ( .IN1(n7106), .IN2(P1_sub_388_n173), 
        .QN(P1_sub_388_n185) );
  OR2X1 P1_sub_388_U184 ( .IN2(n7106), .IN1(P1_sub_388_n173), 
        .Q(P1_sub_388_n186) );
  NAND2X0 P1_sub_388_U183 ( .IN1(P1_sub_388_n185), .IN2(P1_sub_388_n186), 
        .QN(P1_sub_388_n179) );
  NAND2X0 P1_sub_388_U182 ( .IN1(P1_N5165), .IN2(P1_sub_388_n184), 
        .QN(P1_sub_388_n180) );
  OR2X1 P1_sub_388_U181 ( .IN2(P1_N5165), .IN1(P1_sub_388_n184), 
        .Q(P1_sub_388_n182) );
  NAND2X0 P1_sub_388_U180 ( .IN1(P1_sub_388_n182), .IN2(P1_sub_388_n183), 
        .QN(P1_sub_388_n181) );
  NAND2X0 P1_sub_388_U179 ( .IN1(P1_sub_388_n180), .IN2(P1_sub_388_n181), 
        .QN(P1_sub_388_n174) );
  NAND2X0 P1_sub_388_U178 ( .IN1(P1_sub_388_n179), .IN2(P1_sub_388_n174), 
        .QN(P1_sub_388_n177) );
  OR2X1 P1_sub_388_U177 ( .IN2(P1_sub_388_n174), .IN1(P1_sub_388_n179), 
        .Q(P1_sub_388_n178) );
  NAND2X0 P1_sub_388_U176 ( .IN1(P1_sub_388_n177), .IN2(P1_sub_388_n178), 
        .QN(P1_N2617) );
  INVX0 P1_sub_388_U175 ( .ZN(P1_sub_388_n163), .INP(P1_N2376) );
  NAND2X0 P1_sub_388_U174 ( .IN1(n7103), .IN2(P1_sub_388_n163), 
        .QN(P1_sub_388_n175) );
  OR2X1 P1_sub_388_U173 ( .IN2(n7103), .IN1(P1_sub_388_n163), 
        .Q(P1_sub_388_n176) );
  NAND2X0 P1_sub_388_U172 ( .IN1(P1_sub_388_n175), .IN2(P1_sub_388_n176), 
        .QN(P1_sub_388_n169) );
  NAND2X0 P1_sub_388_U171 ( .IN1(n7106), .IN2(P1_sub_388_n174), 
        .QN(P1_sub_388_n170) );
  OR2X1 P1_sub_388_U170 ( .IN2(n7106), .IN1(P1_sub_388_n174), 
        .Q(P1_sub_388_n172) );
  NAND2X0 P1_sub_388_U169 ( .IN1(P1_sub_388_n172), .IN2(P1_sub_388_n173), 
        .QN(P1_sub_388_n171) );
  NAND2X0 P1_sub_388_U168 ( .IN1(P1_sub_388_n170), .IN2(P1_sub_388_n171), 
        .QN(P1_sub_388_n164) );
  NAND2X0 P1_sub_388_U167 ( .IN1(P1_sub_388_n169), .IN2(P1_sub_388_n164), 
        .QN(P1_sub_388_n167) );
  OR2X1 P1_sub_388_U166 ( .IN2(P1_sub_388_n164), .IN1(P1_sub_388_n169), 
        .Q(P1_sub_388_n168) );
  NAND2X0 P1_sub_388_U165 ( .IN1(P1_sub_388_n167), .IN2(P1_sub_388_n168), 
        .QN(P1_N2618) );
  INVX0 P1_sub_388_U164 ( .ZN(P1_sub_388_n145), .INP(P1_N2377) );
  NAND2X0 P1_sub_388_U163 ( .IN1(n7099), .IN2(P1_sub_388_n145), 
        .QN(P1_sub_388_n165) );
  OR2X1 P1_sub_388_U162 ( .IN2(n7099), .IN1(P1_sub_388_n145), 
        .Q(P1_sub_388_n166) );
  NAND2X0 P1_sub_388_U161 ( .IN1(P1_sub_388_n165), .IN2(P1_sub_388_n166), 
        .QN(P1_sub_388_n159) );
  NAND2X0 P1_sub_388_U160 ( .IN1(n7103), .IN2(P1_sub_388_n164), 
        .QN(P1_sub_388_n160) );
  OR2X1 P1_sub_388_U159 ( .IN2(n7103), .IN1(P1_sub_388_n164), 
        .Q(P1_sub_388_n162) );
  NAND2X0 P1_sub_388_U158 ( .IN1(P1_sub_388_n162), .IN2(P1_sub_388_n163), 
        .QN(P1_sub_388_n161) );
  NAND2X0 P1_sub_388_U157 ( .IN1(P1_sub_388_n160), .IN2(P1_sub_388_n161), 
        .QN(P1_sub_388_n146) );
  NAND2X0 P1_sub_388_U156 ( .IN1(P1_sub_388_n159), .IN2(P1_sub_388_n146), 
        .QN(P1_sub_388_n157) );
  OR2X1 P1_sub_388_U155 ( .IN2(P1_sub_388_n146), .IN1(P1_sub_388_n159), 
        .Q(P1_sub_388_n158) );
  NAND2X0 P1_sub_388_U154 ( .IN1(P1_sub_388_n157), .IN2(P1_sub_388_n158), 
        .QN(P1_N2619) );
  NAND2X0 P1_sub_388_U153 ( .IN1(P1_N5150), .IN2(P1_sub_388_n156), 
        .QN(P1_sub_388_n153) );
  NAND2X0 P1_sub_388_U152 ( .IN1(P1_N2359), .IN2(n7048), .QN(P1_sub_388_n154)
         );
  NAND2X0 P1_sub_388_U151 ( .IN1(P1_sub_388_n153), .IN2(P1_sub_388_n154), 
        .QN(P1_sub_388_n151) );
  NAND2X0 P1_sub_388_U150 ( .IN1(P1_sub_388_n151), .IN2(P1_sub_388_n152), 
        .QN(P1_sub_388_n149) );
  OR2X1 P1_sub_388_U149 ( .IN2(P1_sub_388_n152), .IN1(P1_sub_388_n151), 
        .Q(P1_sub_388_n150) );
  NAND2X0 P1_sub_388_U148 ( .IN1(P1_sub_388_n149), .IN2(P1_sub_388_n150), 
        .QN(P1_N2601) );
  INVX0 P1_sub_388_U147 ( .ZN(P1_sub_388_n135), .INP(P1_N2378) );
  NAND2X0 P1_sub_388_U146 ( .IN1(P1_N5169), .IN2(P1_sub_388_n135), 
        .QN(P1_sub_388_n147) );
  OR2X1 P1_sub_388_U145 ( .IN2(P1_N5169), .IN1(P1_sub_388_n135), 
        .Q(P1_sub_388_n148) );
  NAND2X0 P1_sub_388_U144 ( .IN1(P1_sub_388_n147), .IN2(P1_sub_388_n148), 
        .QN(P1_sub_388_n141) );
  NAND2X0 P1_sub_388_U143 ( .IN1(n7099), .IN2(P1_sub_388_n146), 
        .QN(P1_sub_388_n142) );
  OR2X1 P1_sub_388_U142 ( .IN2(n7099), .IN1(P1_sub_388_n146), 
        .Q(P1_sub_388_n144) );
  NAND2X0 P1_sub_388_U141 ( .IN1(P1_sub_388_n144), .IN2(P1_sub_388_n145), 
        .QN(P1_sub_388_n143) );
  NAND2X0 P1_sub_388_U140 ( .IN1(P1_sub_388_n142), .IN2(P1_sub_388_n143), 
        .QN(P1_sub_388_n136) );
  NAND2X0 P1_sub_388_U139 ( .IN1(P1_sub_388_n141), .IN2(P1_sub_388_n136), 
        .QN(P1_sub_388_n139) );
  OR2X1 P1_sub_388_U138 ( .IN2(P1_sub_388_n136), .IN1(P1_sub_388_n141), 
        .Q(P1_sub_388_n140) );
  NAND2X0 P1_sub_388_U137 ( .IN1(P1_sub_388_n139), .IN2(P1_sub_388_n140), 
        .QN(P1_N2620) );
  INVX0 P1_sub_388_U136 ( .ZN(P1_sub_388_n125), .INP(P1_N2379) );
  NAND2X0 P1_sub_388_U135 ( .IN1(P1_N5170), .IN2(P1_sub_388_n125), 
        .QN(P1_sub_388_n137) );
  OR2X1 P1_sub_388_U134 ( .IN2(P1_N5170), .IN1(P1_sub_388_n125), 
        .Q(P1_sub_388_n138) );
  NAND2X0 P1_sub_388_U133 ( .IN1(P1_sub_388_n137), .IN2(P1_sub_388_n138), 
        .QN(P1_sub_388_n131) );
  NAND2X0 P1_sub_388_U132 ( .IN1(P1_N5169), .IN2(P1_sub_388_n136), 
        .QN(P1_sub_388_n132) );
  OR2X1 P1_sub_388_U131 ( .IN2(P1_N5169), .IN1(P1_sub_388_n136), 
        .Q(P1_sub_388_n134) );
  NAND2X0 P1_sub_388_U130 ( .IN1(P1_sub_388_n134), .IN2(P1_sub_388_n135), 
        .QN(P1_sub_388_n133) );
  NAND2X0 P1_sub_388_U129 ( .IN1(P1_sub_388_n132), .IN2(P1_sub_388_n133), 
        .QN(P1_sub_388_n126) );
  NAND2X0 P1_sub_388_U128 ( .IN1(P1_sub_388_n131), .IN2(P1_sub_388_n126), 
        .QN(P1_sub_388_n129) );
  OR2X1 P1_sub_388_U127 ( .IN2(P1_sub_388_n126), .IN1(P1_sub_388_n131), 
        .Q(P1_sub_388_n130) );
  NAND2X0 P1_sub_388_U126 ( .IN1(P1_sub_388_n129), .IN2(P1_sub_388_n130), 
        .QN(P1_N2621) );
  INVX0 P1_sub_388_U125 ( .ZN(P1_sub_388_n115), .INP(P1_N2380) );
  NAND2X0 P1_sub_388_U124 ( .IN1(P1_N5171), .IN2(P1_sub_388_n115), 
        .QN(P1_sub_388_n127) );
  OR2X1 P1_sub_388_U123 ( .IN2(P1_N5171), .IN1(P1_sub_388_n115), 
        .Q(P1_sub_388_n128) );
  NAND2X0 P1_sub_388_U122 ( .IN1(P1_sub_388_n127), .IN2(P1_sub_388_n128), 
        .QN(P1_sub_388_n121) );
  NAND2X0 P1_sub_388_U121 ( .IN1(P1_N5170), .IN2(P1_sub_388_n126), 
        .QN(P1_sub_388_n122) );
  NAND2X0 P1_sub_388_U306 ( .IN1(P1_sub_388_n152), .IN2(P1_sub_388_n280), 
        .QN(P1_N2600) );
  INVX0 P1_sub_388_U305 ( .ZN(P1_sub_388_n243), .INP(P1_N2368) );
  NAND2X0 P1_sub_388_U304 ( .IN1(n7066), .IN2(P1_sub_388_n243), 
        .QN(P1_sub_388_n278) );
  OR2X1 P1_sub_388_U303 ( .IN2(n7066), .IN1(P1_sub_388_n243), 
        .Q(P1_sub_388_n279) );
  NAND2X0 P1_sub_388_U302 ( .IN1(P1_sub_388_n278), .IN2(P1_sub_388_n279), 
        .QN(P1_sub_388_n249) );
  NAND2X0 P1_sub_388_U301 ( .IN1(P1_N5150), .IN2(P1_sub_388_n152), 
        .QN(P1_sub_388_n274) );
  NAND2X0 P1_sub_388_U299 ( .IN1(P1_sub_388_n277), .IN2(n7048), 
        .QN(P1_sub_388_n276) );
  INVX0 P1_sub_388_U298 ( .ZN(P1_sub_388_n156), .INP(P1_N2359) );
  NAND2X0 P1_sub_388_U297 ( .IN1(P1_sub_388_n276), .IN2(P1_sub_388_n156), 
        .QN(P1_sub_388_n275) );
  NAND2X0 P1_sub_388_U296 ( .IN1(P1_sub_388_n274), .IN2(P1_sub_388_n275), 
        .QN(P1_sub_388_n53) );
  NAND2X0 P1_sub_388_U295 ( .IN1(n7046), .IN2(P1_sub_388_n53), 
        .QN(P1_sub_388_n271) );
  OR2X1 P1_sub_388_U294 ( .IN2(n7046), .IN1(P1_sub_388_n53), 
        .Q(P1_sub_388_n273) );
  INVX0 P1_sub_388_U293 ( .ZN(P1_sub_388_n56), .INP(P1_N2360) );
  NAND2X0 P1_sub_388_U292 ( .IN1(P1_sub_388_n273), .IN2(P1_sub_388_n56), 
        .QN(P1_sub_388_n272) );
  NAND2X0 P1_sub_388_U291 ( .IN1(P1_sub_388_n271), .IN2(P1_sub_388_n272), 
        .QN(P1_sub_388_n46) );
  NAND2X0 P1_sub_388_U290 ( .IN1(P1_N5152), .IN2(P1_sub_388_n46), 
        .QN(P1_sub_388_n268) );
  OR2X1 P1_sub_388_U289 ( .IN2(P1_N5152), .IN1(P1_sub_388_n46), 
        .Q(P1_sub_388_n270) );
  INVX0 P1_sub_388_U288 ( .ZN(P1_sub_388_n49), .INP(P1_N2361) );
  NAND2X0 P1_sub_388_U287 ( .IN1(P1_sub_388_n270), .IN2(P1_sub_388_n49), 
        .QN(P1_sub_388_n269) );
  NAND2X0 P1_sub_388_U286 ( .IN1(P1_sub_388_n268), .IN2(P1_sub_388_n269), 
        .QN(P1_sub_388_n39) );
  NAND2X0 P1_sub_388_U285 ( .IN1(n7036), .IN2(P1_sub_388_n39), 
        .QN(P1_sub_388_n265) );
  OR2X1 P1_sub_388_U284 ( .IN2(n7036), .IN1(P1_sub_388_n39), 
        .Q(P1_sub_388_n267) );
  INVX0 P1_sub_388_U283 ( .ZN(P1_sub_388_n42), .INP(P1_N2362) );
  NAND2X0 P1_sub_388_U282 ( .IN1(P1_sub_388_n267), .IN2(P1_sub_388_n42), 
        .QN(P1_sub_388_n266) );
  NAND2X0 P1_sub_388_U281 ( .IN1(P1_sub_388_n265), .IN2(P1_sub_388_n266), 
        .QN(P1_sub_388_n32) );
  NAND2X0 P1_sub_388_U280 ( .IN1(n7081), .IN2(P1_sub_388_n32), 
        .QN(P1_sub_388_n262) );
  OR2X1 P1_sub_388_U279 ( .IN2(n7081), .IN1(P1_sub_388_n32), 
        .Q(P1_sub_388_n264) );
  INVX0 P1_sub_388_U278 ( .ZN(P1_sub_388_n35), .INP(P1_N2363) );
  NAND2X0 P1_sub_388_U277 ( .IN1(P1_sub_388_n264), .IN2(P1_sub_388_n35), 
        .QN(P1_sub_388_n263) );
  NAND2X0 P1_sub_388_U276 ( .IN1(P1_sub_388_n262), .IN2(P1_sub_388_n263), 
        .QN(P1_sub_388_n25) );
  NAND2X0 P1_sub_388_U275 ( .IN1(n7080), .IN2(P1_sub_388_n25), 
        .QN(P1_sub_388_n259) );
  OR2X1 P1_sub_388_U274 ( .IN2(n7080), .IN1(P1_sub_388_n25), 
        .Q(P1_sub_388_n261) );
  INVX0 P1_sub_388_U273 ( .ZN(P1_sub_388_n28), .INP(P1_N2364) );
  NAND2X0 P1_sub_388_U272 ( .IN1(P1_sub_388_n261), .IN2(P1_sub_388_n28), 
        .QN(P1_sub_388_n260) );
  NAND2X0 P1_sub_388_U271 ( .IN1(P1_sub_388_n259), .IN2(P1_sub_388_n260), 
        .QN(P1_sub_388_n18) );
  NAND2X0 P1_sub_388_U270 ( .IN1(P1_N5156), .IN2(P1_sub_388_n18), 
        .QN(P1_sub_388_n256) );
  OR2X1 P1_sub_388_U269 ( .IN2(P1_N5156), .IN1(P1_sub_388_n18), 
        .Q(P1_sub_388_n258) );
  INVX0 P1_sub_388_U268 ( .ZN(P1_sub_388_n21), .INP(P1_N2365) );
  NAND2X0 P1_sub_388_U267 ( .IN1(P1_sub_388_n258), .IN2(P1_sub_388_n21), 
        .QN(P1_sub_388_n257) );
  NAND2X0 P1_sub_388_U266 ( .IN1(P1_sub_388_n256), .IN2(P1_sub_388_n257), 
        .QN(P1_sub_388_n11) );
  NAND2X0 P1_sub_388_U265 ( .IN1(n7072), .IN2(P1_sub_388_n11), 
        .QN(P1_sub_388_n253) );
  OR2X1 P1_sub_388_U264 ( .IN2(n7072), .IN1(P1_sub_388_n11), 
        .Q(P1_sub_388_n255) );
  INVX0 P1_sub_388_U263 ( .ZN(P1_sub_388_n14), .INP(P1_N2366) );
  NAND2X0 P1_sub_388_U262 ( .IN1(P1_sub_388_n255), .IN2(P1_sub_388_n14), 
        .QN(P1_sub_388_n254) );
  NAND2X0 P1_sub_388_U261 ( .IN1(P1_sub_388_n253), .IN2(P1_sub_388_n254), 
        .QN(P1_sub_388_n4) );
  NAND2X0 P1_sub_388_U260 ( .IN1(n7070), .IN2(P1_sub_388_n4), 
        .QN(P1_sub_388_n250) );
  OR2X1 P1_sub_388_U259 ( .IN2(n7070), .IN1(P1_sub_388_n4), 
        .Q(P1_sub_388_n252) );
  INVX0 P1_sub_388_U258 ( .ZN(P1_sub_388_n7), .INP(P1_N2367) );
  NAND2X0 P1_sub_388_U257 ( .IN1(P1_sub_388_n252), .IN2(P1_sub_388_n7), 
        .QN(P1_sub_388_n251) );
  NAND2X0 P1_sub_388_U256 ( .IN1(P1_sub_388_n250), .IN2(P1_sub_388_n251), 
        .QN(P1_sub_388_n244) );
  NAND2X0 P1_sub_388_U255 ( .IN1(P1_sub_388_n249), .IN2(P1_sub_388_n244), 
        .QN(P1_sub_388_n247) );
  OR2X1 P1_sub_388_U254 ( .IN2(P1_sub_388_n244), .IN1(P1_sub_388_n249), 
        .Q(P1_sub_388_n248) );
  NAND2X0 P1_sub_388_U253 ( .IN1(P1_sub_388_n247), .IN2(P1_sub_388_n248), 
        .QN(P1_N2610) );
  INVX0 P1_sub_388_U252 ( .ZN(P1_sub_388_n233), .INP(P1_N2369) );
  NAND2X0 P1_sub_388_U251 ( .IN1(n7062), .IN2(P1_sub_388_n233), 
        .QN(P1_sub_388_n245) );
  OR2X1 P1_sub_388_U250 ( .IN2(n7062), .IN1(P1_sub_388_n233), 
        .Q(P1_sub_388_n246) );
  NAND2X0 P1_sub_388_U249 ( .IN1(P1_sub_388_n245), .IN2(P1_sub_388_n246), 
        .QN(P1_sub_388_n239) );
  NAND2X0 P1_sub_388_U248 ( .IN1(n7066), .IN2(P1_sub_388_n244), 
        .QN(P1_sub_388_n240) );
  OR2X1 P1_sub_388_U247 ( .IN2(n7066), .IN1(P1_sub_388_n244), 
        .Q(P1_sub_388_n242) );
  NAND2X0 P1_sub_388_U246 ( .IN1(P1_sub_388_n242), .IN2(P1_sub_388_n243), 
        .QN(P1_sub_388_n241) );
  NAND2X0 P1_sub_388_U245 ( .IN1(P1_sub_388_n240), .IN2(P1_sub_388_n241), 
        .QN(P1_sub_388_n234) );
  NAND2X0 P1_sub_388_U244 ( .IN1(P1_sub_388_n239), .IN2(P1_sub_388_n234), 
        .QN(P1_sub_388_n237) );
  OR2X1 P1_sub_388_U243 ( .IN2(P1_sub_388_n234), .IN1(P1_sub_388_n239), 
        .Q(P1_sub_388_n238) );
  NAND2X0 P1_sub_388_U242 ( .IN1(P1_sub_388_n237), .IN2(P1_sub_388_n238), 
        .QN(P1_N2611) );
  INVX0 P1_sub_388_U241 ( .ZN(P1_sub_388_n223), .INP(P1_N2370) );
  NAND2X0 P1_sub_388_U240 ( .IN1(n7059), .IN2(P1_sub_388_n223), 
        .QN(P1_sub_388_n235) );
  OR2X1 P1_sub_388_U239 ( .IN2(n7059), .IN1(P1_sub_388_n223), 
        .Q(P1_sub_388_n236) );
  NAND2X0 P1_sub_388_U238 ( .IN1(P1_sub_388_n235), .IN2(P1_sub_388_n236), 
        .QN(P1_sub_388_n229) );
  NAND2X0 P1_sub_388_U237 ( .IN1(n7062), .IN2(P1_sub_388_n234), 
        .QN(P1_sub_388_n230) );
  OR2X1 P1_sub_388_U236 ( .IN2(n7062), .IN1(P1_sub_388_n234), 
        .Q(P1_sub_388_n232) );
  NAND2X0 P1_sub_388_U235 ( .IN1(P1_sub_388_n232), .IN2(P1_sub_388_n233), 
        .QN(P1_sub_388_n231) );
  NAND2X0 P1_sub_388_U234 ( .IN1(P1_sub_388_n230), .IN2(P1_sub_388_n231), 
        .QN(P1_sub_388_n224) );
  NAND2X0 P1_sub_388_U233 ( .IN1(P1_sub_388_n229), .IN2(P1_sub_388_n224), 
        .QN(P1_sub_388_n227) );
  OR2X1 P1_sub_388_U232 ( .IN2(P1_sub_388_n224), .IN1(P1_sub_388_n229), 
        .Q(P1_sub_388_n228) );
  NAND2X0 P1_sub_388_U231 ( .IN1(P1_sub_388_n227), .IN2(P1_sub_388_n228), 
        .QN(P1_N2612) );
  INVX0 P1_sub_388_U230 ( .ZN(P1_sub_388_n213), .INP(P1_N2371) );
  NAND2X0 P1_sub_388_U229 ( .IN1(P1_N5162), .IN2(P1_sub_388_n213), 
        .QN(P1_sub_388_n225) );
  OR2X1 P1_sub_388_U228 ( .IN2(P1_N5162), .IN1(P1_sub_388_n213), 
        .Q(P1_sub_388_n226) );
  NAND2X0 P1_sub_388_U227 ( .IN1(P1_sub_388_n225), .IN2(P1_sub_388_n226), 
        .QN(P1_sub_388_n219) );
  NAND2X0 P1_sub_388_U226 ( .IN1(n7059), .IN2(P1_sub_388_n224), 
        .QN(P1_sub_388_n220) );
  OR2X1 P1_sub_388_U225 ( .IN2(n7059), .IN1(P1_sub_388_n224), 
        .Q(P1_sub_388_n222) );
  NAND2X0 P1_sub_388_U224 ( .IN1(P1_sub_388_n222), .IN2(P1_sub_388_n223), 
        .QN(P1_sub_388_n221) );
  NAND2X0 P1_sub_388_U223 ( .IN1(P1_sub_388_n220), .IN2(P1_sub_388_n221), 
        .QN(P1_sub_388_n214) );
  NAND2X0 P1_sub_388_U222 ( .IN1(P1_sub_388_n219), .IN2(P1_sub_388_n214), 
        .QN(P1_sub_388_n217) );
  OR2X1 P1_sub_388_U221 ( .IN2(P1_sub_388_n214), .IN1(P1_sub_388_n219), 
        .Q(P1_sub_388_n218) );
  NAND2X0 P1_sub_388_U220 ( .IN1(P1_sub_388_n217), .IN2(P1_sub_388_n218), 
        .QN(P1_N2613) );
  INVX0 P1_sub_388_U219 ( .ZN(P1_sub_388_n203), .INP(P1_N2372) );
  NAND2X0 P1_sub_388_U218 ( .IN1(n7116), .IN2(P1_sub_388_n203), 
        .QN(P1_sub_388_n215) );
  OR2X1 P1_sub_388_U217 ( .IN2(n7116), .IN1(P1_sub_388_n203), 
        .Q(P1_sub_388_n216) );
  NAND2X0 P1_sub_388_U216 ( .IN1(P1_sub_388_n215), .IN2(P1_sub_388_n216), 
        .QN(P1_sub_388_n209) );
  NAND2X0 P1_sub_388_U215 ( .IN1(n7055), .IN2(P1_sub_388_n214), 
        .QN(P1_sub_388_n210) );
  OR2X1 P1_sub_388_U214 ( .IN2(n7055), .IN1(P1_sub_388_n214), 
        .Q(P1_sub_388_n212) );
  INVX0 P1_sub_388_U310 ( .ZN(P1_sub_388_n281), .INP(P1_N2358) );
  NOR2X0 P1_sub_388_U309 ( .QN(P1_sub_388_n277), .IN1(P1_sub_388_n281), 
        .IN2(n7034) );
  INVX0 P1_sub_388_U308 ( .ZN(P1_sub_388_n152), .INP(P1_sub_388_n277) );
  NAND2X0 P1_sub_388_U307 ( .IN1(n7034), .IN2(P1_sub_388_n281), 
        .QN(P1_sub_388_n280) );
  OR2X1 P1_sub_408_U58 ( .IN2(P1_N2759), .IN1(n7117), .Q(P1_sub_408_n66) );
  NAND2X0 P1_sub_408_U57 ( .IN1(P1_N2759), .IN2(n7117), .QN(P1_sub_408_n67) );
  NAND2X0 P1_sub_408_U56 ( .IN1(P1_sub_408_n66), .IN2(P1_sub_408_n67), 
        .QN(P1_sub_408_n60) );
  NAND2X0 P1_sub_408_U55 ( .IN1(P1_N5176), .IN2(P1_sub_408_n65), 
        .QN(P1_sub_408_n61) );
  OR2X1 P1_sub_408_U54 ( .IN2(P1_N5176), .IN1(P1_sub_408_n65), 
        .Q(P1_sub_408_n63) );
  NAND2X0 P1_sub_408_U53 ( .IN1(P1_sub_408_n63), .IN2(P1_sub_408_n64), 
        .QN(P1_sub_408_n62) );
  NAND2X0 P1_sub_408_U52 ( .IN1(P1_sub_408_n61), .IN2(P1_sub_408_n62), 
        .QN(P1_sub_408_n59) );
  NAND2X0 P1_sub_408_U51 ( .IN1(P1_sub_408_n60), .IN2(P1_sub_408_n59), 
        .QN(P1_sub_408_n57) );
  OR2X1 P1_sub_408_U50 ( .IN2(P1_sub_408_n60), .IN1(P1_sub_408_n59), 
        .Q(P1_sub_408_n58) );
  NAND2X0 P1_sub_408_U49 ( .IN1(P1_sub_408_n57), .IN2(P1_sub_408_n58), 
        .QN(P1_N3001) );
  NAND2X0 P1_sub_408_U48 ( .IN1(P1_N5151), .IN2(P1_sub_408_n56), 
        .QN(P1_sub_408_n54) );
  OR2X1 P1_sub_408_U47 ( .IN2(P1_N5151), .IN1(P1_sub_408_n56), 
        .Q(P1_sub_408_n55) );
  NAND2X0 P1_sub_408_U46 ( .IN1(P1_sub_408_n54), .IN2(P1_sub_408_n55), 
        .QN(P1_sub_408_n52) );
  NAND2X0 P1_sub_408_U45 ( .IN1(P1_sub_408_n52), .IN2(P1_sub_408_n53), 
        .QN(P1_sub_408_n50) );
  OR2X1 P1_sub_408_U44 ( .IN2(P1_sub_408_n53), .IN1(P1_sub_408_n52), 
        .Q(P1_sub_408_n51) );
  NAND2X0 P1_sub_408_U43 ( .IN1(P1_sub_408_n50), .IN2(P1_sub_408_n51), 
        .QN(P1_N2975) );
  NAND2X0 P1_sub_408_U42 ( .IN1(n7041), .IN2(P1_sub_408_n49), 
        .QN(P1_sub_408_n47) );
  OR2X1 P1_sub_408_U41 ( .IN2(n7041), .IN1(P1_sub_408_n49), .Q(P1_sub_408_n48)
         );
  NAND2X0 P1_sub_408_U40 ( .IN1(P1_sub_408_n47), .IN2(P1_sub_408_n48), 
        .QN(P1_sub_408_n45) );
  NAND2X0 P1_sub_408_U39 ( .IN1(P1_sub_408_n45), .IN2(P1_sub_408_n46), 
        .QN(P1_sub_408_n43) );
  OR2X1 P1_sub_408_U38 ( .IN2(P1_sub_408_n46), .IN1(P1_sub_408_n45), 
        .Q(P1_sub_408_n44) );
  NAND2X0 P1_sub_408_U37 ( .IN1(P1_sub_408_n43), .IN2(P1_sub_408_n44), 
        .QN(P1_N2976) );
  NAND2X0 P1_sub_408_U36 ( .IN1(n7036), .IN2(P1_sub_408_n42), 
        .QN(P1_sub_408_n40) );
  OR2X1 P1_sub_408_U35 ( .IN2(n7036), .IN1(P1_sub_408_n42), .Q(P1_sub_408_n41)
         );
  NAND2X0 P1_sub_408_U34 ( .IN1(P1_sub_408_n40), .IN2(P1_sub_408_n41), 
        .QN(P1_sub_408_n38) );
  NAND2X0 P1_sub_408_U33 ( .IN1(P1_sub_408_n38), .IN2(P1_sub_408_n39), 
        .QN(P1_sub_408_n36) );
  OR2X1 P1_sub_408_U32 ( .IN2(P1_sub_408_n39), .IN1(P1_sub_408_n38), 
        .Q(P1_sub_408_n37) );
  NAND2X0 P1_sub_408_U31 ( .IN1(P1_sub_408_n36), .IN2(P1_sub_408_n37), 
        .QN(P1_N2977) );
  NAND2X0 P1_sub_408_U30 ( .IN1(n7081), .IN2(P1_sub_408_n35), 
        .QN(P1_sub_408_n33) );
  OR2X1 P1_sub_408_U29 ( .IN2(n7081), .IN1(P1_sub_408_n35), .Q(P1_sub_408_n34)
         );
  NAND2X0 P1_sub_408_U28 ( .IN1(P1_sub_408_n33), .IN2(P1_sub_408_n34), 
        .QN(P1_sub_408_n31) );
  NAND2X0 P1_sub_408_U27 ( .IN1(P1_sub_408_n31), .IN2(P1_sub_408_n32), 
        .QN(P1_sub_408_n29) );
  OR2X1 P1_sub_408_U26 ( .IN2(P1_sub_408_n32), .IN1(P1_sub_408_n31), 
        .Q(P1_sub_408_n30) );
  NAND2X0 P1_sub_408_U25 ( .IN1(P1_sub_408_n29), .IN2(P1_sub_408_n30), 
        .QN(P1_N2978) );
  NAND2X0 P1_sub_408_U24 ( .IN1(n7080), .IN2(P1_sub_408_n28), 
        .QN(P1_sub_408_n26) );
  OR2X1 P1_sub_408_U23 ( .IN2(n7080), .IN1(P1_sub_408_n28), .Q(P1_sub_408_n27)
         );
  NAND2X0 P1_sub_408_U22 ( .IN1(P1_sub_408_n26), .IN2(P1_sub_408_n27), 
        .QN(P1_sub_408_n24) );
  NAND2X0 P1_sub_408_U21 ( .IN1(P1_sub_408_n24), .IN2(P1_sub_408_n25), 
        .QN(P1_sub_408_n22) );
  OR2X1 P1_sub_408_U20 ( .IN2(P1_sub_408_n25), .IN1(P1_sub_408_n24), 
        .Q(P1_sub_408_n23) );
  NAND2X0 P1_sub_408_U19 ( .IN1(P1_sub_408_n22), .IN2(P1_sub_408_n23), 
        .QN(P1_N2979) );
  NAND2X0 P1_sub_408_U18 ( .IN1(n7075), .IN2(P1_sub_408_n21), 
        .QN(P1_sub_408_n19) );
  OR2X1 P1_sub_408_U17 ( .IN2(n7075), .IN1(P1_sub_408_n21), .Q(P1_sub_408_n20)
         );
  NAND2X0 P1_sub_408_U16 ( .IN1(P1_sub_408_n19), .IN2(P1_sub_408_n20), 
        .QN(P1_sub_408_n17) );
  NAND2X0 P1_sub_408_U15 ( .IN1(P1_sub_408_n17), .IN2(P1_sub_408_n18), 
        .QN(P1_sub_408_n15) );
  OR2X1 P1_sub_408_U14 ( .IN2(P1_sub_408_n18), .IN1(P1_sub_408_n17), 
        .Q(P1_sub_408_n16) );
  NAND2X0 P1_sub_408_U13 ( .IN1(P1_sub_408_n15), .IN2(P1_sub_408_n16), 
        .QN(P1_N2980) );
  NAND2X0 P1_sub_408_U12 ( .IN1(P1_N5157), .IN2(P1_sub_408_n14), 
        .QN(P1_sub_408_n12) );
  OR2X1 P1_sub_408_U11 ( .IN2(P1_N5157), .IN1(P1_sub_408_n14), 
        .Q(P1_sub_408_n13) );
  NAND2X0 P1_sub_408_U10 ( .IN1(P1_sub_408_n12), .IN2(P1_sub_408_n13), 
        .QN(P1_sub_408_n10) );
  NAND2X0 P1_sub_408_U9 ( .IN1(P1_sub_408_n10), .IN2(P1_sub_408_n11), 
        .QN(P1_sub_408_n8) );
  OR2X1 P1_sub_408_U8 ( .IN2(P1_sub_408_n11), .IN1(P1_sub_408_n10), 
        .Q(P1_sub_408_n9) );
  NAND2X0 P1_sub_408_U7 ( .IN1(P1_sub_408_n8), .IN2(P1_sub_408_n9), 
        .QN(P1_N2981) );
  NAND2X0 P1_sub_408_U6 ( .IN1(P1_N5158), .IN2(P1_sub_408_n7), 
        .QN(P1_sub_408_n5) );
  OR2X1 P1_sub_408_U5 ( .IN2(P1_N5158), .IN1(P1_sub_408_n7), .Q(P1_sub_408_n6)
         );
  NAND2X0 P1_sub_408_U4 ( .IN1(P1_sub_408_n5), .IN2(P1_sub_408_n6), 
        .QN(P1_sub_408_n3) );
  NAND2X0 P1_sub_408_U3 ( .IN1(P1_sub_408_n3), .IN2(P1_sub_408_n4), 
        .QN(P1_sub_408_n1) );
  OR2X1 P1_sub_408_U2 ( .IN2(P1_sub_408_n4), .IN1(P1_sub_408_n3), 
        .Q(P1_sub_408_n2) );
  NAND2X0 P1_sub_408_U1 ( .IN1(P1_sub_408_n1), .IN2(P1_sub_408_n2), 
        .QN(P1_N2982) );
  NAND2X0 P1_sub_408_U151 ( .IN1(P1_sub_408_n153), .IN2(P1_sub_408_n154), 
        .QN(P1_sub_408_n151) );
  NAND2X0 P1_sub_408_U150 ( .IN1(P1_sub_408_n151), .IN2(P1_sub_408_n152), 
        .QN(P1_sub_408_n149) );
  OR2X1 P1_sub_408_U149 ( .IN2(P1_sub_408_n152), .IN1(P1_sub_408_n151), 
        .Q(P1_sub_408_n150) );
  NAND2X0 P1_sub_408_U148 ( .IN1(P1_sub_408_n149), .IN2(P1_sub_408_n150), 
        .QN(P1_N2974) );
  INVX0 P1_sub_408_U147 ( .ZN(P1_sub_408_n135), .INP(P1_N2751) );
  NAND2X0 P1_sub_408_U146 ( .IN1(n7096), .IN2(P1_sub_408_n135), 
        .QN(P1_sub_408_n147) );
  OR2X1 P1_sub_408_U145 ( .IN2(n7096), .IN1(P1_sub_408_n135), 
        .Q(P1_sub_408_n148) );
  NAND2X0 P1_sub_408_U144 ( .IN1(P1_sub_408_n147), .IN2(P1_sub_408_n148), 
        .QN(P1_sub_408_n141) );
  NAND2X0 P1_sub_408_U143 ( .IN1(P1_N5168), .IN2(P1_sub_408_n146), 
        .QN(P1_sub_408_n142) );
  OR2X1 P1_sub_408_U142 ( .IN2(P1_N5168), .IN1(P1_sub_408_n146), 
        .Q(P1_sub_408_n144) );
  NAND2X0 P1_sub_408_U141 ( .IN1(P1_sub_408_n144), .IN2(P1_sub_408_n145), 
        .QN(P1_sub_408_n143) );
  NAND2X0 P1_sub_408_U140 ( .IN1(P1_sub_408_n142), .IN2(P1_sub_408_n143), 
        .QN(P1_sub_408_n136) );
  NAND2X0 P1_sub_408_U139 ( .IN1(P1_sub_408_n141), .IN2(P1_sub_408_n136), 
        .QN(P1_sub_408_n139) );
  OR2X1 P1_sub_408_U138 ( .IN2(P1_sub_408_n136), .IN1(P1_sub_408_n141), 
        .Q(P1_sub_408_n140) );
  NAND2X0 P1_sub_408_U137 ( .IN1(P1_sub_408_n139), .IN2(P1_sub_408_n140), 
        .QN(P1_N2993) );
  INVX0 P1_sub_408_U136 ( .ZN(P1_sub_408_n125), .INP(P1_N2752) );
  NAND2X0 P1_sub_408_U135 ( .IN1(P1_N5170), .IN2(P1_sub_408_n125), 
        .QN(P1_sub_408_n137) );
  OR2X1 P1_sub_408_U134 ( .IN2(P1_N5170), .IN1(P1_sub_408_n125), 
        .Q(P1_sub_408_n138) );
  NAND2X0 P1_sub_408_U133 ( .IN1(P1_sub_408_n137), .IN2(P1_sub_408_n138), 
        .QN(P1_sub_408_n131) );
  NAND2X0 P1_sub_408_U132 ( .IN1(n7096), .IN2(P1_sub_408_n136), 
        .QN(P1_sub_408_n132) );
  OR2X1 P1_sub_408_U131 ( .IN2(n7096), .IN1(P1_sub_408_n136), 
        .Q(P1_sub_408_n134) );
  NAND2X0 P1_sub_408_U130 ( .IN1(P1_sub_408_n134), .IN2(P1_sub_408_n135), 
        .QN(P1_sub_408_n133) );
  NAND2X0 P1_sub_408_U129 ( .IN1(P1_sub_408_n132), .IN2(P1_sub_408_n133), 
        .QN(P1_sub_408_n126) );
  NAND2X0 P1_sub_408_U128 ( .IN1(P1_sub_408_n131), .IN2(P1_sub_408_n126), 
        .QN(P1_sub_408_n129) );
  OR2X1 P1_sub_408_U127 ( .IN2(P1_sub_408_n126), .IN1(P1_sub_408_n131), 
        .Q(P1_sub_408_n130) );
  NAND2X0 P1_sub_408_U126 ( .IN1(P1_sub_408_n129), .IN2(P1_sub_408_n130), 
        .QN(P1_N2994) );
  INVX0 P1_sub_408_U125 ( .ZN(P1_sub_408_n115), .INP(P1_N2753) );
  NAND2X0 P1_sub_408_U124 ( .IN1(n7089), .IN2(P1_sub_408_n115), 
        .QN(P1_sub_408_n127) );
  OR2X1 P1_sub_408_U123 ( .IN2(n7089), .IN1(P1_sub_408_n115), 
        .Q(P1_sub_408_n128) );
  NAND2X0 P1_sub_408_U122 ( .IN1(P1_sub_408_n127), .IN2(P1_sub_408_n128), 
        .QN(P1_sub_408_n121) );
  NAND2X0 P1_sub_408_U121 ( .IN1(P1_N5170), .IN2(P1_sub_408_n126), 
        .QN(P1_sub_408_n122) );
  OR2X1 P1_sub_408_U120 ( .IN2(P1_N5170), .IN1(P1_sub_408_n126), 
        .Q(P1_sub_408_n124) );
  NAND2X0 P1_sub_408_U119 ( .IN1(P1_sub_408_n124), .IN2(P1_sub_408_n125), 
        .QN(P1_sub_408_n123) );
  NAND2X0 P1_sub_408_U118 ( .IN1(P1_sub_408_n122), .IN2(P1_sub_408_n123), 
        .QN(P1_sub_408_n116) );
  NAND2X0 P1_sub_408_U117 ( .IN1(P1_sub_408_n121), .IN2(P1_sub_408_n116), 
        .QN(P1_sub_408_n119) );
  OR2X1 P1_sub_408_U116 ( .IN2(P1_sub_408_n116), .IN1(P1_sub_408_n121), 
        .Q(P1_sub_408_n120) );
  NAND2X0 P1_sub_408_U115 ( .IN1(P1_sub_408_n119), .IN2(P1_sub_408_n120), 
        .QN(P1_N2995) );
  INVX0 P1_sub_408_U114 ( .ZN(P1_sub_408_n105), .INP(P1_N2754) );
  NAND2X0 P1_sub_408_U113 ( .IN1(P1_N5172), .IN2(P1_sub_408_n105), 
        .QN(P1_sub_408_n117) );
  OR2X1 P1_sub_408_U112 ( .IN2(P1_N5172), .IN1(P1_sub_408_n105), 
        .Q(P1_sub_408_n118) );
  NAND2X0 P1_sub_408_U111 ( .IN1(P1_sub_408_n117), .IN2(P1_sub_408_n118), 
        .QN(P1_sub_408_n111) );
  NAND2X0 P1_sub_408_U110 ( .IN1(n7089), .IN2(P1_sub_408_n116), 
        .QN(P1_sub_408_n112) );
  OR2X1 P1_sub_408_U109 ( .IN2(n7089), .IN1(P1_sub_408_n116), 
        .Q(P1_sub_408_n114) );
  NAND2X0 P1_sub_408_U108 ( .IN1(P1_sub_408_n114), .IN2(P1_sub_408_n115), 
        .QN(P1_sub_408_n113) );
  NAND2X0 P1_sub_408_U107 ( .IN1(P1_sub_408_n112), .IN2(P1_sub_408_n113), 
        .QN(P1_sub_408_n106) );
  NAND2X0 P1_sub_408_U106 ( .IN1(P1_sub_408_n111), .IN2(P1_sub_408_n106), 
        .QN(P1_sub_408_n109) );
  OR2X1 P1_sub_408_U105 ( .IN2(P1_sub_408_n106), .IN1(P1_sub_408_n111), 
        .Q(P1_sub_408_n110) );
  NAND2X0 P1_sub_408_U104 ( .IN1(P1_sub_408_n109), .IN2(P1_sub_408_n110), 
        .QN(P1_N2996) );
  INVX0 P1_sub_408_U103 ( .ZN(P1_sub_408_n95), .INP(P1_N2755) );
  NAND2X0 P1_sub_408_U102 ( .IN1(n7138), .IN2(P1_sub_408_n95), 
        .QN(P1_sub_408_n107) );
  OR2X1 P1_sub_408_U101 ( .IN2(n7138), .IN1(P1_sub_408_n95), 
        .Q(P1_sub_408_n108) );
  NAND2X0 P1_sub_408_U100 ( .IN1(P1_sub_408_n107), .IN2(P1_sub_408_n108), 
        .QN(P1_sub_408_n101) );
  NAND2X0 P1_sub_408_U99 ( .IN1(P1_N5172), .IN2(P1_sub_408_n106), 
        .QN(P1_sub_408_n102) );
  OR2X1 P1_sub_408_U98 ( .IN2(P1_N5172), .IN1(P1_sub_408_n106), 
        .Q(P1_sub_408_n104) );
  NAND2X0 P1_sub_408_U97 ( .IN1(P1_sub_408_n104), .IN2(P1_sub_408_n105), 
        .QN(P1_sub_408_n103) );
  NAND2X0 P1_sub_408_U96 ( .IN1(P1_sub_408_n102), .IN2(P1_sub_408_n103), 
        .QN(P1_sub_408_n96) );
  NAND2X0 P1_sub_408_U95 ( .IN1(P1_sub_408_n101), .IN2(P1_sub_408_n96), 
        .QN(P1_sub_408_n99) );
  OR2X1 P1_sub_408_U94 ( .IN2(P1_sub_408_n96), .IN1(P1_sub_408_n101), 
        .Q(P1_sub_408_n100) );
  NAND2X0 P1_sub_408_U93 ( .IN1(P1_sub_408_n99), .IN2(P1_sub_408_n100), 
        .QN(P1_N2997) );
  INVX0 P1_sub_408_U92 ( .ZN(P1_sub_408_n85), .INP(P1_N2756) );
  NAND2X0 P1_sub_408_U91 ( .IN1(n7129), .IN2(P1_sub_408_n85), 
        .QN(P1_sub_408_n97) );
  OR2X1 P1_sub_408_U90 ( .IN2(n7129), .IN1(P1_sub_408_n85), .Q(P1_sub_408_n98)
         );
  NAND2X0 P1_sub_408_U89 ( .IN1(P1_sub_408_n97), .IN2(P1_sub_408_n98), 
        .QN(P1_sub_408_n91) );
  NAND2X0 P1_sub_408_U88 ( .IN1(n7138), .IN2(P1_sub_408_n96), 
        .QN(P1_sub_408_n92) );
  OR2X1 P1_sub_408_U87 ( .IN2(n7138), .IN1(P1_sub_408_n96), .Q(P1_sub_408_n94)
         );
  NAND2X0 P1_sub_408_U86 ( .IN1(P1_sub_408_n94), .IN2(P1_sub_408_n95), 
        .QN(P1_sub_408_n93) );
  NAND2X0 P1_sub_408_U85 ( .IN1(P1_sub_408_n92), .IN2(P1_sub_408_n93), 
        .QN(P1_sub_408_n86) );
  NAND2X0 P1_sub_408_U84 ( .IN1(P1_sub_408_n91), .IN2(P1_sub_408_n86), 
        .QN(P1_sub_408_n89) );
  OR2X1 P1_sub_408_U83 ( .IN2(P1_sub_408_n86), .IN1(P1_sub_408_n91), 
        .Q(P1_sub_408_n90) );
  NAND2X0 P1_sub_408_U82 ( .IN1(P1_sub_408_n89), .IN2(P1_sub_408_n90), 
        .QN(P1_N2998) );
  INVX0 P1_sub_408_U81 ( .ZN(P1_sub_408_n75), .INP(P1_N2757) );
  NAND2X0 P1_sub_408_U80 ( .IN1(P1_N5175), .IN2(P1_sub_408_n75), 
        .QN(P1_sub_408_n87) );
  OR2X1 P1_sub_408_U79 ( .IN2(P1_N5175), .IN1(P1_sub_408_n75), 
        .Q(P1_sub_408_n88) );
  NAND2X0 P1_sub_408_U78 ( .IN1(P1_sub_408_n87), .IN2(P1_sub_408_n88), 
        .QN(P1_sub_408_n81) );
  NAND2X0 P1_sub_408_U77 ( .IN1(n7129), .IN2(P1_sub_408_n86), 
        .QN(P1_sub_408_n82) );
  OR2X1 P1_sub_408_U76 ( .IN2(n7129), .IN1(P1_sub_408_n86), .Q(P1_sub_408_n84)
         );
  NAND2X0 P1_sub_408_U75 ( .IN1(P1_sub_408_n84), .IN2(P1_sub_408_n85), 
        .QN(P1_sub_408_n83) );
  NAND2X0 P1_sub_408_U74 ( .IN1(P1_sub_408_n82), .IN2(P1_sub_408_n83), 
        .QN(P1_sub_408_n76) );
  NAND2X0 P1_sub_408_U73 ( .IN1(P1_sub_408_n81), .IN2(P1_sub_408_n76), 
        .QN(P1_sub_408_n79) );
  OR2X1 P1_sub_408_U72 ( .IN2(P1_sub_408_n76), .IN1(P1_sub_408_n81), 
        .Q(P1_sub_408_n80) );
  NAND2X0 P1_sub_408_U71 ( .IN1(P1_sub_408_n79), .IN2(P1_sub_408_n80), 
        .QN(P1_N2999) );
  INVX0 P1_sub_408_U70 ( .ZN(P1_sub_408_n64), .INP(P1_N2758) );
  NAND2X0 P1_sub_408_U69 ( .IN1(P1_N5176), .IN2(P1_sub_408_n64), 
        .QN(P1_sub_408_n77) );
  OR2X1 P1_sub_408_U68 ( .IN2(P1_N5176), .IN1(P1_sub_408_n64), 
        .Q(P1_sub_408_n78) );
  NAND2X0 P1_sub_408_U67 ( .IN1(P1_sub_408_n77), .IN2(P1_sub_408_n78), 
        .QN(P1_sub_408_n71) );
  NAND2X0 P1_sub_408_U66 ( .IN1(P1_N5175), .IN2(P1_sub_408_n76), 
        .QN(P1_sub_408_n72) );
  OR2X1 P1_sub_408_U65 ( .IN2(P1_N5175), .IN1(P1_sub_408_n76), 
        .Q(P1_sub_408_n74) );
  NAND2X0 P1_sub_408_U64 ( .IN1(P1_sub_408_n74), .IN2(P1_sub_408_n75), 
        .QN(P1_sub_408_n73) );
  NAND2X0 P1_sub_408_U63 ( .IN1(P1_sub_408_n72), .IN2(P1_sub_408_n73), 
        .QN(P1_sub_408_n65) );
  NAND2X0 P1_sub_408_U62 ( .IN1(P1_sub_408_n71), .IN2(P1_sub_408_n65), 
        .QN(P1_sub_408_n69) );
  OR2X1 P1_sub_408_U61 ( .IN2(P1_sub_408_n65), .IN1(P1_sub_408_n71), 
        .Q(P1_sub_408_n70) );
  NAND2X0 P1_sub_408_U60 ( .IN1(P1_sub_408_n69), .IN2(P1_sub_408_n70), 
        .QN(P1_N3000) );
  NAND2X0 P1_sub_408_U244 ( .IN1(P1_sub_408_n239), .IN2(P1_sub_408_n234), 
        .QN(P1_sub_408_n237) );
  OR2X1 P1_sub_408_U243 ( .IN2(P1_sub_408_n234), .IN1(P1_sub_408_n239), 
        .Q(P1_sub_408_n238) );
  NAND2X0 P1_sub_408_U242 ( .IN1(P1_sub_408_n237), .IN2(P1_sub_408_n238), 
        .QN(P1_N2984) );
  INVX0 P1_sub_408_U241 ( .ZN(P1_sub_408_n223), .INP(P1_N2743) );
  NAND2X0 P1_sub_408_U240 ( .IN1(n7059), .IN2(P1_sub_408_n223), 
        .QN(P1_sub_408_n235) );
  OR2X1 P1_sub_408_U239 ( .IN2(n7059), .IN1(P1_sub_408_n223), 
        .Q(P1_sub_408_n236) );
  NAND2X0 P1_sub_408_U238 ( .IN1(P1_sub_408_n235), .IN2(P1_sub_408_n236), 
        .QN(P1_sub_408_n229) );
  NAND2X0 P1_sub_408_U237 ( .IN1(P1_N5160), .IN2(P1_sub_408_n234), 
        .QN(P1_sub_408_n230) );
  OR2X1 P1_sub_408_U236 ( .IN2(P1_N5160), .IN1(P1_sub_408_n234), 
        .Q(P1_sub_408_n232) );
  NAND2X0 P1_sub_408_U235 ( .IN1(P1_sub_408_n232), .IN2(P1_sub_408_n233), 
        .QN(P1_sub_408_n231) );
  NAND2X0 P1_sub_408_U234 ( .IN1(P1_sub_408_n230), .IN2(P1_sub_408_n231), 
        .QN(P1_sub_408_n224) );
  NAND2X0 P1_sub_408_U233 ( .IN1(P1_sub_408_n229), .IN2(P1_sub_408_n224), 
        .QN(P1_sub_408_n227) );
  OR2X1 P1_sub_408_U232 ( .IN2(P1_sub_408_n224), .IN1(P1_sub_408_n229), 
        .Q(P1_sub_408_n228) );
  NAND2X0 P1_sub_408_U231 ( .IN1(P1_sub_408_n227), .IN2(P1_sub_408_n228), 
        .QN(P1_N2985) );
  INVX0 P1_sub_408_U230 ( .ZN(P1_sub_408_n213), .INP(P1_N2744) );
  NAND2X0 P1_sub_408_U229 ( .IN1(P1_N5162), .IN2(P1_sub_408_n213), 
        .QN(P1_sub_408_n225) );
  OR2X1 P1_sub_408_U228 ( .IN2(P1_N5162), .IN1(P1_sub_408_n213), 
        .Q(P1_sub_408_n226) );
  NAND2X0 P1_sub_408_U227 ( .IN1(P1_sub_408_n225), .IN2(P1_sub_408_n226), 
        .QN(P1_sub_408_n219) );
  NAND2X0 P1_sub_408_U226 ( .IN1(n7059), .IN2(P1_sub_408_n224), 
        .QN(P1_sub_408_n220) );
  OR2X1 P1_sub_408_U225 ( .IN2(n7059), .IN1(P1_sub_408_n224), 
        .Q(P1_sub_408_n222) );
  NAND2X0 P1_sub_408_U224 ( .IN1(P1_sub_408_n222), .IN2(P1_sub_408_n223), 
        .QN(P1_sub_408_n221) );
  NAND2X0 P1_sub_408_U223 ( .IN1(P1_sub_408_n220), .IN2(P1_sub_408_n221), 
        .QN(P1_sub_408_n214) );
  NAND2X0 P1_sub_408_U222 ( .IN1(P1_sub_408_n219), .IN2(P1_sub_408_n214), 
        .QN(P1_sub_408_n217) );
  OR2X1 P1_sub_408_U221 ( .IN2(P1_sub_408_n214), .IN1(P1_sub_408_n219), 
        .Q(P1_sub_408_n218) );
  NAND2X0 P1_sub_408_U220 ( .IN1(P1_sub_408_n217), .IN2(P1_sub_408_n218), 
        .QN(P1_N2986) );
  INVX0 P1_sub_408_U219 ( .ZN(P1_sub_408_n203), .INP(P1_N2745) );
  NAND2X0 P1_sub_408_U218 ( .IN1(n7116), .IN2(P1_sub_408_n203), 
        .QN(P1_sub_408_n215) );
  OR2X1 P1_sub_408_U217 ( .IN2(n7116), .IN1(P1_sub_408_n203), 
        .Q(P1_sub_408_n216) );
  NAND2X0 P1_sub_408_U216 ( .IN1(P1_sub_408_n215), .IN2(P1_sub_408_n216), 
        .QN(P1_sub_408_n209) );
  NAND2X0 P1_sub_408_U215 ( .IN1(P1_N5162), .IN2(P1_sub_408_n214), 
        .QN(P1_sub_408_n210) );
  OR2X1 P1_sub_408_U214 ( .IN2(P1_N5162), .IN1(P1_sub_408_n214), 
        .Q(P1_sub_408_n212) );
  NAND2X0 P1_sub_408_U213 ( .IN1(P1_sub_408_n212), .IN2(P1_sub_408_n213), 
        .QN(P1_sub_408_n211) );
  NAND2X0 P1_sub_408_U212 ( .IN1(P1_sub_408_n210), .IN2(P1_sub_408_n211), 
        .QN(P1_sub_408_n204) );
  NAND2X0 P1_sub_408_U211 ( .IN1(P1_sub_408_n209), .IN2(P1_sub_408_n204), 
        .QN(P1_sub_408_n207) );
  OR2X1 P1_sub_408_U210 ( .IN2(P1_sub_408_n204), .IN1(P1_sub_408_n209), 
        .Q(P1_sub_408_n208) );
  NAND2X0 P1_sub_408_U209 ( .IN1(P1_sub_408_n207), .IN2(P1_sub_408_n208), 
        .QN(P1_N2987) );
  INVX0 P1_sub_408_U208 ( .ZN(P1_sub_408_n193), .INP(P1_N2746) );
  NAND2X0 P1_sub_408_U207 ( .IN1(P1_N5164), .IN2(P1_sub_408_n193), 
        .QN(P1_sub_408_n205) );
  OR2X1 P1_sub_408_U206 ( .IN2(P1_N5164), .IN1(P1_sub_408_n193), 
        .Q(P1_sub_408_n206) );
  NAND2X0 P1_sub_408_U205 ( .IN1(P1_sub_408_n205), .IN2(P1_sub_408_n206), 
        .QN(P1_sub_408_n199) );
  NAND2X0 P1_sub_408_U204 ( .IN1(n7116), .IN2(P1_sub_408_n204), 
        .QN(P1_sub_408_n200) );
  OR2X1 P1_sub_408_U203 ( .IN2(n7116), .IN1(P1_sub_408_n204), 
        .Q(P1_sub_408_n202) );
  NAND2X0 P1_sub_408_U202 ( .IN1(P1_sub_408_n202), .IN2(P1_sub_408_n203), 
        .QN(P1_sub_408_n201) );
  NAND2X0 P1_sub_408_U201 ( .IN1(P1_sub_408_n200), .IN2(P1_sub_408_n201), 
        .QN(P1_sub_408_n194) );
  NAND2X0 P1_sub_408_U200 ( .IN1(P1_sub_408_n199), .IN2(P1_sub_408_n194), 
        .QN(P1_sub_408_n197) );
  OR2X1 P1_sub_408_U199 ( .IN2(P1_sub_408_n194), .IN1(P1_sub_408_n199), 
        .Q(P1_sub_408_n198) );
  NAND2X0 P1_sub_408_U198 ( .IN1(P1_sub_408_n197), .IN2(P1_sub_408_n198), 
        .QN(P1_N2988) );
  INVX0 P1_sub_408_U197 ( .ZN(P1_sub_408_n183), .INP(P1_N2747) );
  NAND2X0 P1_sub_408_U196 ( .IN1(P1_N5165), .IN2(P1_sub_408_n183), 
        .QN(P1_sub_408_n195) );
  OR2X1 P1_sub_408_U195 ( .IN2(P1_N5165), .IN1(P1_sub_408_n183), 
        .Q(P1_sub_408_n196) );
  NAND2X0 P1_sub_408_U194 ( .IN1(P1_sub_408_n195), .IN2(P1_sub_408_n196), 
        .QN(P1_sub_408_n189) );
  NAND2X0 P1_sub_408_U193 ( .IN1(P1_N5164), .IN2(P1_sub_408_n194), 
        .QN(P1_sub_408_n190) );
  OR2X1 P1_sub_408_U192 ( .IN2(P1_N5164), .IN1(P1_sub_408_n194), 
        .Q(P1_sub_408_n192) );
  NAND2X0 P1_sub_408_U191 ( .IN1(P1_sub_408_n192), .IN2(P1_sub_408_n193), 
        .QN(P1_sub_408_n191) );
  NAND2X0 P1_sub_408_U190 ( .IN1(P1_sub_408_n190), .IN2(P1_sub_408_n191), 
        .QN(P1_sub_408_n184) );
  NAND2X0 P1_sub_408_U189 ( .IN1(P1_sub_408_n189), .IN2(P1_sub_408_n184), 
        .QN(P1_sub_408_n187) );
  OR2X1 P1_sub_408_U188 ( .IN2(P1_sub_408_n184), .IN1(P1_sub_408_n189), 
        .Q(P1_sub_408_n188) );
  NAND2X0 P1_sub_408_U187 ( .IN1(P1_sub_408_n187), .IN2(P1_sub_408_n188), 
        .QN(P1_N2989) );
  INVX0 P1_sub_408_U186 ( .ZN(P1_sub_408_n173), .INP(P1_N2748) );
  NAND2X0 P1_sub_408_U185 ( .IN1(n7106), .IN2(P1_sub_408_n173), 
        .QN(P1_sub_408_n185) );
  OR2X1 P1_sub_408_U184 ( .IN2(n7106), .IN1(P1_sub_408_n173), 
        .Q(P1_sub_408_n186) );
  NAND2X0 P1_sub_408_U183 ( .IN1(P1_sub_408_n185), .IN2(P1_sub_408_n186), 
        .QN(P1_sub_408_n179) );
  NAND2X0 P1_sub_408_U182 ( .IN1(P1_N5165), .IN2(P1_sub_408_n184), 
        .QN(P1_sub_408_n180) );
  OR2X1 P1_sub_408_U181 ( .IN2(P1_N5165), .IN1(P1_sub_408_n184), 
        .Q(P1_sub_408_n182) );
  NAND2X0 P1_sub_408_U180 ( .IN1(P1_sub_408_n182), .IN2(P1_sub_408_n183), 
        .QN(P1_sub_408_n181) );
  NAND2X0 P1_sub_408_U179 ( .IN1(P1_sub_408_n180), .IN2(P1_sub_408_n181), 
        .QN(P1_sub_408_n174) );
  NAND2X0 P1_sub_408_U178 ( .IN1(P1_sub_408_n179), .IN2(P1_sub_408_n174), 
        .QN(P1_sub_408_n177) );
  OR2X1 P1_sub_408_U177 ( .IN2(P1_sub_408_n174), .IN1(P1_sub_408_n179), 
        .Q(P1_sub_408_n178) );
  NAND2X0 P1_sub_408_U176 ( .IN1(P1_sub_408_n177), .IN2(P1_sub_408_n178), 
        .QN(P1_N2990) );
  INVX0 P1_sub_408_U175 ( .ZN(P1_sub_408_n163), .INP(P1_N2749) );
  NAND2X0 P1_sub_408_U174 ( .IN1(n7103), .IN2(P1_sub_408_n163), 
        .QN(P1_sub_408_n175) );
  OR2X1 P1_sub_408_U173 ( .IN2(n7103), .IN1(P1_sub_408_n163), 
        .Q(P1_sub_408_n176) );
  NAND2X0 P1_sub_408_U172 ( .IN1(P1_sub_408_n175), .IN2(P1_sub_408_n176), 
        .QN(P1_sub_408_n169) );
  NAND2X0 P1_sub_408_U171 ( .IN1(n7106), .IN2(P1_sub_408_n174), 
        .QN(P1_sub_408_n170) );
  OR2X1 P1_sub_408_U170 ( .IN2(n7106), .IN1(P1_sub_408_n174), 
        .Q(P1_sub_408_n172) );
  NAND2X0 P1_sub_408_U169 ( .IN1(P1_sub_408_n172), .IN2(P1_sub_408_n173), 
        .QN(P1_sub_408_n171) );
  NAND2X0 P1_sub_408_U168 ( .IN1(P1_sub_408_n170), .IN2(P1_sub_408_n171), 
        .QN(P1_sub_408_n164) );
  NAND2X0 P1_sub_408_U167 ( .IN1(P1_sub_408_n169), .IN2(P1_sub_408_n164), 
        .QN(P1_sub_408_n167) );
  OR2X1 P1_sub_408_U166 ( .IN2(P1_sub_408_n164), .IN1(P1_sub_408_n169), 
        .Q(P1_sub_408_n168) );
  NAND2X0 P1_sub_408_U165 ( .IN1(P1_sub_408_n167), .IN2(P1_sub_408_n168), 
        .QN(P1_N2991) );
  INVX0 P1_sub_408_U164 ( .ZN(P1_sub_408_n145), .INP(P1_N2750) );
  NAND2X0 P1_sub_408_U163 ( .IN1(P1_N5168), .IN2(P1_sub_408_n145), 
        .QN(P1_sub_408_n165) );
  OR2X1 P1_sub_408_U162 ( .IN2(P1_N5168), .IN1(P1_sub_408_n145), 
        .Q(P1_sub_408_n166) );
  NAND2X0 P1_sub_408_U161 ( .IN1(P1_sub_408_n165), .IN2(P1_sub_408_n166), 
        .QN(P1_sub_408_n159) );
  NAND2X0 P1_sub_408_U160 ( .IN1(P1_N5167), .IN2(P1_sub_408_n164), 
        .QN(P1_sub_408_n160) );
  OR2X1 P1_sub_408_U159 ( .IN2(n7103), .IN1(P1_sub_408_n164), 
        .Q(P1_sub_408_n162) );
  NAND2X0 P1_sub_408_U158 ( .IN1(P1_sub_408_n162), .IN2(P1_sub_408_n163), 
        .QN(P1_sub_408_n161) );
  NAND2X0 P1_sub_408_U157 ( .IN1(P1_sub_408_n160), .IN2(P1_sub_408_n161), 
        .QN(P1_sub_408_n146) );
  NAND2X0 P1_sub_408_U156 ( .IN1(P1_sub_408_n159), .IN2(P1_sub_408_n146), 
        .QN(P1_sub_408_n157) );
  OR2X1 P1_sub_408_U155 ( .IN2(P1_sub_408_n146), .IN1(P1_sub_408_n159), 
        .Q(P1_sub_408_n158) );
  NAND2X0 P1_sub_408_U154 ( .IN1(P1_sub_408_n157), .IN2(P1_sub_408_n158), 
        .QN(P1_N2992) );
  NAND2X0 P1_sub_408_U153 ( .IN1(P1_N5150), .IN2(P1_sub_408_n156), 
        .QN(P1_sub_408_n153) );
  NAND2X0 P1_sub_408_U152 ( .IN1(P1_N2732), .IN2(n7048), .QN(P1_sub_408_n154)
         );
  INVX0 P1_sub_408_U310 ( .ZN(P1_sub_408_n281), .INP(P1_N2731) );
  NOR2X0 P1_sub_408_U309 ( .QN(P1_sub_408_n277), .IN1(P1_sub_408_n281), 
        .IN2(n7034) );
  INVX0 P1_sub_408_U308 ( .ZN(P1_sub_408_n152), .INP(P1_sub_408_n277) );
  NAND2X0 P1_sub_408_U307 ( .IN1(n7034), .IN2(P1_sub_408_n281), 
        .QN(P1_sub_408_n280) );
  NAND2X0 P1_sub_408_U306 ( .IN1(P1_sub_408_n152), .IN2(P1_sub_408_n280), 
        .QN(P1_N2973) );
  INVX0 P1_sub_408_U305 ( .ZN(P1_sub_408_n243), .INP(P1_N2741) );
  NAND2X0 P1_sub_408_U304 ( .IN1(n7066), .IN2(P1_sub_408_n243), 
        .QN(P1_sub_408_n278) );
  OR2X1 P1_sub_408_U303 ( .IN2(n7066), .IN1(P1_sub_408_n243), 
        .Q(P1_sub_408_n279) );
  NAND2X0 P1_sub_408_U302 ( .IN1(P1_sub_408_n278), .IN2(P1_sub_408_n279), 
        .QN(P1_sub_408_n249) );
  NAND2X0 P1_sub_408_U301 ( .IN1(P1_N5150), .IN2(P1_sub_408_n152), 
        .QN(P1_sub_408_n274) );
  NAND2X0 P1_sub_408_U299 ( .IN1(P1_sub_408_n277), .IN2(n7048), 
        .QN(P1_sub_408_n276) );
  INVX0 P1_sub_408_U298 ( .ZN(P1_sub_408_n156), .INP(P1_N2732) );
  NAND2X0 P1_sub_408_U297 ( .IN1(P1_sub_408_n276), .IN2(P1_sub_408_n156), 
        .QN(P1_sub_408_n275) );
  NAND2X0 P1_sub_408_U296 ( .IN1(P1_sub_408_n274), .IN2(P1_sub_408_n275), 
        .QN(P1_sub_408_n53) );
  NAND2X0 P1_sub_408_U295 ( .IN1(n7046), .IN2(P1_sub_408_n53), 
        .QN(P1_sub_408_n271) );
  OR2X1 P1_sub_408_U294 ( .IN2(n7046), .IN1(P1_sub_408_n53), 
        .Q(P1_sub_408_n273) );
  INVX0 P1_sub_408_U293 ( .ZN(P1_sub_408_n56), .INP(P1_N2733) );
  NAND2X0 P1_sub_408_U292 ( .IN1(P1_sub_408_n273), .IN2(P1_sub_408_n56), 
        .QN(P1_sub_408_n272) );
  NAND2X0 P1_sub_408_U291 ( .IN1(P1_sub_408_n271), .IN2(P1_sub_408_n272), 
        .QN(P1_sub_408_n46) );
  NAND2X0 P1_sub_408_U290 ( .IN1(n7041), .IN2(P1_sub_408_n46), 
        .QN(P1_sub_408_n268) );
  OR2X1 P1_sub_408_U289 ( .IN2(n7041), .IN1(P1_sub_408_n46), 
        .Q(P1_sub_408_n270) );
  INVX0 P1_sub_408_U288 ( .ZN(P1_sub_408_n49), .INP(P1_N2734) );
  NAND2X0 P1_sub_408_U287 ( .IN1(P1_sub_408_n270), .IN2(P1_sub_408_n49), 
        .QN(P1_sub_408_n269) );
  NAND2X0 P1_sub_408_U286 ( .IN1(P1_sub_408_n268), .IN2(P1_sub_408_n269), 
        .QN(P1_sub_408_n39) );
  NAND2X0 P1_sub_408_U285 ( .IN1(n7036), .IN2(P1_sub_408_n39), 
        .QN(P1_sub_408_n265) );
  OR2X1 P1_sub_408_U284 ( .IN2(n7036), .IN1(P1_sub_408_n39), 
        .Q(P1_sub_408_n267) );
  INVX0 P1_sub_408_U283 ( .ZN(P1_sub_408_n42), .INP(P1_N2735) );
  NAND2X0 P1_sub_408_U282 ( .IN1(P1_sub_408_n267), .IN2(P1_sub_408_n42), 
        .QN(P1_sub_408_n266) );
  NAND2X0 P1_sub_408_U281 ( .IN1(P1_sub_408_n265), .IN2(P1_sub_408_n266), 
        .QN(P1_sub_408_n32) );
  NAND2X0 P1_sub_408_U280 ( .IN1(n7081), .IN2(P1_sub_408_n32), 
        .QN(P1_sub_408_n262) );
  OR2X1 P1_sub_408_U279 ( .IN2(n7081), .IN1(P1_sub_408_n32), 
        .Q(P1_sub_408_n264) );
  INVX0 P1_sub_408_U278 ( .ZN(P1_sub_408_n35), .INP(P1_N2736) );
  NAND2X0 P1_sub_408_U277 ( .IN1(P1_sub_408_n264), .IN2(P1_sub_408_n35), 
        .QN(P1_sub_408_n263) );
  NAND2X0 P1_sub_408_U276 ( .IN1(P1_sub_408_n262), .IN2(P1_sub_408_n263), 
        .QN(P1_sub_408_n25) );
  NAND2X0 P1_sub_408_U275 ( .IN1(n7080), .IN2(P1_sub_408_n25), 
        .QN(P1_sub_408_n259) );
  OR2X1 P1_sub_408_U274 ( .IN2(n7080), .IN1(P1_sub_408_n25), 
        .Q(P1_sub_408_n261) );
  INVX0 P1_sub_408_U273 ( .ZN(P1_sub_408_n28), .INP(P1_N2737) );
  NAND2X0 P1_sub_408_U272 ( .IN1(P1_sub_408_n261), .IN2(P1_sub_408_n28), 
        .QN(P1_sub_408_n260) );
  NAND2X0 P1_sub_408_U271 ( .IN1(P1_sub_408_n259), .IN2(P1_sub_408_n260), 
        .QN(P1_sub_408_n18) );
  NAND2X0 P1_sub_408_U270 ( .IN1(n7075), .IN2(P1_sub_408_n18), 
        .QN(P1_sub_408_n256) );
  OR2X1 P1_sub_408_U269 ( .IN2(n7075), .IN1(P1_sub_408_n18), 
        .Q(P1_sub_408_n258) );
  INVX0 P1_sub_408_U268 ( .ZN(P1_sub_408_n21), .INP(P1_N2738) );
  NAND2X0 P1_sub_408_U267 ( .IN1(P1_sub_408_n258), .IN2(P1_sub_408_n21), 
        .QN(P1_sub_408_n257) );
  NAND2X0 P1_sub_408_U266 ( .IN1(P1_sub_408_n256), .IN2(P1_sub_408_n257), 
        .QN(P1_sub_408_n11) );
  NAND2X0 P1_sub_408_U265 ( .IN1(P1_N5157), .IN2(P1_sub_408_n11), 
        .QN(P1_sub_408_n253) );
  OR2X1 P1_sub_408_U264 ( .IN2(P1_N5157), .IN1(P1_sub_408_n11), 
        .Q(P1_sub_408_n255) );
  INVX0 P1_sub_408_U263 ( .ZN(P1_sub_408_n14), .INP(P1_N2739) );
  NAND2X0 P1_sub_408_U262 ( .IN1(P1_sub_408_n255), .IN2(P1_sub_408_n14), 
        .QN(P1_sub_408_n254) );
  NAND2X0 P1_sub_408_U261 ( .IN1(P1_sub_408_n253), .IN2(P1_sub_408_n254), 
        .QN(P1_sub_408_n4) );
  NAND2X0 P1_sub_408_U260 ( .IN1(P1_N5158), .IN2(P1_sub_408_n4), 
        .QN(P1_sub_408_n250) );
  OR2X1 P1_sub_408_U259 ( .IN2(P1_N5158), .IN1(P1_sub_408_n4), 
        .Q(P1_sub_408_n252) );
  INVX0 P1_sub_408_U258 ( .ZN(P1_sub_408_n7), .INP(P1_N2740) );
  NAND2X0 P1_sub_408_U257 ( .IN1(P1_sub_408_n252), .IN2(P1_sub_408_n7), 
        .QN(P1_sub_408_n251) );
  NAND2X0 P1_sub_408_U256 ( .IN1(P1_sub_408_n250), .IN2(P1_sub_408_n251), 
        .QN(P1_sub_408_n244) );
  NAND2X0 P1_sub_408_U255 ( .IN1(P1_sub_408_n249), .IN2(P1_sub_408_n244), 
        .QN(P1_sub_408_n247) );
  OR2X1 P1_sub_408_U254 ( .IN2(P1_sub_408_n244), .IN1(P1_sub_408_n249), 
        .Q(P1_sub_408_n248) );
  NAND2X0 P1_sub_408_U253 ( .IN1(P1_sub_408_n247), .IN2(P1_sub_408_n248), 
        .QN(P1_N2983) );
  INVX0 P1_sub_408_U252 ( .ZN(P1_sub_408_n233), .INP(P1_N2742) );
  NAND2X0 P1_sub_408_U251 ( .IN1(P1_N5160), .IN2(P1_sub_408_n233), 
        .QN(P1_sub_408_n245) );
  OR2X1 P1_sub_408_U250 ( .IN2(P1_N5160), .IN1(P1_sub_408_n233), 
        .Q(P1_sub_408_n246) );
  NAND2X0 P1_sub_408_U249 ( .IN1(P1_sub_408_n245), .IN2(P1_sub_408_n246), 
        .QN(P1_sub_408_n239) );
  NAND2X0 P1_sub_408_U248 ( .IN1(n7066), .IN2(P1_sub_408_n244), 
        .QN(P1_sub_408_n240) );
  OR2X1 P1_sub_408_U247 ( .IN2(n7066), .IN1(P1_sub_408_n244), 
        .Q(P1_sub_408_n242) );
  NAND2X0 P1_sub_408_U246 ( .IN1(P1_sub_408_n242), .IN2(P1_sub_408_n243), 
        .QN(P1_sub_408_n241) );
  NAND2X0 P1_sub_408_U245 ( .IN1(P1_sub_408_n240), .IN2(P1_sub_408_n241), 
        .QN(P1_sub_408_n234) );
  OR2X1 P1_add_428_U88 ( .IN2(n7129), .IN1(P1_add_428_n87), .Q(P1_add_428_n86)
         );
  NAND2X0 P1_add_428_U87 ( .IN1(P1_N3129), .IN2(P1_add_428_n86), 
        .QN(P1_add_428_n85) );
  NAND2X0 P1_add_428_U86 ( .IN1(P1_add_428_n84), .IN2(P1_add_428_n85), 
        .QN(P1_add_428_n77) );
  OR2X1 P1_add_428_U84 ( .IN2(P1_N3130), .IN1(n7125), .Q(P1_add_428_n81) );
  NAND2X0 P1_add_428_U83 ( .IN1(P1_N3130), .IN2(n7125), .QN(P1_add_428_n82) );
  NAND2X0 P1_add_428_U82 ( .IN1(P1_add_428_n81), .IN2(P1_add_428_n82), 
        .QN(P1_add_428_n80) );
  NOR2X0 P1_add_428_U81 ( .QN(P1_add_428_n78), .IN1(P1_add_428_n77), 
        .IN2(P1_add_428_n80) );
  AND2X1 P1_add_428_U80 ( .IN1(P1_add_428_n77), .IN2(P1_add_428_n80), 
        .Q(P1_add_428_n79) );
  NOR2X0 P1_add_428_U79 ( .QN(P1_N3372), .IN1(P1_add_428_n78), 
        .IN2(P1_add_428_n79) );
  NAND2X0 P1_add_428_U78 ( .IN1(P1_N5175), .IN2(P1_add_428_n77), 
        .QN(P1_add_428_n74) );
  OR2X1 P1_add_428_U77 ( .IN2(P1_N5175), .IN1(P1_add_428_n77), 
        .Q(P1_add_428_n76) );
  NAND2X0 P1_add_428_U76 ( .IN1(P1_N3130), .IN2(P1_add_428_n76), 
        .QN(P1_add_428_n75) );
  NAND2X0 P1_add_428_U75 ( .IN1(P1_add_428_n74), .IN2(P1_add_428_n75), 
        .QN(P1_add_428_n64) );
  OR2X1 P1_add_428_U73 ( .IN2(P1_N3131), .IN1(n7119), .Q(P1_add_428_n71) );
  NAND2X0 P1_add_428_U72 ( .IN1(P1_N3131), .IN2(n7119), .QN(P1_add_428_n72) );
  NAND2X0 P1_add_428_U71 ( .IN1(P1_add_428_n71), .IN2(P1_add_428_n72), 
        .QN(P1_add_428_n70) );
  NOR2X0 P1_add_428_U70 ( .QN(P1_add_428_n68), .IN1(P1_add_428_n64), 
        .IN2(P1_add_428_n70) );
  AND2X1 P1_add_428_U69 ( .IN1(P1_add_428_n64), .IN2(P1_add_428_n70), 
        .Q(P1_add_428_n69) );
  NOR2X0 P1_add_428_U68 ( .QN(P1_N3373), .IN1(P1_add_428_n68), 
        .IN2(P1_add_428_n69) );
  OR2X1 P1_add_428_U66 ( .IN2(P1_N3132), .IN1(n7117), .Q(P1_add_428_n65) );
  NAND2X0 P1_add_428_U65 ( .IN1(P1_N3132), .IN2(n7117), .QN(P1_add_428_n66) );
  NAND2X0 P1_add_428_U64 ( .IN1(P1_add_428_n65), .IN2(P1_add_428_n66), 
        .QN(P1_add_428_n60) );
  NAND2X0 P1_add_428_U63 ( .IN1(n7122), .IN2(P1_add_428_n64), 
        .QN(P1_add_428_n61) );
  OR2X1 P1_add_428_U62 ( .IN2(n7122), .IN1(P1_add_428_n64), .Q(P1_add_428_n63)
         );
  NAND2X0 P1_add_428_U61 ( .IN1(P1_N3131), .IN2(P1_add_428_n63), 
        .QN(P1_add_428_n62) );
  NAND2X0 P1_add_428_U60 ( .IN1(P1_add_428_n61), .IN2(P1_add_428_n62), 
        .QN(P1_add_428_n59) );
  NOR2X0 P1_add_428_U59 ( .QN(P1_add_428_n57), .IN1(P1_add_428_n60), 
        .IN2(P1_add_428_n59) );
  AND2X1 P1_add_428_U58 ( .IN1(P1_add_428_n59), .IN2(P1_add_428_n60), 
        .Q(P1_add_428_n58) );
  NOR2X0 P1_add_428_U57 ( .QN(P1_N3374), .IN1(P1_add_428_n57), 
        .IN2(P1_add_428_n58) );
  OR2X1 P1_add_428_U55 ( .IN2(P1_N3106), .IN1(n7045), .Q(P1_add_428_n54) );
  NAND2X0 P1_add_428_U54 ( .IN1(P1_N3106), .IN2(n7045), .QN(P1_add_428_n55) );
  NAND2X0 P1_add_428_U53 ( .IN1(P1_add_428_n54), .IN2(P1_add_428_n55), 
        .QN(P1_add_428_n53) );
  NOR2X0 P1_add_428_U52 ( .QN(P1_add_428_n50), .IN1(P1_add_428_n52), 
        .IN2(P1_add_428_n53) );
  AND2X1 P1_add_428_U51 ( .IN1(P1_add_428_n52), .IN2(P1_add_428_n53), 
        .Q(P1_add_428_n51) );
  NOR2X0 P1_add_428_U50 ( .QN(P1_N3348), .IN1(P1_add_428_n50), 
        .IN2(P1_add_428_n51) );
  OR2X1 P1_add_428_U48 ( .IN2(P1_N3107), .IN1(n7043), .Q(P1_add_428_n47) );
  NAND2X0 P1_add_428_U47 ( .IN1(P1_N3107), .IN2(n7043), .QN(P1_add_428_n48) );
  NAND2X0 P1_add_428_U46 ( .IN1(P1_add_428_n47), .IN2(P1_add_428_n48), 
        .QN(P1_add_428_n46) );
  NOR2X0 P1_add_428_U45 ( .QN(P1_add_428_n43), .IN1(P1_add_428_n45), 
        .IN2(P1_add_428_n46) );
  AND2X1 P1_add_428_U44 ( .IN1(P1_add_428_n45), .IN2(P1_add_428_n46), 
        .Q(P1_add_428_n44) );
  NOR2X0 P1_add_428_U43 ( .QN(P1_N3349), .IN1(P1_add_428_n43), 
        .IN2(P1_add_428_n44) );
  OR2X1 P1_add_428_U41 ( .IN2(P1_N3108), .IN1(n7037), .Q(P1_add_428_n40) );
  NAND2X0 P1_add_428_U40 ( .IN1(P1_N3108), .IN2(n7037), .QN(P1_add_428_n41) );
  NAND2X0 P1_add_428_U39 ( .IN1(P1_add_428_n40), .IN2(P1_add_428_n41), 
        .QN(P1_add_428_n39) );
  NOR2X0 P1_add_428_U38 ( .QN(P1_add_428_n36), .IN1(P1_add_428_n38), 
        .IN2(P1_add_428_n39) );
  AND2X1 P1_add_428_U37 ( .IN1(P1_add_428_n38), .IN2(P1_add_428_n39), 
        .Q(P1_add_428_n37) );
  NOR2X0 P1_add_428_U36 ( .QN(P1_N3350), .IN1(P1_add_428_n36), 
        .IN2(P1_add_428_n37) );
  OR2X1 P1_add_428_U34 ( .IN2(P1_N3109), .IN1(n7082), .Q(P1_add_428_n33) );
  NAND2X0 P1_add_428_U33 ( .IN1(P1_N3109), .IN2(n7082), .QN(P1_add_428_n34) );
  NAND2X0 P1_add_428_U32 ( .IN1(P1_add_428_n33), .IN2(P1_add_428_n34), 
        .QN(P1_add_428_n32) );
  NOR2X0 P1_add_428_U31 ( .QN(P1_add_428_n29), .IN1(P1_add_428_n31), 
        .IN2(P1_add_428_n32) );
  AND2X1 P1_add_428_U30 ( .IN1(P1_add_428_n31), .IN2(P1_add_428_n32), 
        .Q(P1_add_428_n30) );
  NOR2X0 P1_add_428_U29 ( .QN(P1_N3351), .IN1(P1_add_428_n29), 
        .IN2(P1_add_428_n30) );
  OR2X1 P1_add_428_U27 ( .IN2(P1_N3110), .IN1(n7079), .Q(P1_add_428_n26) );
  NAND2X0 P1_add_428_U26 ( .IN1(P1_N3110), .IN2(n7079), .QN(P1_add_428_n27) );
  NAND2X0 P1_add_428_U25 ( .IN1(P1_add_428_n26), .IN2(P1_add_428_n27), 
        .QN(P1_add_428_n25) );
  NOR2X0 P1_add_428_U24 ( .QN(P1_add_428_n22), .IN1(P1_add_428_n24), 
        .IN2(P1_add_428_n25) );
  AND2X1 P1_add_428_U23 ( .IN1(P1_add_428_n24), .IN2(P1_add_428_n25), 
        .Q(P1_add_428_n23) );
  NOR2X0 P1_add_428_U22 ( .QN(P1_N3352), .IN1(P1_add_428_n22), 
        .IN2(P1_add_428_n23) );
  OR2X1 P1_add_428_U20 ( .IN2(P1_N3111), .IN1(n7076), .Q(P1_add_428_n19) );
  NAND2X0 P1_add_428_U19 ( .IN1(P1_N3111), .IN2(n7076), .QN(P1_add_428_n20) );
  NAND2X0 P1_add_428_U18 ( .IN1(P1_add_428_n19), .IN2(P1_add_428_n20), 
        .QN(P1_add_428_n18) );
  NOR2X0 P1_add_428_U17 ( .QN(P1_add_428_n15), .IN1(P1_add_428_n17), 
        .IN2(P1_add_428_n18) );
  AND2X1 P1_add_428_U16 ( .IN1(P1_add_428_n17), .IN2(P1_add_428_n18), 
        .Q(P1_add_428_n16) );
  NOR2X0 P1_add_428_U15 ( .QN(P1_N3353), .IN1(P1_add_428_n15), 
        .IN2(P1_add_428_n16) );
  OR2X1 P1_add_428_U13 ( .IN2(P1_N3112), .IN1(n7073), .Q(P1_add_428_n12) );
  NAND2X0 P1_add_428_U12 ( .IN1(P1_N3112), .IN2(n7073), .QN(P1_add_428_n13) );
  NAND2X0 P1_add_428_U11 ( .IN1(P1_add_428_n12), .IN2(P1_add_428_n13), 
        .QN(P1_add_428_n11) );
  NOR2X0 P1_add_428_U10 ( .QN(P1_add_428_n8), .IN1(P1_add_428_n10), 
        .IN2(P1_add_428_n11) );
  AND2X1 P1_add_428_U9 ( .IN1(P1_add_428_n10), .IN2(P1_add_428_n11), 
        .Q(P1_add_428_n9) );
  NOR2X0 P1_add_428_U8 ( .QN(P1_N3354), .IN1(P1_add_428_n8), 
        .IN2(P1_add_428_n9) );
  OR2X1 P1_add_428_U6 ( .IN2(P1_N3113), .IN1(n7071), .Q(P1_add_428_n5) );
  NAND2X0 P1_add_428_U5 ( .IN1(P1_N3113), .IN2(n7071), .QN(P1_add_428_n6) );
  NAND2X0 P1_add_428_U4 ( .IN1(P1_add_428_n5), .IN2(P1_add_428_n6), 
        .QN(P1_add_428_n4) );
  NOR2X0 P1_add_428_U3 ( .QN(P1_add_428_n1), .IN1(P1_add_428_n3), 
        .IN2(P1_add_428_n4) );
  AND2X1 P1_add_428_U2 ( .IN1(P1_add_428_n3), .IN2(P1_add_428_n4), 
        .Q(P1_add_428_n2) );
  NOR2X0 P1_add_428_U1 ( .QN(P1_N3355), .IN1(P1_add_428_n1), 
        .IN2(P1_add_428_n2) );
  NAND2X0 P1_add_428_U181 ( .IN1(P1_N3121), .IN2(P1_add_428_n173), 
        .QN(P1_add_428_n172) );
  NAND2X0 P1_add_428_U180 ( .IN1(P1_add_428_n171), .IN2(P1_add_428_n172), 
        .QN(P1_add_428_n164) );
  OR2X1 P1_add_428_U178 ( .IN2(P1_N3122), .IN1(n7102), .Q(P1_add_428_n168) );
  NAND2X0 P1_add_428_U177 ( .IN1(P1_N3122), .IN2(n7102), .QN(P1_add_428_n169)
         );
  NAND2X0 P1_add_428_U176 ( .IN1(P1_add_428_n168), .IN2(P1_add_428_n169), 
        .QN(P1_add_428_n167) );
  NOR2X0 P1_add_428_U175 ( .QN(P1_add_428_n165), .IN1(P1_add_428_n164), 
        .IN2(P1_add_428_n167) );
  AND2X1 P1_add_428_U174 ( .IN1(P1_add_428_n164), .IN2(P1_add_428_n167), 
        .Q(P1_add_428_n166) );
  NOR2X0 P1_add_428_U173 ( .QN(P1_N3364), .IN1(P1_add_428_n165), 
        .IN2(P1_add_428_n166) );
  NAND2X0 P1_add_428_U172 ( .IN1(P1_N5167), .IN2(P1_add_428_n164), 
        .QN(P1_add_428_n161) );
  OR2X1 P1_add_428_U171 ( .IN2(P1_N5167), .IN1(P1_add_428_n164), 
        .Q(P1_add_428_n163) );
  NAND2X0 P1_add_428_U170 ( .IN1(P1_N3122), .IN2(P1_add_428_n163), 
        .QN(P1_add_428_n162) );
  NAND2X0 P1_add_428_U169 ( .IN1(P1_add_428_n161), .IN2(P1_add_428_n162), 
        .QN(P1_add_428_n147) );
  OR2X1 P1_add_428_U167 ( .IN2(P1_N3123), .IN1(n7098), .Q(P1_add_428_n158) );
  NAND2X0 P1_add_428_U166 ( .IN1(P1_N3123), .IN2(n7098), .QN(P1_add_428_n159)
         );
  NAND2X0 P1_add_428_U165 ( .IN1(P1_add_428_n158), .IN2(P1_add_428_n159), 
        .QN(P1_add_428_n157) );
  NOR2X0 P1_add_428_U164 ( .QN(P1_add_428_n155), .IN1(P1_add_428_n147), 
        .IN2(P1_add_428_n157) );
  AND2X1 P1_add_428_U163 ( .IN1(P1_add_428_n147), .IN2(P1_add_428_n157), 
        .Q(P1_add_428_n156) );
  NOR2X0 P1_add_428_U162 ( .QN(P1_N3365), .IN1(P1_add_428_n155), 
        .IN2(P1_add_428_n156) );
  OR2X1 P1_add_428_U161 ( .IN2(P1_N3105), .IN1(n7051), .Q(P1_add_428_n152) );
  NAND2X0 P1_add_428_U160 ( .IN1(P1_N3105), .IN2(n7051), .QN(P1_add_428_n153)
         );
  NAND2X0 P1_add_428_U159 ( .IN1(P1_add_428_n152), .IN2(P1_add_428_n153), 
        .QN(P1_add_428_n150) );
  NAND2X0 P1_add_428_U158 ( .IN1(P1_add_428_n150), .IN2(P1_add_428_n151), 
        .QN(P1_add_428_n148) );
  OR2X1 P1_add_428_U157 ( .IN2(P1_add_428_n151), .IN1(P1_add_428_n150), 
        .Q(P1_add_428_n149) );
  NAND2X0 P1_add_428_U156 ( .IN1(P1_add_428_n148), .IN2(P1_add_428_n149), 
        .QN(P1_N3347) );
  NAND2X0 P1_add_428_U155 ( .IN1(n7099), .IN2(P1_add_428_n147), 
        .QN(P1_add_428_n144) );
  OR2X1 P1_add_428_U154 ( .IN2(n7099), .IN1(P1_add_428_n147), 
        .Q(P1_add_428_n146) );
  NAND2X0 P1_add_428_U153 ( .IN1(P1_N3123), .IN2(P1_add_428_n146), 
        .QN(P1_add_428_n145) );
  NAND2X0 P1_add_428_U152 ( .IN1(P1_add_428_n144), .IN2(P1_add_428_n145), 
        .QN(P1_add_428_n137) );
  OR2X1 P1_add_428_U150 ( .IN2(P1_N3124), .IN1(n7095), .Q(P1_add_428_n141) );
  NAND2X0 P1_add_428_U149 ( .IN1(P1_N3124), .IN2(n7095), .QN(P1_add_428_n142)
         );
  NAND2X0 P1_add_428_U148 ( .IN1(P1_add_428_n141), .IN2(P1_add_428_n142), 
        .QN(P1_add_428_n140) );
  NOR2X0 P1_add_428_U147 ( .QN(P1_add_428_n138), .IN1(P1_add_428_n137), 
        .IN2(P1_add_428_n140) );
  AND2X1 P1_add_428_U146 ( .IN1(P1_add_428_n137), .IN2(P1_add_428_n140), 
        .Q(P1_add_428_n139) );
  NOR2X0 P1_add_428_U145 ( .QN(P1_N3366), .IN1(P1_add_428_n138), 
        .IN2(P1_add_428_n139) );
  NAND2X0 P1_add_428_U144 ( .IN1(P1_N5169), .IN2(P1_add_428_n137), 
        .QN(P1_add_428_n134) );
  OR2X1 P1_add_428_U143 ( .IN2(P1_N5169), .IN1(P1_add_428_n137), 
        .Q(P1_add_428_n136) );
  NAND2X0 P1_add_428_U142 ( .IN1(P1_N3124), .IN2(P1_add_428_n136), 
        .QN(P1_add_428_n135) );
  NAND2X0 P1_add_428_U141 ( .IN1(P1_add_428_n134), .IN2(P1_add_428_n135), 
        .QN(P1_add_428_n127) );
  OR2X1 P1_add_428_U139 ( .IN2(P1_N3125), .IN1(n7092), .Q(P1_add_428_n131) );
  NAND2X0 P1_add_428_U138 ( .IN1(P1_N3125), .IN2(n7092), .QN(P1_add_428_n132)
         );
  NAND2X0 P1_add_428_U137 ( .IN1(P1_add_428_n131), .IN2(P1_add_428_n132), 
        .QN(P1_add_428_n130) );
  NOR2X0 P1_add_428_U136 ( .QN(P1_add_428_n128), .IN1(P1_add_428_n127), 
        .IN2(P1_add_428_n130) );
  AND2X1 P1_add_428_U135 ( .IN1(P1_add_428_n127), .IN2(P1_add_428_n130), 
        .Q(P1_add_428_n129) );
  NOR2X0 P1_add_428_U134 ( .QN(P1_N3367), .IN1(P1_add_428_n128), 
        .IN2(P1_add_428_n129) );
  NAND2X0 P1_add_428_U133 ( .IN1(n7093), .IN2(P1_add_428_n127), 
        .QN(P1_add_428_n124) );
  OR2X1 P1_add_428_U132 ( .IN2(n7093), .IN1(P1_add_428_n127), 
        .Q(P1_add_428_n126) );
  NAND2X0 P1_add_428_U131 ( .IN1(P1_N3125), .IN2(P1_add_428_n126), 
        .QN(P1_add_428_n125) );
  NAND2X0 P1_add_428_U130 ( .IN1(P1_add_428_n124), .IN2(P1_add_428_n125), 
        .QN(P1_add_428_n117) );
  OR2X1 P1_add_428_U128 ( .IN2(P1_N3126), .IN1(n7090), .Q(P1_add_428_n121) );
  NAND2X0 P1_add_428_U127 ( .IN1(P1_N3126), .IN2(n7090), .QN(P1_add_428_n122)
         );
  NAND2X0 P1_add_428_U126 ( .IN1(P1_add_428_n121), .IN2(P1_add_428_n122), 
        .QN(P1_add_428_n120) );
  NOR2X0 P1_add_428_U125 ( .QN(P1_add_428_n118), .IN1(P1_add_428_n117), 
        .IN2(P1_add_428_n120) );
  AND2X1 P1_add_428_U124 ( .IN1(P1_add_428_n117), .IN2(P1_add_428_n120), 
        .Q(P1_add_428_n119) );
  NOR2X0 P1_add_428_U123 ( .QN(P1_N3368), .IN1(P1_add_428_n118), 
        .IN2(P1_add_428_n119) );
  NAND2X0 P1_add_428_U122 ( .IN1(P1_N5171), .IN2(P1_add_428_n117), 
        .QN(P1_add_428_n114) );
  OR2X1 P1_add_428_U121 ( .IN2(P1_N5171), .IN1(P1_add_428_n117), 
        .Q(P1_add_428_n116) );
  NAND2X0 P1_add_428_U120 ( .IN1(P1_N3126), .IN2(P1_add_428_n116), 
        .QN(P1_add_428_n115) );
  NAND2X0 P1_add_428_U119 ( .IN1(P1_add_428_n114), .IN2(P1_add_428_n115), 
        .QN(P1_add_428_n107) );
  OR2X1 P1_add_428_U117 ( .IN2(P1_N3127), .IN1(n7144), .Q(P1_add_428_n111) );
  NAND2X0 P1_add_428_U116 ( .IN1(P1_N3127), .IN2(n7144), .QN(P1_add_428_n112)
         );
  NAND2X0 P1_add_428_U115 ( .IN1(P1_add_428_n111), .IN2(P1_add_428_n112), 
        .QN(P1_add_428_n110) );
  NOR2X0 P1_add_428_U114 ( .QN(P1_add_428_n108), .IN1(P1_add_428_n107), 
        .IN2(P1_add_428_n110) );
  AND2X1 P1_add_428_U113 ( .IN1(P1_add_428_n107), .IN2(P1_add_428_n110), 
        .Q(P1_add_428_n109) );
  NOR2X0 P1_add_428_U112 ( .QN(P1_N3369), .IN1(P1_add_428_n108), 
        .IN2(P1_add_428_n109) );
  NAND2X0 P1_add_428_U111 ( .IN1(n7141), .IN2(P1_add_428_n107), 
        .QN(P1_add_428_n104) );
  OR2X1 P1_add_428_U110 ( .IN2(n7141), .IN1(P1_add_428_n107), 
        .Q(P1_add_428_n106) );
  NAND2X0 P1_add_428_U109 ( .IN1(P1_N3127), .IN2(P1_add_428_n106), 
        .QN(P1_add_428_n105) );
  NAND2X0 P1_add_428_U108 ( .IN1(P1_add_428_n104), .IN2(P1_add_428_n105), 
        .QN(P1_add_428_n97) );
  OR2X1 P1_add_428_U106 ( .IN2(P1_N3128), .IN1(n7136), .Q(P1_add_428_n101) );
  NAND2X0 P1_add_428_U105 ( .IN1(P1_N3128), .IN2(n7136), .QN(P1_add_428_n102)
         );
  NAND2X0 P1_add_428_U104 ( .IN1(P1_add_428_n101), .IN2(P1_add_428_n102), 
        .QN(P1_add_428_n100) );
  NOR2X0 P1_add_428_U103 ( .QN(P1_add_428_n98), .IN1(P1_add_428_n97), 
        .IN2(P1_add_428_n100) );
  AND2X1 P1_add_428_U102 ( .IN1(P1_add_428_n97), .IN2(P1_add_428_n100), 
        .Q(P1_add_428_n99) );
  NOR2X0 P1_add_428_U101 ( .QN(P1_N3370), .IN1(P1_add_428_n98), 
        .IN2(P1_add_428_n99) );
  NAND2X0 P1_add_428_U100 ( .IN1(P1_N5173), .IN2(P1_add_428_n97), 
        .QN(P1_add_428_n94) );
  OR2X1 P1_add_428_U99 ( .IN2(P1_N5173), .IN1(P1_add_428_n97), 
        .Q(P1_add_428_n96) );
  NAND2X0 P1_add_428_U98 ( .IN1(P1_N3128), .IN2(P1_add_428_n96), 
        .QN(P1_add_428_n95) );
  NAND2X0 P1_add_428_U97 ( .IN1(P1_add_428_n94), .IN2(P1_add_428_n95), 
        .QN(P1_add_428_n87) );
  OR2X1 P1_add_428_U95 ( .IN2(P1_N3129), .IN1(n7130), .Q(P1_add_428_n91) );
  NAND2X0 P1_add_428_U94 ( .IN1(P1_N3129), .IN2(n7130), .QN(P1_add_428_n92) );
  NAND2X0 P1_add_428_U93 ( .IN1(P1_add_428_n91), .IN2(P1_add_428_n92), 
        .QN(P1_add_428_n90) );
  NOR2X0 P1_add_428_U92 ( .QN(P1_add_428_n88), .IN1(P1_add_428_n87), 
        .IN2(P1_add_428_n90) );
  AND2X1 P1_add_428_U91 ( .IN1(P1_add_428_n87), .IN2(P1_add_428_n90), 
        .Q(P1_add_428_n89) );
  NOR2X0 P1_add_428_U90 ( .QN(P1_N3371), .IN1(P1_add_428_n88), 
        .IN2(P1_add_428_n89) );
  NAND2X0 P1_add_428_U89 ( .IN1(n7129), .IN2(P1_add_428_n87), 
        .QN(P1_add_428_n84) );
  OR2X1 P1_add_428_U274 ( .IN2(n7072), .IN1(P1_add_428_n10), 
        .Q(P1_add_428_n256) );
  NAND2X0 P1_add_428_U273 ( .IN1(P1_N3112), .IN2(P1_add_428_n256), 
        .QN(P1_add_428_n255) );
  NAND2X0 P1_add_428_U272 ( .IN1(P1_add_428_n254), .IN2(P1_add_428_n255), 
        .QN(P1_add_428_n3) );
  NAND2X0 P1_add_428_U271 ( .IN1(P1_N5158), .IN2(P1_add_428_n3), 
        .QN(P1_add_428_n251) );
  OR2X1 P1_add_428_U270 ( .IN2(P1_N5158), .IN1(P1_add_428_n3), 
        .Q(P1_add_428_n253) );
  NAND2X0 P1_add_428_U269 ( .IN1(P1_N3113), .IN2(P1_add_428_n253), 
        .QN(P1_add_428_n252) );
  NAND2X0 P1_add_428_U268 ( .IN1(P1_add_428_n251), .IN2(P1_add_428_n252), 
        .QN(P1_add_428_n244) );
  OR2X1 P1_add_428_U266 ( .IN2(P1_N3114), .IN1(n7067), .Q(P1_add_428_n248) );
  NAND2X0 P1_add_428_U265 ( .IN1(P1_N3114), .IN2(n7067), .QN(P1_add_428_n249)
         );
  NAND2X0 P1_add_428_U264 ( .IN1(P1_add_428_n248), .IN2(P1_add_428_n249), 
        .QN(P1_add_428_n247) );
  NOR2X0 P1_add_428_U263 ( .QN(P1_add_428_n245), .IN1(P1_add_428_n244), 
        .IN2(P1_add_428_n247) );
  AND2X1 P1_add_428_U262 ( .IN1(P1_add_428_n244), .IN2(P1_add_428_n247), 
        .Q(P1_add_428_n246) );
  NOR2X0 P1_add_428_U261 ( .QN(P1_N3356), .IN1(P1_add_428_n245), 
        .IN2(P1_add_428_n246) );
  NAND2X0 P1_add_428_U260 ( .IN1(P1_N5159), .IN2(P1_add_428_n244), 
        .QN(P1_add_428_n241) );
  OR2X1 P1_add_428_U259 ( .IN2(P1_N5159), .IN1(P1_add_428_n244), 
        .Q(P1_add_428_n243) );
  NAND2X0 P1_add_428_U258 ( .IN1(P1_N3114), .IN2(P1_add_428_n243), 
        .QN(P1_add_428_n242) );
  NAND2X0 P1_add_428_U257 ( .IN1(P1_add_428_n241), .IN2(P1_add_428_n242), 
        .QN(P1_add_428_n234) );
  OR2X1 P1_add_428_U255 ( .IN2(P1_N3115), .IN1(n7063), .Q(P1_add_428_n238) );
  NAND2X0 P1_add_428_U254 ( .IN1(P1_N3115), .IN2(n7063), .QN(P1_add_428_n239)
         );
  NAND2X0 P1_add_428_U253 ( .IN1(P1_add_428_n238), .IN2(P1_add_428_n239), 
        .QN(P1_add_428_n237) );
  NOR2X0 P1_add_428_U252 ( .QN(P1_add_428_n235), .IN1(P1_add_428_n234), 
        .IN2(P1_add_428_n237) );
  AND2X1 P1_add_428_U251 ( .IN1(P1_add_428_n234), .IN2(P1_add_428_n237), 
        .Q(P1_add_428_n236) );
  NOR2X0 P1_add_428_U250 ( .QN(P1_N3357), .IN1(P1_add_428_n235), 
        .IN2(P1_add_428_n236) );
  NAND2X0 P1_add_428_U249 ( .IN1(P1_N5160), .IN2(P1_add_428_n234), 
        .QN(P1_add_428_n231) );
  OR2X1 P1_add_428_U248 ( .IN2(P1_N5160), .IN1(P1_add_428_n234), 
        .Q(P1_add_428_n233) );
  NAND2X0 P1_add_428_U247 ( .IN1(P1_N3115), .IN2(P1_add_428_n233), 
        .QN(P1_add_428_n232) );
  NAND2X0 P1_add_428_U246 ( .IN1(P1_add_428_n231), .IN2(P1_add_428_n232), 
        .QN(P1_add_428_n224) );
  OR2X1 P1_add_428_U244 ( .IN2(P1_N3116), .IN1(n7058), .Q(P1_add_428_n228) );
  NAND2X0 P1_add_428_U243 ( .IN1(P1_N3116), .IN2(n7058), .QN(P1_add_428_n229)
         );
  NAND2X0 P1_add_428_U242 ( .IN1(P1_add_428_n228), .IN2(P1_add_428_n229), 
        .QN(P1_add_428_n227) );
  NOR2X0 P1_add_428_U241 ( .QN(P1_add_428_n225), .IN1(P1_add_428_n224), 
        .IN2(P1_add_428_n227) );
  AND2X1 P1_add_428_U240 ( .IN1(P1_add_428_n224), .IN2(P1_add_428_n227), 
        .Q(P1_add_428_n226) );
  NOR2X0 P1_add_428_U239 ( .QN(P1_N3358), .IN1(P1_add_428_n225), 
        .IN2(P1_add_428_n226) );
  NAND2X0 P1_add_428_U238 ( .IN1(P1_N5161), .IN2(P1_add_428_n224), 
        .QN(P1_add_428_n221) );
  OR2X1 P1_add_428_U237 ( .IN2(P1_N5161), .IN1(P1_add_428_n224), 
        .Q(P1_add_428_n223) );
  NAND2X0 P1_add_428_U236 ( .IN1(P1_N3116), .IN2(P1_add_428_n223), 
        .QN(P1_add_428_n222) );
  NAND2X0 P1_add_428_U235 ( .IN1(P1_add_428_n221), .IN2(P1_add_428_n222), 
        .QN(P1_add_428_n214) );
  OR2X1 P1_add_428_U233 ( .IN2(P1_N3117), .IN1(n7056), .Q(P1_add_428_n218) );
  NAND2X0 P1_add_428_U232 ( .IN1(P1_N3117), .IN2(n7056), .QN(P1_add_428_n219)
         );
  NAND2X0 P1_add_428_U231 ( .IN1(P1_add_428_n218), .IN2(P1_add_428_n219), 
        .QN(P1_add_428_n217) );
  NOR2X0 P1_add_428_U230 ( .QN(P1_add_428_n215), .IN1(P1_add_428_n214), 
        .IN2(P1_add_428_n217) );
  AND2X1 P1_add_428_U229 ( .IN1(P1_add_428_n214), .IN2(P1_add_428_n217), 
        .Q(P1_add_428_n216) );
  NOR2X0 P1_add_428_U228 ( .QN(P1_N3359), .IN1(P1_add_428_n215), 
        .IN2(P1_add_428_n216) );
  NAND2X0 P1_add_428_U227 ( .IN1(P1_N5162), .IN2(P1_add_428_n214), 
        .QN(P1_add_428_n211) );
  OR2X1 P1_add_428_U226 ( .IN2(P1_N5162), .IN1(P1_add_428_n214), 
        .Q(P1_add_428_n213) );
  NAND2X0 P1_add_428_U225 ( .IN1(P1_N3117), .IN2(P1_add_428_n213), 
        .QN(P1_add_428_n212) );
  NAND2X0 P1_add_428_U224 ( .IN1(P1_add_428_n211), .IN2(P1_add_428_n212), 
        .QN(P1_add_428_n204) );
  OR2X1 P1_add_428_U222 ( .IN2(P1_N3118), .IN1(n7115), .Q(P1_add_428_n208) );
  NAND2X0 P1_add_428_U221 ( .IN1(P1_N3118), .IN2(n7115), .QN(P1_add_428_n209)
         );
  NAND2X0 P1_add_428_U220 ( .IN1(P1_add_428_n208), .IN2(P1_add_428_n209), 
        .QN(P1_add_428_n207) );
  NOR2X0 P1_add_428_U219 ( .QN(P1_add_428_n205), .IN1(P1_add_428_n204), 
        .IN2(P1_add_428_n207) );
  AND2X1 P1_add_428_U218 ( .IN1(P1_add_428_n204), .IN2(P1_add_428_n207), 
        .Q(P1_add_428_n206) );
  NOR2X0 P1_add_428_U217 ( .QN(P1_N3360), .IN1(P1_add_428_n205), 
        .IN2(P1_add_428_n206) );
  NAND2X0 P1_add_428_U216 ( .IN1(n7116), .IN2(P1_add_428_n204), 
        .QN(P1_add_428_n201) );
  OR2X1 P1_add_428_U215 ( .IN2(n7116), .IN1(P1_add_428_n204), 
        .Q(P1_add_428_n203) );
  NAND2X0 P1_add_428_U214 ( .IN1(P1_N3118), .IN2(P1_add_428_n203), 
        .QN(P1_add_428_n202) );
  NAND2X0 P1_add_428_U213 ( .IN1(P1_add_428_n201), .IN2(P1_add_428_n202), 
        .QN(P1_add_428_n194) );
  OR2X1 P1_add_428_U211 ( .IN2(P1_N3119), .IN1(n7112), .Q(P1_add_428_n198) );
  NAND2X0 P1_add_428_U210 ( .IN1(P1_N3119), .IN2(n7112), .QN(P1_add_428_n199)
         );
  NAND2X0 P1_add_428_U209 ( .IN1(P1_add_428_n198), .IN2(P1_add_428_n199), 
        .QN(P1_add_428_n197) );
  NOR2X0 P1_add_428_U208 ( .QN(P1_add_428_n195), .IN1(P1_add_428_n194), 
        .IN2(P1_add_428_n197) );
  AND2X1 P1_add_428_U207 ( .IN1(P1_add_428_n194), .IN2(P1_add_428_n197), 
        .Q(P1_add_428_n196) );
  NOR2X0 P1_add_428_U206 ( .QN(P1_N3361), .IN1(P1_add_428_n195), 
        .IN2(P1_add_428_n196) );
  NAND2X0 P1_add_428_U205 ( .IN1(P1_N5164), .IN2(P1_add_428_n194), 
        .QN(P1_add_428_n191) );
  OR2X1 P1_add_428_U204 ( .IN2(P1_N5164), .IN1(P1_add_428_n194), 
        .Q(P1_add_428_n193) );
  NAND2X0 P1_add_428_U203 ( .IN1(P1_N3119), .IN2(P1_add_428_n193), 
        .QN(P1_add_428_n192) );
  NAND2X0 P1_add_428_U202 ( .IN1(P1_add_428_n191), .IN2(P1_add_428_n192), 
        .QN(P1_add_428_n184) );
  OR2X1 P1_add_428_U200 ( .IN2(P1_N3120), .IN1(n7109), .Q(P1_add_428_n188) );
  NAND2X0 P1_add_428_U199 ( .IN1(P1_N3120), .IN2(n7109), .QN(P1_add_428_n189)
         );
  NAND2X0 P1_add_428_U198 ( .IN1(P1_add_428_n188), .IN2(P1_add_428_n189), 
        .QN(P1_add_428_n187) );
  NOR2X0 P1_add_428_U197 ( .QN(P1_add_428_n185), .IN1(P1_add_428_n184), 
        .IN2(P1_add_428_n187) );
  AND2X1 P1_add_428_U196 ( .IN1(P1_add_428_n184), .IN2(P1_add_428_n187), 
        .Q(P1_add_428_n186) );
  NOR2X0 P1_add_428_U195 ( .QN(P1_N3362), .IN1(P1_add_428_n185), 
        .IN2(P1_add_428_n186) );
  NAND2X0 P1_add_428_U194 ( .IN1(P1_N5165), .IN2(P1_add_428_n184), 
        .QN(P1_add_428_n181) );
  OR2X1 P1_add_428_U193 ( .IN2(P1_N5165), .IN1(P1_add_428_n184), 
        .Q(P1_add_428_n183) );
  NAND2X0 P1_add_428_U192 ( .IN1(P1_N3120), .IN2(P1_add_428_n183), 
        .QN(P1_add_428_n182) );
  NAND2X0 P1_add_428_U191 ( .IN1(P1_add_428_n181), .IN2(P1_add_428_n182), 
        .QN(P1_add_428_n174) );
  OR2X1 P1_add_428_U189 ( .IN2(P1_N3121), .IN1(n7105), .Q(P1_add_428_n178) );
  NAND2X0 P1_add_428_U188 ( .IN1(P1_N3121), .IN2(n7105), .QN(P1_add_428_n179)
         );
  NAND2X0 P1_add_428_U187 ( .IN1(P1_add_428_n178), .IN2(P1_add_428_n179), 
        .QN(P1_add_428_n177) );
  NOR2X0 P1_add_428_U186 ( .QN(P1_add_428_n175), .IN1(P1_add_428_n174), 
        .IN2(P1_add_428_n177) );
  AND2X1 P1_add_428_U185 ( .IN1(P1_add_428_n174), .IN2(P1_add_428_n177), 
        .Q(P1_add_428_n176) );
  NOR2X0 P1_add_428_U184 ( .QN(P1_N3363), .IN1(P1_add_428_n175), 
        .IN2(P1_add_428_n176) );
  NAND2X0 P1_add_428_U183 ( .IN1(n7106), .IN2(P1_add_428_n174), 
        .QN(P1_add_428_n171) );
  OR2X1 P1_add_428_U182 ( .IN2(n7106), .IN1(P1_add_428_n174), 
        .Q(P1_add_428_n173) );
  OR2X1 P1_add_428_U308 ( .IN2(P1_N3104), .IN1(n4803), .Q(P1_add_428_n278) );
  NAND2X0 P1_add_428_U307 ( .IN1(P1_N3104), .IN2(n4803), .QN(P1_add_428_n279)
         );
  NAND2X0 P1_add_428_U306 ( .IN1(P1_add_428_n278), .IN2(P1_add_428_n279), 
        .QN(P1_N3346) );
  NAND2X0 P1_add_428_U304 ( .IN1(P1_N3104), .IN2(n7034), .QN(P1_add_428_n151)
         );
  OR2X1 P1_add_428_U303 ( .IN2(P1_add_428_n151), .IN1(n7051), 
        .Q(P1_add_428_n275) );
  NAND2X0 P1_add_428_U302 ( .IN1(n7051), .IN2(P1_add_428_n151), 
        .QN(P1_add_428_n277) );
  NAND2X0 P1_add_428_U301 ( .IN1(P1_N3105), .IN2(P1_add_428_n277), 
        .QN(P1_add_428_n276) );
  NAND2X0 P1_add_428_U300 ( .IN1(P1_add_428_n275), .IN2(P1_add_428_n276), 
        .QN(P1_add_428_n52) );
  NAND2X0 P1_add_428_U299 ( .IN1(P1_N5151), .IN2(P1_add_428_n52), 
        .QN(P1_add_428_n272) );
  OR2X1 P1_add_428_U298 ( .IN2(P1_N5151), .IN1(P1_add_428_n52), 
        .Q(P1_add_428_n274) );
  NAND2X0 P1_add_428_U297 ( .IN1(P1_N3106), .IN2(P1_add_428_n274), 
        .QN(P1_add_428_n273) );
  NAND2X0 P1_add_428_U296 ( .IN1(P1_add_428_n272), .IN2(P1_add_428_n273), 
        .QN(P1_add_428_n45) );
  NAND2X0 P1_add_428_U295 ( .IN1(P1_N5152), .IN2(P1_add_428_n45), 
        .QN(P1_add_428_n269) );
  OR2X1 P1_add_428_U294 ( .IN2(P1_N5152), .IN1(P1_add_428_n45), 
        .Q(P1_add_428_n271) );
  NAND2X0 P1_add_428_U293 ( .IN1(P1_N3107), .IN2(P1_add_428_n271), 
        .QN(P1_add_428_n270) );
  NAND2X0 P1_add_428_U292 ( .IN1(P1_add_428_n269), .IN2(P1_add_428_n270), 
        .QN(P1_add_428_n38) );
  NAND2X0 P1_add_428_U291 ( .IN1(n7036), .IN2(P1_add_428_n38), 
        .QN(P1_add_428_n266) );
  OR2X1 P1_add_428_U290 ( .IN2(n7036), .IN1(P1_add_428_n38), 
        .Q(P1_add_428_n268) );
  NAND2X0 P1_add_428_U289 ( .IN1(P1_N3108), .IN2(P1_add_428_n268), 
        .QN(P1_add_428_n267) );
  NAND2X0 P1_add_428_U288 ( .IN1(P1_add_428_n266), .IN2(P1_add_428_n267), 
        .QN(P1_add_428_n31) );
  NAND2X0 P1_add_428_U287 ( .IN1(n7081), .IN2(P1_add_428_n31), 
        .QN(P1_add_428_n263) );
  OR2X1 P1_add_428_U286 ( .IN2(n7081), .IN1(P1_add_428_n31), 
        .Q(P1_add_428_n265) );
  NAND2X0 P1_add_428_U285 ( .IN1(P1_N3109), .IN2(P1_add_428_n265), 
        .QN(P1_add_428_n264) );
  NAND2X0 P1_add_428_U284 ( .IN1(P1_add_428_n263), .IN2(P1_add_428_n264), 
        .QN(P1_add_428_n24) );
  NAND2X0 P1_add_428_U283 ( .IN1(P1_N5155), .IN2(P1_add_428_n24), 
        .QN(P1_add_428_n260) );
  OR2X1 P1_add_428_U282 ( .IN2(P1_N5155), .IN1(P1_add_428_n24), 
        .Q(P1_add_428_n262) );
  NAND2X0 P1_add_428_U281 ( .IN1(P1_N3110), .IN2(P1_add_428_n262), 
        .QN(P1_add_428_n261) );
  NAND2X0 P1_add_428_U280 ( .IN1(P1_add_428_n260), .IN2(P1_add_428_n261), 
        .QN(P1_add_428_n17) );
  NAND2X0 P1_add_428_U279 ( .IN1(n7075), .IN2(P1_add_428_n17), 
        .QN(P1_add_428_n257) );
  OR2X1 P1_add_428_U278 ( .IN2(n7075), .IN1(P1_add_428_n17), 
        .Q(P1_add_428_n259) );
  NAND2X0 P1_add_428_U277 ( .IN1(P1_N3111), .IN2(P1_add_428_n259), 
        .QN(P1_add_428_n258) );
  NAND2X0 P1_add_428_U276 ( .IN1(P1_add_428_n257), .IN2(P1_add_428_n258), 
        .QN(P1_add_428_n10) );
  NAND2X0 P1_add_428_U275 ( .IN1(n7072), .IN2(P1_add_428_n10), 
        .QN(P1_add_428_n254) );
  OR2X1 P1_sub_448_U26 ( .IN2(P1_sub_448_n32), .IN1(P1_sub_448_n31), 
        .Q(P1_sub_448_n30) );
  NAND2X0 P1_sub_448_U25 ( .IN1(P1_sub_448_n29), .IN2(P1_sub_448_n30), 
        .QN(P1_N3724) );
  NAND2X0 P1_sub_448_U24 ( .IN1(n7080), .IN2(P1_sub_448_n28), 
        .QN(P1_sub_448_n26) );
  OR2X1 P1_sub_448_U23 ( .IN2(n7080), .IN1(P1_sub_448_n28), .Q(P1_sub_448_n27)
         );
  NAND2X0 P1_sub_448_U22 ( .IN1(P1_sub_448_n26), .IN2(P1_sub_448_n27), 
        .QN(P1_sub_448_n24) );
  NAND2X0 P1_sub_448_U21 ( .IN1(P1_sub_448_n24), .IN2(P1_sub_448_n25), 
        .QN(P1_sub_448_n22) );
  OR2X1 P1_sub_448_U20 ( .IN2(P1_sub_448_n25), .IN1(P1_sub_448_n24), 
        .Q(P1_sub_448_n23) );
  NAND2X0 P1_sub_448_U19 ( .IN1(P1_sub_448_n22), .IN2(P1_sub_448_n23), 
        .QN(P1_N3725) );
  NAND2X0 P1_sub_448_U18 ( .IN1(n7075), .IN2(P1_sub_448_n21), 
        .QN(P1_sub_448_n19) );
  OR2X1 P1_sub_448_U17 ( .IN2(n7075), .IN1(P1_sub_448_n21), .Q(P1_sub_448_n20)
         );
  NAND2X0 P1_sub_448_U16 ( .IN1(P1_sub_448_n19), .IN2(P1_sub_448_n20), 
        .QN(P1_sub_448_n17) );
  NAND2X0 P1_sub_448_U15 ( .IN1(P1_sub_448_n17), .IN2(P1_sub_448_n18), 
        .QN(P1_sub_448_n15) );
  OR2X1 P1_sub_448_U14 ( .IN2(P1_sub_448_n18), .IN1(P1_sub_448_n17), 
        .Q(P1_sub_448_n16) );
  NAND2X0 P1_sub_448_U13 ( .IN1(P1_sub_448_n15), .IN2(P1_sub_448_n16), 
        .QN(P1_N3726) );
  NAND2X0 P1_sub_448_U12 ( .IN1(P1_N5157), .IN2(P1_sub_448_n14), 
        .QN(P1_sub_448_n12) );
  OR2X1 P1_sub_448_U11 ( .IN2(P1_N5157), .IN1(P1_sub_448_n14), 
        .Q(P1_sub_448_n13) );
  NAND2X0 P1_sub_448_U10 ( .IN1(P1_sub_448_n12), .IN2(P1_sub_448_n13), 
        .QN(P1_sub_448_n10) );
  NAND2X0 P1_sub_448_U9 ( .IN1(P1_sub_448_n10), .IN2(P1_sub_448_n11), 
        .QN(P1_sub_448_n8) );
  OR2X1 P1_sub_448_U8 ( .IN2(P1_sub_448_n11), .IN1(P1_sub_448_n10), 
        .Q(P1_sub_448_n9) );
  NAND2X0 P1_sub_448_U7 ( .IN1(P1_sub_448_n8), .IN2(P1_sub_448_n9), 
        .QN(P1_N3727) );
  NAND2X0 P1_sub_448_U6 ( .IN1(P1_N5158), .IN2(P1_sub_448_n7), 
        .QN(P1_sub_448_n5) );
  OR2X1 P1_sub_448_U5 ( .IN2(P1_N5158), .IN1(P1_sub_448_n7), .Q(P1_sub_448_n6)
         );
  NAND2X0 P1_sub_448_U4 ( .IN1(P1_sub_448_n5), .IN2(P1_sub_448_n6), 
        .QN(P1_sub_448_n3) );
  NAND2X0 P1_sub_448_U3 ( .IN1(P1_sub_448_n3), .IN2(P1_sub_448_n4), 
        .QN(P1_sub_448_n1) );
  OR2X1 P1_sub_448_U2 ( .IN2(P1_sub_448_n4), .IN1(P1_sub_448_n3), 
        .Q(P1_sub_448_n2) );
  NAND2X0 P1_sub_448_U1 ( .IN1(P1_sub_448_n1), .IN2(P1_sub_448_n2), 
        .QN(P1_N3728) );
  NAND2X0 P1_sub_448_U119 ( .IN1(P1_sub_448_n124), .IN2(P1_sub_448_n125), 
        .QN(P1_sub_448_n123) );
  NAND2X0 P1_sub_448_U118 ( .IN1(P1_sub_448_n122), .IN2(P1_sub_448_n123), 
        .QN(P1_sub_448_n116) );
  NAND2X0 P1_sub_448_U117 ( .IN1(P1_sub_448_n121), .IN2(P1_sub_448_n116), 
        .QN(P1_sub_448_n119) );
  OR2X1 P1_sub_448_U116 ( .IN2(P1_sub_448_n116), .IN1(P1_sub_448_n121), 
        .Q(P1_sub_448_n120) );
  NAND2X0 P1_sub_448_U115 ( .IN1(P1_sub_448_n119), .IN2(P1_sub_448_n120), 
        .QN(P1_N3741) );
  INVX0 P1_sub_448_U114 ( .ZN(P1_sub_448_n105), .INP(P1_N3500) );
  NAND2X0 P1_sub_448_U113 ( .IN1(P1_N5172), .IN2(P1_sub_448_n105), 
        .QN(P1_sub_448_n117) );
  OR2X1 P1_sub_448_U112 ( .IN2(P1_N5172), .IN1(P1_sub_448_n105), 
        .Q(P1_sub_448_n118) );
  NAND2X0 P1_sub_448_U111 ( .IN1(P1_sub_448_n117), .IN2(P1_sub_448_n118), 
        .QN(P1_sub_448_n111) );
  NAND2X0 P1_sub_448_U110 ( .IN1(n7089), .IN2(P1_sub_448_n116), 
        .QN(P1_sub_448_n112) );
  OR2X1 P1_sub_448_U109 ( .IN2(n7089), .IN1(P1_sub_448_n116), 
        .Q(P1_sub_448_n114) );
  NAND2X0 P1_sub_448_U108 ( .IN1(P1_sub_448_n114), .IN2(P1_sub_448_n115), 
        .QN(P1_sub_448_n113) );
  NAND2X0 P1_sub_448_U107 ( .IN1(P1_sub_448_n112), .IN2(P1_sub_448_n113), 
        .QN(P1_sub_448_n106) );
  NAND2X0 P1_sub_448_U106 ( .IN1(P1_sub_448_n111), .IN2(P1_sub_448_n106), 
        .QN(P1_sub_448_n109) );
  OR2X1 P1_sub_448_U105 ( .IN2(P1_sub_448_n106), .IN1(P1_sub_448_n111), 
        .Q(P1_sub_448_n110) );
  NAND2X0 P1_sub_448_U104 ( .IN1(P1_sub_448_n109), .IN2(P1_sub_448_n110), 
        .QN(P1_N3742) );
  INVX0 P1_sub_448_U103 ( .ZN(P1_sub_448_n95), .INP(P1_N3501) );
  NAND2X0 P1_sub_448_U102 ( .IN1(P1_N5173), .IN2(P1_sub_448_n95), 
        .QN(P1_sub_448_n107) );
  OR2X1 P1_sub_448_U101 ( .IN2(P1_N5173), .IN1(P1_sub_448_n95), 
        .Q(P1_sub_448_n108) );
  NAND2X0 P1_sub_448_U100 ( .IN1(P1_sub_448_n107), .IN2(P1_sub_448_n108), 
        .QN(P1_sub_448_n101) );
  NAND2X0 P1_sub_448_U99 ( .IN1(P1_N5172), .IN2(P1_sub_448_n106), 
        .QN(P1_sub_448_n102) );
  OR2X1 P1_sub_448_U98 ( .IN2(P1_N5172), .IN1(P1_sub_448_n106), 
        .Q(P1_sub_448_n104) );
  NAND2X0 P1_sub_448_U97 ( .IN1(P1_sub_448_n104), .IN2(P1_sub_448_n105), 
        .QN(P1_sub_448_n103) );
  NAND2X0 P1_sub_448_U96 ( .IN1(P1_sub_448_n102), .IN2(P1_sub_448_n103), 
        .QN(P1_sub_448_n96) );
  NAND2X0 P1_sub_448_U95 ( .IN1(P1_sub_448_n101), .IN2(P1_sub_448_n96), 
        .QN(P1_sub_448_n99) );
  OR2X1 P1_sub_448_U94 ( .IN2(P1_sub_448_n96), .IN1(P1_sub_448_n101), 
        .Q(P1_sub_448_n100) );
  NAND2X0 P1_sub_448_U93 ( .IN1(P1_sub_448_n99), .IN2(P1_sub_448_n100), 
        .QN(P1_N3743) );
  INVX0 P1_sub_448_U92 ( .ZN(P1_sub_448_n85), .INP(P1_N3502) );
  NAND2X0 P1_sub_448_U91 ( .IN1(n7129), .IN2(P1_sub_448_n85), 
        .QN(P1_sub_448_n97) );
  OR2X1 P1_sub_448_U90 ( .IN2(n7129), .IN1(P1_sub_448_n85), .Q(P1_sub_448_n98)
         );
  NAND2X0 P1_sub_448_U89 ( .IN1(P1_sub_448_n97), .IN2(P1_sub_448_n98), 
        .QN(P1_sub_448_n91) );
  NAND2X0 P1_sub_448_U88 ( .IN1(P1_N5173), .IN2(P1_sub_448_n96), 
        .QN(P1_sub_448_n92) );
  OR2X1 P1_sub_448_U87 ( .IN2(P1_N5173), .IN1(P1_sub_448_n96), 
        .Q(P1_sub_448_n94) );
  NAND2X0 P1_sub_448_U86 ( .IN1(P1_sub_448_n94), .IN2(P1_sub_448_n95), 
        .QN(P1_sub_448_n93) );
  NAND2X0 P1_sub_448_U85 ( .IN1(P1_sub_448_n92), .IN2(P1_sub_448_n93), 
        .QN(P1_sub_448_n86) );
  NAND2X0 P1_sub_448_U84 ( .IN1(P1_sub_448_n91), .IN2(P1_sub_448_n86), 
        .QN(P1_sub_448_n89) );
  OR2X1 P1_sub_448_U83 ( .IN2(P1_sub_448_n86), .IN1(P1_sub_448_n91), 
        .Q(P1_sub_448_n90) );
  NAND2X0 P1_sub_448_U82 ( .IN1(P1_sub_448_n89), .IN2(P1_sub_448_n90), 
        .QN(P1_N3744) );
  INVX0 P1_sub_448_U81 ( .ZN(P1_sub_448_n75), .INP(P1_N3503) );
  NAND2X0 P1_sub_448_U80 ( .IN1(P1_N5175), .IN2(P1_sub_448_n75), 
        .QN(P1_sub_448_n87) );
  OR2X1 P1_sub_448_U79 ( .IN2(P1_N5175), .IN1(P1_sub_448_n75), 
        .Q(P1_sub_448_n88) );
  NAND2X0 P1_sub_448_U78 ( .IN1(P1_sub_448_n87), .IN2(P1_sub_448_n88), 
        .QN(P1_sub_448_n81) );
  NAND2X0 P1_sub_448_U77 ( .IN1(n7129), .IN2(P1_sub_448_n86), 
        .QN(P1_sub_448_n82) );
  OR2X1 P1_sub_448_U76 ( .IN2(n7129), .IN1(P1_sub_448_n86), .Q(P1_sub_448_n84)
         );
  NAND2X0 P1_sub_448_U75 ( .IN1(P1_sub_448_n84), .IN2(P1_sub_448_n85), 
        .QN(P1_sub_448_n83) );
  NAND2X0 P1_sub_448_U74 ( .IN1(P1_sub_448_n82), .IN2(P1_sub_448_n83), 
        .QN(P1_sub_448_n76) );
  NAND2X0 P1_sub_448_U73 ( .IN1(P1_sub_448_n81), .IN2(P1_sub_448_n76), 
        .QN(P1_sub_448_n79) );
  OR2X1 P1_sub_448_U72 ( .IN2(P1_sub_448_n76), .IN1(P1_sub_448_n81), 
        .Q(P1_sub_448_n80) );
  NAND2X0 P1_sub_448_U71 ( .IN1(P1_sub_448_n79), .IN2(P1_sub_448_n80), 
        .QN(P1_N3745) );
  INVX0 P1_sub_448_U70 ( .ZN(P1_sub_448_n64), .INP(P1_N3504) );
  NAND2X0 P1_sub_448_U69 ( .IN1(n7122), .IN2(P1_sub_448_n64), 
        .QN(P1_sub_448_n77) );
  OR2X1 P1_sub_448_U68 ( .IN2(n7122), .IN1(P1_sub_448_n64), .Q(P1_sub_448_n78)
         );
  NAND2X0 P1_sub_448_U67 ( .IN1(P1_sub_448_n77), .IN2(P1_sub_448_n78), 
        .QN(P1_sub_448_n71) );
  NAND2X0 P1_sub_448_U66 ( .IN1(P1_N5175), .IN2(P1_sub_448_n76), 
        .QN(P1_sub_448_n72) );
  OR2X1 P1_sub_448_U65 ( .IN2(P1_N5175), .IN1(P1_sub_448_n76), 
        .Q(P1_sub_448_n74) );
  NAND2X0 P1_sub_448_U64 ( .IN1(P1_sub_448_n74), .IN2(P1_sub_448_n75), 
        .QN(P1_sub_448_n73) );
  NAND2X0 P1_sub_448_U63 ( .IN1(P1_sub_448_n72), .IN2(P1_sub_448_n73), 
        .QN(P1_sub_448_n65) );
  NAND2X0 P1_sub_448_U62 ( .IN1(P1_sub_448_n71), .IN2(P1_sub_448_n65), 
        .QN(P1_sub_448_n69) );
  OR2X1 P1_sub_448_U61 ( .IN2(P1_sub_448_n65), .IN1(P1_sub_448_n71), 
        .Q(P1_sub_448_n70) );
  NAND2X0 P1_sub_448_U60 ( .IN1(P1_sub_448_n69), .IN2(P1_sub_448_n70), 
        .QN(P1_N3746) );
  OR2X1 P1_sub_448_U58 ( .IN2(P1_N3505), .IN1(n7117), .Q(P1_sub_448_n66) );
  NAND2X0 P1_sub_448_U57 ( .IN1(P1_N3505), .IN2(n7117), .QN(P1_sub_448_n67) );
  NAND2X0 P1_sub_448_U56 ( .IN1(P1_sub_448_n66), .IN2(P1_sub_448_n67), 
        .QN(P1_sub_448_n60) );
  NAND2X0 P1_sub_448_U55 ( .IN1(n7122), .IN2(P1_sub_448_n65), 
        .QN(P1_sub_448_n61) );
  OR2X1 P1_sub_448_U54 ( .IN2(n7122), .IN1(P1_sub_448_n65), .Q(P1_sub_448_n63)
         );
  NAND2X0 P1_sub_448_U53 ( .IN1(P1_sub_448_n63), .IN2(P1_sub_448_n64), 
        .QN(P1_sub_448_n62) );
  NAND2X0 P1_sub_448_U52 ( .IN1(P1_sub_448_n61), .IN2(P1_sub_448_n62), 
        .QN(P1_sub_448_n59) );
  NAND2X0 P1_sub_448_U51 ( .IN1(P1_sub_448_n60), .IN2(P1_sub_448_n59), 
        .QN(P1_sub_448_n57) );
  OR2X1 P1_sub_448_U50 ( .IN2(P1_sub_448_n60), .IN1(P1_sub_448_n59), 
        .Q(P1_sub_448_n58) );
  NAND2X0 P1_sub_448_U49 ( .IN1(P1_sub_448_n57), .IN2(P1_sub_448_n58), 
        .QN(P1_N3747) );
  NAND2X0 P1_sub_448_U48 ( .IN1(n7046), .IN2(P1_sub_448_n56), 
        .QN(P1_sub_448_n54) );
  OR2X1 P1_sub_448_U47 ( .IN2(n7046), .IN1(P1_sub_448_n56), .Q(P1_sub_448_n55)
         );
  NAND2X0 P1_sub_448_U46 ( .IN1(P1_sub_448_n54), .IN2(P1_sub_448_n55), 
        .QN(P1_sub_448_n52) );
  NAND2X0 P1_sub_448_U45 ( .IN1(P1_sub_448_n52), .IN2(P1_sub_448_n53), 
        .QN(P1_sub_448_n50) );
  OR2X1 P1_sub_448_U44 ( .IN2(P1_sub_448_n53), .IN1(P1_sub_448_n52), 
        .Q(P1_sub_448_n51) );
  NAND2X0 P1_sub_448_U43 ( .IN1(P1_sub_448_n50), .IN2(P1_sub_448_n51), 
        .QN(P1_N3721) );
  NAND2X0 P1_sub_448_U42 ( .IN1(P1_N5152), .IN2(P1_sub_448_n49), 
        .QN(P1_sub_448_n47) );
  OR2X1 P1_sub_448_U41 ( .IN2(P1_N5152), .IN1(P1_sub_448_n49), 
        .Q(P1_sub_448_n48) );
  NAND2X0 P1_sub_448_U40 ( .IN1(P1_sub_448_n47), .IN2(P1_sub_448_n48), 
        .QN(P1_sub_448_n45) );
  NAND2X0 P1_sub_448_U39 ( .IN1(P1_sub_448_n45), .IN2(P1_sub_448_n46), 
        .QN(P1_sub_448_n43) );
  OR2X1 P1_sub_448_U38 ( .IN2(P1_sub_448_n46), .IN1(P1_sub_448_n45), 
        .Q(P1_sub_448_n44) );
  NAND2X0 P1_sub_448_U37 ( .IN1(P1_sub_448_n43), .IN2(P1_sub_448_n44), 
        .QN(P1_N3722) );
  NAND2X0 P1_sub_448_U36 ( .IN1(n7036), .IN2(P1_sub_448_n42), 
        .QN(P1_sub_448_n40) );
  OR2X1 P1_sub_448_U35 ( .IN2(n7036), .IN1(P1_sub_448_n42), .Q(P1_sub_448_n41)
         );
  NAND2X0 P1_sub_448_U34 ( .IN1(P1_sub_448_n40), .IN2(P1_sub_448_n41), 
        .QN(P1_sub_448_n38) );
  NAND2X0 P1_sub_448_U33 ( .IN1(P1_sub_448_n38), .IN2(P1_sub_448_n39), 
        .QN(P1_sub_448_n36) );
  OR2X1 P1_sub_448_U32 ( .IN2(P1_sub_448_n39), .IN1(P1_sub_448_n38), 
        .Q(P1_sub_448_n37) );
  NAND2X0 P1_sub_448_U31 ( .IN1(P1_sub_448_n36), .IN2(P1_sub_448_n37), 
        .QN(P1_N3723) );
  NAND2X0 P1_sub_448_U30 ( .IN1(n7081), .IN2(P1_sub_448_n35), 
        .QN(P1_sub_448_n33) );
  OR2X1 P1_sub_448_U29 ( .IN2(n7081), .IN1(P1_sub_448_n35), .Q(P1_sub_448_n34)
         );
  NAND2X0 P1_sub_448_U28 ( .IN1(P1_sub_448_n33), .IN2(P1_sub_448_n34), 
        .QN(P1_sub_448_n31) );
  NAND2X0 P1_sub_448_U27 ( .IN1(P1_sub_448_n31), .IN2(P1_sub_448_n32), 
        .QN(P1_sub_448_n29) );
  NAND2X0 P1_sub_448_U212 ( .IN1(P1_sub_448_n210), .IN2(P1_sub_448_n211), 
        .QN(P1_sub_448_n204) );
  NAND2X0 P1_sub_448_U211 ( .IN1(P1_sub_448_n209), .IN2(P1_sub_448_n204), 
        .QN(P1_sub_448_n207) );
  OR2X1 P1_sub_448_U210 ( .IN2(P1_sub_448_n204), .IN1(P1_sub_448_n209), 
        .Q(P1_sub_448_n208) );
  NAND2X0 P1_sub_448_U209 ( .IN1(P1_sub_448_n207), .IN2(P1_sub_448_n208), 
        .QN(P1_N3733) );
  INVX0 P1_sub_448_U208 ( .ZN(P1_sub_448_n193), .INP(P1_N3492) );
  NAND2X0 P1_sub_448_U207 ( .IN1(n7113), .IN2(P1_sub_448_n193), 
        .QN(P1_sub_448_n205) );
  OR2X1 P1_sub_448_U206 ( .IN2(n7113), .IN1(P1_sub_448_n193), 
        .Q(P1_sub_448_n206) );
  NAND2X0 P1_sub_448_U205 ( .IN1(P1_sub_448_n205), .IN2(P1_sub_448_n206), 
        .QN(P1_sub_448_n199) );
  NAND2X0 P1_sub_448_U204 ( .IN1(n7116), .IN2(P1_sub_448_n204), 
        .QN(P1_sub_448_n200) );
  OR2X1 P1_sub_448_U203 ( .IN2(n7116), .IN1(P1_sub_448_n204), 
        .Q(P1_sub_448_n202) );
  NAND2X0 P1_sub_448_U202 ( .IN1(P1_sub_448_n202), .IN2(P1_sub_448_n203), 
        .QN(P1_sub_448_n201) );
  NAND2X0 P1_sub_448_U201 ( .IN1(P1_sub_448_n200), .IN2(P1_sub_448_n201), 
        .QN(P1_sub_448_n194) );
  NAND2X0 P1_sub_448_U200 ( .IN1(P1_sub_448_n199), .IN2(P1_sub_448_n194), 
        .QN(P1_sub_448_n197) );
  OR2X1 P1_sub_448_U199 ( .IN2(P1_sub_448_n194), .IN1(P1_sub_448_n199), 
        .Q(P1_sub_448_n198) );
  NAND2X0 P1_sub_448_U198 ( .IN1(P1_sub_448_n197), .IN2(P1_sub_448_n198), 
        .QN(P1_N3734) );
  INVX0 P1_sub_448_U197 ( .ZN(P1_sub_448_n183), .INP(P1_N3493) );
  NAND2X0 P1_sub_448_U196 ( .IN1(n7110), .IN2(P1_sub_448_n183), 
        .QN(P1_sub_448_n195) );
  OR2X1 P1_sub_448_U195 ( .IN2(n7110), .IN1(P1_sub_448_n183), 
        .Q(P1_sub_448_n196) );
  NAND2X0 P1_sub_448_U194 ( .IN1(P1_sub_448_n195), .IN2(P1_sub_448_n196), 
        .QN(P1_sub_448_n189) );
  NAND2X0 P1_sub_448_U193 ( .IN1(n7113), .IN2(P1_sub_448_n194), 
        .QN(P1_sub_448_n190) );
  OR2X1 P1_sub_448_U192 ( .IN2(n7113), .IN1(P1_sub_448_n194), 
        .Q(P1_sub_448_n192) );
  NAND2X0 P1_sub_448_U191 ( .IN1(P1_sub_448_n192), .IN2(P1_sub_448_n193), 
        .QN(P1_sub_448_n191) );
  NAND2X0 P1_sub_448_U190 ( .IN1(P1_sub_448_n190), .IN2(P1_sub_448_n191), 
        .QN(P1_sub_448_n184) );
  NAND2X0 P1_sub_448_U189 ( .IN1(P1_sub_448_n189), .IN2(P1_sub_448_n184), 
        .QN(P1_sub_448_n187) );
  OR2X1 P1_sub_448_U188 ( .IN2(P1_sub_448_n184), .IN1(P1_sub_448_n189), 
        .Q(P1_sub_448_n188) );
  NAND2X0 P1_sub_448_U187 ( .IN1(P1_sub_448_n187), .IN2(P1_sub_448_n188), 
        .QN(P1_N3735) );
  INVX0 P1_sub_448_U186 ( .ZN(P1_sub_448_n173), .INP(P1_N3494) );
  NAND2X0 P1_sub_448_U185 ( .IN1(P1_N5166), .IN2(P1_sub_448_n173), 
        .QN(P1_sub_448_n185) );
  OR2X1 P1_sub_448_U184 ( .IN2(P1_N5166), .IN1(P1_sub_448_n173), 
        .Q(P1_sub_448_n186) );
  NAND2X0 P1_sub_448_U183 ( .IN1(P1_sub_448_n185), .IN2(P1_sub_448_n186), 
        .QN(P1_sub_448_n179) );
  NAND2X0 P1_sub_448_U182 ( .IN1(n7110), .IN2(P1_sub_448_n184), 
        .QN(P1_sub_448_n180) );
  OR2X1 P1_sub_448_U181 ( .IN2(n7110), .IN1(P1_sub_448_n184), 
        .Q(P1_sub_448_n182) );
  NAND2X0 P1_sub_448_U180 ( .IN1(P1_sub_448_n182), .IN2(P1_sub_448_n183), 
        .QN(P1_sub_448_n181) );
  NAND2X0 P1_sub_448_U179 ( .IN1(P1_sub_448_n180), .IN2(P1_sub_448_n181), 
        .QN(P1_sub_448_n174) );
  NAND2X0 P1_sub_448_U178 ( .IN1(P1_sub_448_n179), .IN2(P1_sub_448_n174), 
        .QN(P1_sub_448_n177) );
  OR2X1 P1_sub_448_U177 ( .IN2(P1_sub_448_n174), .IN1(P1_sub_448_n179), 
        .Q(P1_sub_448_n178) );
  NAND2X0 P1_sub_448_U176 ( .IN1(P1_sub_448_n177), .IN2(P1_sub_448_n178), 
        .QN(P1_N3736) );
  INVX0 P1_sub_448_U175 ( .ZN(P1_sub_448_n163), .INP(P1_N3495) );
  NAND2X0 P1_sub_448_U174 ( .IN1(n7103), .IN2(P1_sub_448_n163), 
        .QN(P1_sub_448_n175) );
  OR2X1 P1_sub_448_U173 ( .IN2(n7103), .IN1(P1_sub_448_n163), 
        .Q(P1_sub_448_n176) );
  NAND2X0 P1_sub_448_U172 ( .IN1(P1_sub_448_n175), .IN2(P1_sub_448_n176), 
        .QN(P1_sub_448_n169) );
  NAND2X0 P1_sub_448_U171 ( .IN1(P1_N5166), .IN2(P1_sub_448_n174), 
        .QN(P1_sub_448_n170) );
  OR2X1 P1_sub_448_U170 ( .IN2(P1_N5166), .IN1(P1_sub_448_n174), 
        .Q(P1_sub_448_n172) );
  NAND2X0 P1_sub_448_U169 ( .IN1(P1_sub_448_n172), .IN2(P1_sub_448_n173), 
        .QN(P1_sub_448_n171) );
  NAND2X0 P1_sub_448_U168 ( .IN1(P1_sub_448_n170), .IN2(P1_sub_448_n171), 
        .QN(P1_sub_448_n164) );
  NAND2X0 P1_sub_448_U167 ( .IN1(P1_sub_448_n169), .IN2(P1_sub_448_n164), 
        .QN(P1_sub_448_n167) );
  OR2X1 P1_sub_448_U166 ( .IN2(P1_sub_448_n164), .IN1(P1_sub_448_n169), 
        .Q(P1_sub_448_n168) );
  NAND2X0 P1_sub_448_U165 ( .IN1(P1_sub_448_n167), .IN2(P1_sub_448_n168), 
        .QN(P1_N3737) );
  INVX0 P1_sub_448_U164 ( .ZN(P1_sub_448_n145), .INP(P1_N3496) );
  NAND2X0 P1_sub_448_U163 ( .IN1(P1_N5168), .IN2(P1_sub_448_n145), 
        .QN(P1_sub_448_n165) );
  OR2X1 P1_sub_448_U162 ( .IN2(P1_N5168), .IN1(P1_sub_448_n145), 
        .Q(P1_sub_448_n166) );
  NAND2X0 P1_sub_448_U161 ( .IN1(P1_sub_448_n165), .IN2(P1_sub_448_n166), 
        .QN(P1_sub_448_n159) );
  NAND2X0 P1_sub_448_U160 ( .IN1(n7103), .IN2(P1_sub_448_n164), 
        .QN(P1_sub_448_n160) );
  OR2X1 P1_sub_448_U159 ( .IN2(n7103), .IN1(P1_sub_448_n164), 
        .Q(P1_sub_448_n162) );
  NAND2X0 P1_sub_448_U158 ( .IN1(P1_sub_448_n162), .IN2(P1_sub_448_n163), 
        .QN(P1_sub_448_n161) );
  NAND2X0 P1_sub_448_U157 ( .IN1(P1_sub_448_n160), .IN2(P1_sub_448_n161), 
        .QN(P1_sub_448_n146) );
  NAND2X0 P1_sub_448_U156 ( .IN1(P1_sub_448_n159), .IN2(P1_sub_448_n146), 
        .QN(P1_sub_448_n157) );
  OR2X1 P1_sub_448_U155 ( .IN2(P1_sub_448_n146), .IN1(P1_sub_448_n159), 
        .Q(P1_sub_448_n158) );
  NAND2X0 P1_sub_448_U154 ( .IN1(P1_sub_448_n157), .IN2(P1_sub_448_n158), 
        .QN(P1_N3738) );
  NAND2X0 P1_sub_448_U153 ( .IN1(P1_N5150), .IN2(P1_sub_448_n156), 
        .QN(P1_sub_448_n153) );
  NAND2X0 P1_sub_448_U152 ( .IN1(P1_N3478), .IN2(n7048), .QN(P1_sub_448_n154)
         );
  NAND2X0 P1_sub_448_U151 ( .IN1(P1_sub_448_n153), .IN2(P1_sub_448_n154), 
        .QN(P1_sub_448_n151) );
  NAND2X0 P1_sub_448_U150 ( .IN1(P1_sub_448_n151), .IN2(P1_sub_448_n152), 
        .QN(P1_sub_448_n149) );
  OR2X1 P1_sub_448_U149 ( .IN2(P1_sub_448_n152), .IN1(P1_sub_448_n151), 
        .Q(P1_sub_448_n150) );
  NAND2X0 P1_sub_448_U148 ( .IN1(P1_sub_448_n149), .IN2(P1_sub_448_n150), 
        .QN(P1_N3720) );
  INVX0 P1_sub_448_U147 ( .ZN(P1_sub_448_n135), .INP(P1_N3497) );
  NAND2X0 P1_sub_448_U146 ( .IN1(n7096), .IN2(P1_sub_448_n135), 
        .QN(P1_sub_448_n147) );
  OR2X1 P1_sub_448_U145 ( .IN2(n7096), .IN1(P1_sub_448_n135), 
        .Q(P1_sub_448_n148) );
  NAND2X0 P1_sub_448_U144 ( .IN1(P1_sub_448_n147), .IN2(P1_sub_448_n148), 
        .QN(P1_sub_448_n141) );
  NAND2X0 P1_sub_448_U143 ( .IN1(P1_N5168), .IN2(P1_sub_448_n146), 
        .QN(P1_sub_448_n142) );
  OR2X1 P1_sub_448_U142 ( .IN2(P1_N5168), .IN1(P1_sub_448_n146), 
        .Q(P1_sub_448_n144) );
  NAND2X0 P1_sub_448_U141 ( .IN1(P1_sub_448_n144), .IN2(P1_sub_448_n145), 
        .QN(P1_sub_448_n143) );
  NAND2X0 P1_sub_448_U140 ( .IN1(P1_sub_448_n142), .IN2(P1_sub_448_n143), 
        .QN(P1_sub_448_n136) );
  NAND2X0 P1_sub_448_U139 ( .IN1(P1_sub_448_n141), .IN2(P1_sub_448_n136), 
        .QN(P1_sub_448_n139) );
  OR2X1 P1_sub_448_U138 ( .IN2(P1_sub_448_n136), .IN1(P1_sub_448_n141), 
        .Q(P1_sub_448_n140) );
  NAND2X0 P1_sub_448_U137 ( .IN1(P1_sub_448_n139), .IN2(P1_sub_448_n140), 
        .QN(P1_N3739) );
  INVX0 P1_sub_448_U136 ( .ZN(P1_sub_448_n125), .INP(P1_N3498) );
  NAND2X0 P1_sub_448_U135 ( .IN1(n7093), .IN2(P1_sub_448_n125), 
        .QN(P1_sub_448_n137) );
  OR2X1 P1_sub_448_U134 ( .IN2(n7093), .IN1(P1_sub_448_n125), 
        .Q(P1_sub_448_n138) );
  NAND2X0 P1_sub_448_U133 ( .IN1(P1_sub_448_n137), .IN2(P1_sub_448_n138), 
        .QN(P1_sub_448_n131) );
  NAND2X0 P1_sub_448_U132 ( .IN1(n7096), .IN2(P1_sub_448_n136), 
        .QN(P1_sub_448_n132) );
  OR2X1 P1_sub_448_U131 ( .IN2(n7096), .IN1(P1_sub_448_n136), 
        .Q(P1_sub_448_n134) );
  NAND2X0 P1_sub_448_U130 ( .IN1(P1_sub_448_n134), .IN2(P1_sub_448_n135), 
        .QN(P1_sub_448_n133) );
  NAND2X0 P1_sub_448_U129 ( .IN1(P1_sub_448_n132), .IN2(P1_sub_448_n133), 
        .QN(P1_sub_448_n126) );
  NAND2X0 P1_sub_448_U128 ( .IN1(P1_sub_448_n131), .IN2(P1_sub_448_n126), 
        .QN(P1_sub_448_n129) );
  OR2X1 P1_sub_448_U127 ( .IN2(P1_sub_448_n126), .IN1(P1_sub_448_n131), 
        .Q(P1_sub_448_n130) );
  NAND2X0 P1_sub_448_U126 ( .IN1(P1_sub_448_n129), .IN2(P1_sub_448_n130), 
        .QN(P1_N3740) );
  INVX0 P1_sub_448_U125 ( .ZN(P1_sub_448_n115), .INP(P1_N3499) );
  NAND2X0 P1_sub_448_U124 ( .IN1(n7089), .IN2(P1_sub_448_n115), 
        .QN(P1_sub_448_n127) );
  OR2X1 P1_sub_448_U123 ( .IN2(n7089), .IN1(P1_sub_448_n115), 
        .Q(P1_sub_448_n128) );
  NAND2X0 P1_sub_448_U122 ( .IN1(P1_sub_448_n127), .IN2(P1_sub_448_n128), 
        .QN(P1_sub_448_n121) );
  NAND2X0 P1_sub_448_U121 ( .IN1(n7093), .IN2(P1_sub_448_n126), 
        .QN(P1_sub_448_n122) );
  OR2X1 P1_sub_448_U120 ( .IN2(n7093), .IN1(P1_sub_448_n126), 
        .Q(P1_sub_448_n124) );
  INVX0 P1_sub_448_U305 ( .ZN(P1_sub_448_n243), .INP(P1_N3487) );
  NAND2X0 P1_sub_448_U304 ( .IN1(P1_N5159), .IN2(P1_sub_448_n243), 
        .QN(P1_sub_448_n278) );
  OR2X1 P1_sub_448_U303 ( .IN2(P1_N5159), .IN1(P1_sub_448_n243), 
        .Q(P1_sub_448_n279) );
  NAND2X0 P1_sub_448_U302 ( .IN1(P1_sub_448_n278), .IN2(P1_sub_448_n279), 
        .QN(P1_sub_448_n249) );
  NAND2X0 P1_sub_448_U301 ( .IN1(P1_N5150), .IN2(P1_sub_448_n152), 
        .QN(P1_sub_448_n274) );
  NAND2X0 P1_sub_448_U299 ( .IN1(P1_sub_448_n277), .IN2(n7048), 
        .QN(P1_sub_448_n276) );
  INVX0 P1_sub_448_U298 ( .ZN(P1_sub_448_n156), .INP(P1_N3478) );
  NAND2X0 P1_sub_448_U297 ( .IN1(P1_sub_448_n276), .IN2(P1_sub_448_n156), 
        .QN(P1_sub_448_n275) );
  NAND2X0 P1_sub_448_U296 ( .IN1(P1_sub_448_n274), .IN2(P1_sub_448_n275), 
        .QN(P1_sub_448_n53) );
  NAND2X0 P1_sub_448_U295 ( .IN1(n7046), .IN2(P1_sub_448_n53), 
        .QN(P1_sub_448_n271) );
  OR2X1 P1_sub_448_U294 ( .IN2(n7046), .IN1(P1_sub_448_n53), 
        .Q(P1_sub_448_n273) );
  INVX0 P1_sub_448_U293 ( .ZN(P1_sub_448_n56), .INP(P1_N3479) );
  NAND2X0 P1_sub_448_U292 ( .IN1(P1_sub_448_n273), .IN2(P1_sub_448_n56), 
        .QN(P1_sub_448_n272) );
  NAND2X0 P1_sub_448_U291 ( .IN1(P1_sub_448_n271), .IN2(P1_sub_448_n272), 
        .QN(P1_sub_448_n46) );
  NAND2X0 P1_sub_448_U290 ( .IN1(P1_N5152), .IN2(P1_sub_448_n46), 
        .QN(P1_sub_448_n268) );
  OR2X1 P1_sub_448_U289 ( .IN2(P1_N5152), .IN1(P1_sub_448_n46), 
        .Q(P1_sub_448_n270) );
  INVX0 P1_sub_448_U288 ( .ZN(P1_sub_448_n49), .INP(P1_N3480) );
  NAND2X0 P1_sub_448_U287 ( .IN1(P1_sub_448_n270), .IN2(P1_sub_448_n49), 
        .QN(P1_sub_448_n269) );
  NAND2X0 P1_sub_448_U286 ( .IN1(P1_sub_448_n268), .IN2(P1_sub_448_n269), 
        .QN(P1_sub_448_n39) );
  NAND2X0 P1_sub_448_U285 ( .IN1(n7036), .IN2(P1_sub_448_n39), 
        .QN(P1_sub_448_n265) );
  OR2X1 P1_sub_448_U284 ( .IN2(n7036), .IN1(P1_sub_448_n39), 
        .Q(P1_sub_448_n267) );
  INVX0 P1_sub_448_U283 ( .ZN(P1_sub_448_n42), .INP(P1_N3481) );
  NAND2X0 P1_sub_448_U282 ( .IN1(P1_sub_448_n267), .IN2(P1_sub_448_n42), 
        .QN(P1_sub_448_n266) );
  NAND2X0 P1_sub_448_U281 ( .IN1(P1_sub_448_n265), .IN2(P1_sub_448_n266), 
        .QN(P1_sub_448_n32) );
  NAND2X0 P1_sub_448_U280 ( .IN1(n7081), .IN2(P1_sub_448_n32), 
        .QN(P1_sub_448_n262) );
  OR2X1 P1_sub_448_U279 ( .IN2(n7081), .IN1(P1_sub_448_n32), 
        .Q(P1_sub_448_n264) );
  INVX0 P1_sub_448_U278 ( .ZN(P1_sub_448_n35), .INP(P1_N3482) );
  NAND2X0 P1_sub_448_U277 ( .IN1(P1_sub_448_n264), .IN2(P1_sub_448_n35), 
        .QN(P1_sub_448_n263) );
  NAND2X0 P1_sub_448_U276 ( .IN1(P1_sub_448_n262), .IN2(P1_sub_448_n263), 
        .QN(P1_sub_448_n25) );
  NAND2X0 P1_sub_448_U275 ( .IN1(n7080), .IN2(P1_sub_448_n25), 
        .QN(P1_sub_448_n259) );
  OR2X1 P1_sub_448_U274 ( .IN2(n7080), .IN1(P1_sub_448_n25), 
        .Q(P1_sub_448_n261) );
  INVX0 P1_sub_448_U273 ( .ZN(P1_sub_448_n28), .INP(P1_N3483) );
  NAND2X0 P1_sub_448_U272 ( .IN1(P1_sub_448_n261), .IN2(P1_sub_448_n28), 
        .QN(P1_sub_448_n260) );
  NAND2X0 P1_sub_448_U271 ( .IN1(P1_sub_448_n259), .IN2(P1_sub_448_n260), 
        .QN(P1_sub_448_n18) );
  NAND2X0 P1_sub_448_U270 ( .IN1(n7075), .IN2(P1_sub_448_n18), 
        .QN(P1_sub_448_n256) );
  OR2X1 P1_sub_448_U269 ( .IN2(n7075), .IN1(P1_sub_448_n18), 
        .Q(P1_sub_448_n258) );
  INVX0 P1_sub_448_U268 ( .ZN(P1_sub_448_n21), .INP(P1_N3484) );
  NAND2X0 P1_sub_448_U267 ( .IN1(P1_sub_448_n258), .IN2(P1_sub_448_n21), 
        .QN(P1_sub_448_n257) );
  NAND2X0 P1_sub_448_U266 ( .IN1(P1_sub_448_n256), .IN2(P1_sub_448_n257), 
        .QN(P1_sub_448_n11) );
  NAND2X0 P1_sub_448_U265 ( .IN1(P1_N5157), .IN2(P1_sub_448_n11), 
        .QN(P1_sub_448_n253) );
  OR2X1 P1_sub_448_U264 ( .IN2(P1_N5157), .IN1(P1_sub_448_n11), 
        .Q(P1_sub_448_n255) );
  INVX0 P1_sub_448_U263 ( .ZN(P1_sub_448_n14), .INP(P1_N3485) );
  NAND2X0 P1_sub_448_U262 ( .IN1(P1_sub_448_n255), .IN2(P1_sub_448_n14), 
        .QN(P1_sub_448_n254) );
  NAND2X0 P1_sub_448_U261 ( .IN1(P1_sub_448_n253), .IN2(P1_sub_448_n254), 
        .QN(P1_sub_448_n4) );
  NAND2X0 P1_sub_448_U260 ( .IN1(P1_N5158), .IN2(P1_sub_448_n4), 
        .QN(P1_sub_448_n250) );
  OR2X1 P1_sub_448_U259 ( .IN2(P1_N5158), .IN1(P1_sub_448_n4), 
        .Q(P1_sub_448_n252) );
  INVX0 P1_sub_448_U258 ( .ZN(P1_sub_448_n7), .INP(P1_N3486) );
  NAND2X0 P1_sub_448_U257 ( .IN1(P1_sub_448_n252), .IN2(P1_sub_448_n7), 
        .QN(P1_sub_448_n251) );
  NAND2X0 P1_sub_448_U256 ( .IN1(P1_sub_448_n250), .IN2(P1_sub_448_n251), 
        .QN(P1_sub_448_n244) );
  NAND2X0 P1_sub_448_U255 ( .IN1(P1_sub_448_n249), .IN2(P1_sub_448_n244), 
        .QN(P1_sub_448_n247) );
  OR2X1 P1_sub_448_U254 ( .IN2(P1_sub_448_n244), .IN1(P1_sub_448_n249), 
        .Q(P1_sub_448_n248) );
  NAND2X0 P1_sub_448_U253 ( .IN1(P1_sub_448_n247), .IN2(P1_sub_448_n248), 
        .QN(P1_N3729) );
  INVX0 P1_sub_448_U252 ( .ZN(P1_sub_448_n233), .INP(P1_N3488) );
  NAND2X0 P1_sub_448_U251 ( .IN1(n7062), .IN2(P1_sub_448_n233), 
        .QN(P1_sub_448_n245) );
  OR2X1 P1_sub_448_U250 ( .IN2(n7062), .IN1(P1_sub_448_n233), 
        .Q(P1_sub_448_n246) );
  NAND2X0 P1_sub_448_U249 ( .IN1(P1_sub_448_n245), .IN2(P1_sub_448_n246), 
        .QN(P1_sub_448_n239) );
  NAND2X0 P1_sub_448_U248 ( .IN1(n7066), .IN2(P1_sub_448_n244), 
        .QN(P1_sub_448_n240) );
  OR2X1 P1_sub_448_U247 ( .IN2(P1_N5159), .IN1(P1_sub_448_n244), 
        .Q(P1_sub_448_n242) );
  NAND2X0 P1_sub_448_U246 ( .IN1(P1_sub_448_n242), .IN2(P1_sub_448_n243), 
        .QN(P1_sub_448_n241) );
  NAND2X0 P1_sub_448_U245 ( .IN1(P1_sub_448_n240), .IN2(P1_sub_448_n241), 
        .QN(P1_sub_448_n234) );
  NAND2X0 P1_sub_448_U244 ( .IN1(P1_sub_448_n239), .IN2(P1_sub_448_n234), 
        .QN(P1_sub_448_n237) );
  OR2X1 P1_sub_448_U243 ( .IN2(P1_sub_448_n234), .IN1(P1_sub_448_n239), 
        .Q(P1_sub_448_n238) );
  NAND2X0 P1_sub_448_U242 ( .IN1(P1_sub_448_n237), .IN2(P1_sub_448_n238), 
        .QN(P1_N3730) );
  INVX0 P1_sub_448_U241 ( .ZN(P1_sub_448_n223), .INP(P1_N3489) );
  NAND2X0 P1_sub_448_U240 ( .IN1(n7059), .IN2(P1_sub_448_n223), 
        .QN(P1_sub_448_n235) );
  OR2X1 P1_sub_448_U239 ( .IN2(n7059), .IN1(P1_sub_448_n223), 
        .Q(P1_sub_448_n236) );
  NAND2X0 P1_sub_448_U238 ( .IN1(P1_sub_448_n235), .IN2(P1_sub_448_n236), 
        .QN(P1_sub_448_n229) );
  NAND2X0 P1_sub_448_U237 ( .IN1(n7062), .IN2(P1_sub_448_n234), 
        .QN(P1_sub_448_n230) );
  OR2X1 P1_sub_448_U236 ( .IN2(n7062), .IN1(P1_sub_448_n234), 
        .Q(P1_sub_448_n232) );
  NAND2X0 P1_sub_448_U235 ( .IN1(P1_sub_448_n232), .IN2(P1_sub_448_n233), 
        .QN(P1_sub_448_n231) );
  NAND2X0 P1_sub_448_U234 ( .IN1(P1_sub_448_n230), .IN2(P1_sub_448_n231), 
        .QN(P1_sub_448_n224) );
  NAND2X0 P1_sub_448_U233 ( .IN1(P1_sub_448_n229), .IN2(P1_sub_448_n224), 
        .QN(P1_sub_448_n227) );
  OR2X1 P1_sub_448_U232 ( .IN2(P1_sub_448_n224), .IN1(P1_sub_448_n229), 
        .Q(P1_sub_448_n228) );
  NAND2X0 P1_sub_448_U231 ( .IN1(P1_sub_448_n227), .IN2(P1_sub_448_n228), 
        .QN(P1_N3731) );
  INVX0 P1_sub_448_U230 ( .ZN(P1_sub_448_n213), .INP(P1_N3490) );
  NAND2X0 P1_sub_448_U229 ( .IN1(n7055), .IN2(P1_sub_448_n213), 
        .QN(P1_sub_448_n225) );
  OR2X1 P1_sub_448_U228 ( .IN2(n7055), .IN1(P1_sub_448_n213), 
        .Q(P1_sub_448_n226) );
  NAND2X0 P1_sub_448_U227 ( .IN1(P1_sub_448_n225), .IN2(P1_sub_448_n226), 
        .QN(P1_sub_448_n219) );
  NAND2X0 P1_sub_448_U226 ( .IN1(n7059), .IN2(P1_sub_448_n224), 
        .QN(P1_sub_448_n220) );
  OR2X1 P1_sub_448_U225 ( .IN2(n7059), .IN1(P1_sub_448_n224), 
        .Q(P1_sub_448_n222) );
  NAND2X0 P1_sub_448_U224 ( .IN1(P1_sub_448_n222), .IN2(P1_sub_448_n223), 
        .QN(P1_sub_448_n221) );
  NAND2X0 P1_sub_448_U223 ( .IN1(P1_sub_448_n220), .IN2(P1_sub_448_n221), 
        .QN(P1_sub_448_n214) );
  NAND2X0 P1_sub_448_U222 ( .IN1(P1_sub_448_n219), .IN2(P1_sub_448_n214), 
        .QN(P1_sub_448_n217) );
  OR2X1 P1_sub_448_U221 ( .IN2(P1_sub_448_n214), .IN1(P1_sub_448_n219), 
        .Q(P1_sub_448_n218) );
  NAND2X0 P1_sub_448_U220 ( .IN1(P1_sub_448_n217), .IN2(P1_sub_448_n218), 
        .QN(P1_N3732) );
  INVX0 P1_sub_448_U219 ( .ZN(P1_sub_448_n203), .INP(P1_N3491) );
  NAND2X0 P1_sub_448_U218 ( .IN1(n7116), .IN2(P1_sub_448_n203), 
        .QN(P1_sub_448_n215) );
  OR2X1 P1_sub_448_U217 ( .IN2(n7116), .IN1(P1_sub_448_n203), 
        .Q(P1_sub_448_n216) );
  NAND2X0 P1_sub_448_U216 ( .IN1(P1_sub_448_n215), .IN2(P1_sub_448_n216), 
        .QN(P1_sub_448_n209) );
  NAND2X0 P1_sub_448_U215 ( .IN1(n7055), .IN2(P1_sub_448_n214), 
        .QN(P1_sub_448_n210) );
  OR2X1 P1_sub_448_U214 ( .IN2(n7055), .IN1(P1_sub_448_n214), 
        .Q(P1_sub_448_n212) );
  NAND2X0 P1_sub_448_U213 ( .IN1(P1_sub_448_n212), .IN2(P1_sub_448_n213), 
        .QN(P1_sub_448_n211) );
  INVX0 P1_sub_448_U310 ( .ZN(P1_sub_448_n281), .INP(P1_N3477) );
  NOR2X0 P1_sub_448_U309 ( .QN(P1_sub_448_n277), .IN1(P1_sub_448_n281), 
        .IN2(n7034) );
  INVX0 P1_sub_448_U308 ( .ZN(P1_sub_448_n152), .INP(P1_sub_448_n277) );
  NAND2X0 P1_sub_448_U307 ( .IN1(n7034), .IN2(P1_sub_448_n281), 
        .QN(P1_sub_448_n280) );
  NAND2X0 P1_sub_448_U306 ( .IN1(P1_sub_448_n152), .IN2(P1_sub_448_n280), 
        .QN(P1_N3719) );
  OR2X1 P1_add_468_U55 ( .IN2(P1_N3852), .IN1(n7045), .Q(P1_add_468_n54) );
  NAND2X0 P1_add_468_U54 ( .IN1(P1_N3852), .IN2(n7045), .QN(P1_add_468_n55) );
  NAND2X0 P1_add_468_U53 ( .IN1(P1_add_468_n54), .IN2(P1_add_468_n55), 
        .QN(P1_add_468_n53) );
  NOR2X0 P1_add_468_U52 ( .QN(P1_add_468_n50), .IN1(P1_add_468_n52), 
        .IN2(P1_add_468_n53) );
  AND2X1 P1_add_468_U51 ( .IN1(P1_add_468_n52), .IN2(P1_add_468_n53), 
        .Q(P1_add_468_n51) );
  NOR2X0 P1_add_468_U50 ( .QN(P1_N4094), .IN1(P1_add_468_n50), 
        .IN2(P1_add_468_n51) );
  OR2X1 P1_add_468_U48 ( .IN2(P1_N3853), .IN1(n7043), .Q(P1_add_468_n47) );
  NAND2X0 P1_add_468_U47 ( .IN1(P1_N3853), .IN2(n7043), .QN(P1_add_468_n48) );
  NAND2X0 P1_add_468_U46 ( .IN1(P1_add_468_n47), .IN2(P1_add_468_n48), 
        .QN(P1_add_468_n46) );
  NOR2X0 P1_add_468_U45 ( .QN(P1_add_468_n43), .IN1(P1_add_468_n45), 
        .IN2(P1_add_468_n46) );
  AND2X1 P1_add_468_U44 ( .IN1(P1_add_468_n45), .IN2(P1_add_468_n46), 
        .Q(P1_add_468_n44) );
  NOR2X0 P1_add_468_U43 ( .QN(P1_N4095), .IN1(P1_add_468_n43), 
        .IN2(P1_add_468_n44) );
  OR2X1 P1_add_468_U41 ( .IN2(P1_N3854), .IN1(n7037), .Q(P1_add_468_n40) );
  NAND2X0 P1_add_468_U40 ( .IN1(P1_N3854), .IN2(n7037), .QN(P1_add_468_n41) );
  NAND2X0 P1_add_468_U39 ( .IN1(P1_add_468_n40), .IN2(P1_add_468_n41), 
        .QN(P1_add_468_n39) );
  NOR2X0 P1_add_468_U38 ( .QN(P1_add_468_n36), .IN1(P1_add_468_n38), 
        .IN2(P1_add_468_n39) );
  AND2X1 P1_add_468_U37 ( .IN1(P1_add_468_n38), .IN2(P1_add_468_n39), 
        .Q(P1_add_468_n37) );
  NOR2X0 P1_add_468_U36 ( .QN(P1_N4096), .IN1(P1_add_468_n36), 
        .IN2(P1_add_468_n37) );
  OR2X1 P1_add_468_U34 ( .IN2(P1_N3855), .IN1(n7082), .Q(P1_add_468_n33) );
  NAND2X0 P1_add_468_U33 ( .IN1(P1_N3855), .IN2(n7082), .QN(P1_add_468_n34) );
  NAND2X0 P1_add_468_U32 ( .IN1(P1_add_468_n33), .IN2(P1_add_468_n34), 
        .QN(P1_add_468_n32) );
  NOR2X0 P1_add_468_U31 ( .QN(P1_add_468_n29), .IN1(P1_add_468_n31), 
        .IN2(P1_add_468_n32) );
  AND2X1 P1_add_468_U30 ( .IN1(P1_add_468_n31), .IN2(P1_add_468_n32), 
        .Q(P1_add_468_n30) );
  NOR2X0 P1_add_468_U29 ( .QN(P1_N4097), .IN1(P1_add_468_n29), 
        .IN2(P1_add_468_n30) );
  OR2X1 P1_add_468_U27 ( .IN2(P1_N3856), .IN1(n7079), .Q(P1_add_468_n26) );
  NAND2X0 P1_add_468_U26 ( .IN1(P1_N3856), .IN2(n7079), .QN(P1_add_468_n27) );
  NAND2X0 P1_add_468_U25 ( .IN1(P1_add_468_n26), .IN2(P1_add_468_n27), 
        .QN(P1_add_468_n25) );
  NOR2X0 P1_add_468_U24 ( .QN(P1_add_468_n22), .IN1(P1_add_468_n24), 
        .IN2(P1_add_468_n25) );
  AND2X1 P1_add_468_U23 ( .IN1(P1_add_468_n24), .IN2(P1_add_468_n25), 
        .Q(P1_add_468_n23) );
  NOR2X0 P1_add_468_U22 ( .QN(P1_N4098), .IN1(P1_add_468_n22), 
        .IN2(P1_add_468_n23) );
  OR2X1 P1_add_468_U20 ( .IN2(P1_N3857), .IN1(n7076), .Q(P1_add_468_n19) );
  NAND2X0 P1_add_468_U19 ( .IN1(P1_N3857), .IN2(n7076), .QN(P1_add_468_n20) );
  NAND2X0 P1_add_468_U18 ( .IN1(P1_add_468_n19), .IN2(P1_add_468_n20), 
        .QN(P1_add_468_n18) );
  NOR2X0 P1_add_468_U17 ( .QN(P1_add_468_n15), .IN1(P1_add_468_n17), 
        .IN2(P1_add_468_n18) );
  AND2X1 P1_add_468_U16 ( .IN1(P1_add_468_n17), .IN2(P1_add_468_n18), 
        .Q(P1_add_468_n16) );
  NOR2X0 P1_add_468_U15 ( .QN(P1_N4099), .IN1(P1_add_468_n15), 
        .IN2(P1_add_468_n16) );
  OR2X1 P1_add_468_U13 ( .IN2(P1_N3858), .IN1(n7073), .Q(P1_add_468_n12) );
  NAND2X0 P1_add_468_U12 ( .IN1(P1_N3858), .IN2(n7073), .QN(P1_add_468_n13) );
  NAND2X0 P1_add_468_U11 ( .IN1(P1_add_468_n12), .IN2(P1_add_468_n13), 
        .QN(P1_add_468_n11) );
  NOR2X0 P1_add_468_U10 ( .QN(P1_add_468_n8), .IN1(P1_add_468_n10), 
        .IN2(P1_add_468_n11) );
  AND2X1 P1_add_468_U9 ( .IN1(P1_add_468_n10), .IN2(P1_add_468_n11), 
        .Q(P1_add_468_n9) );
  NOR2X0 P1_add_468_U8 ( .QN(P1_N4100), .IN1(P1_add_468_n8), 
        .IN2(P1_add_468_n9) );
  OR2X1 P1_add_468_U6 ( .IN2(P1_N3859), .IN1(n7071), .Q(P1_add_468_n5) );
  NAND2X0 P1_add_468_U5 ( .IN1(P1_N3859), .IN2(n7071), .QN(P1_add_468_n6) );
  NAND2X0 P1_add_468_U4 ( .IN1(P1_add_468_n5), .IN2(P1_add_468_n6), 
        .QN(P1_add_468_n4) );
  NOR2X0 P1_add_468_U3 ( .QN(P1_add_468_n1), .IN1(P1_add_468_n3), 
        .IN2(P1_add_468_n4) );
  AND2X1 P1_add_468_U2 ( .IN1(P1_add_468_n3), .IN2(P1_add_468_n4), 
        .Q(P1_add_468_n2) );
  NOR2X0 P1_add_468_U1 ( .QN(P1_N4101), .IN1(P1_add_468_n1), 
        .IN2(P1_add_468_n2) );
  NAND2X0 P1_add_468_U149 ( .IN1(P1_N3870), .IN2(n7095), .QN(P1_add_468_n142)
         );
  NAND2X0 P1_add_468_U148 ( .IN1(P1_add_468_n141), .IN2(P1_add_468_n142), 
        .QN(P1_add_468_n140) );
  NOR2X0 P1_add_468_U147 ( .QN(P1_add_468_n138), .IN1(P1_add_468_n137), 
        .IN2(P1_add_468_n140) );
  AND2X1 P1_add_468_U146 ( .IN1(P1_add_468_n137), .IN2(P1_add_468_n140), 
        .Q(P1_add_468_n139) );
  NOR2X0 P1_add_468_U145 ( .QN(P1_N4112), .IN1(P1_add_468_n138), 
        .IN2(P1_add_468_n139) );
  NAND2X0 P1_add_468_U144 ( .IN1(P1_N5169), .IN2(P1_add_468_n137), 
        .QN(P1_add_468_n134) );
  OR2X1 P1_add_468_U143 ( .IN2(P1_N5169), .IN1(P1_add_468_n137), 
        .Q(P1_add_468_n136) );
  NAND2X0 P1_add_468_U142 ( .IN1(P1_N3870), .IN2(P1_add_468_n136), 
        .QN(P1_add_468_n135) );
  NAND2X0 P1_add_468_U141 ( .IN1(P1_add_468_n134), .IN2(P1_add_468_n135), 
        .QN(P1_add_468_n127) );
  OR2X1 P1_add_468_U139 ( .IN2(P1_N3871), .IN1(n7092), .Q(P1_add_468_n131) );
  NAND2X0 P1_add_468_U138 ( .IN1(P1_N3871), .IN2(n7092), .QN(P1_add_468_n132)
         );
  NAND2X0 P1_add_468_U137 ( .IN1(P1_add_468_n131), .IN2(P1_add_468_n132), 
        .QN(P1_add_468_n130) );
  NOR2X0 P1_add_468_U136 ( .QN(P1_add_468_n128), .IN1(P1_add_468_n127), 
        .IN2(P1_add_468_n130) );
  AND2X1 P1_add_468_U135 ( .IN1(P1_add_468_n127), .IN2(P1_add_468_n130), 
        .Q(P1_add_468_n129) );
  NOR2X0 P1_add_468_U134 ( .QN(P1_N4113), .IN1(P1_add_468_n128), 
        .IN2(P1_add_468_n129) );
  NAND2X0 P1_add_468_U133 ( .IN1(n7093), .IN2(P1_add_468_n127), 
        .QN(P1_add_468_n124) );
  OR2X1 P1_add_468_U132 ( .IN2(n7093), .IN1(P1_add_468_n127), 
        .Q(P1_add_468_n126) );
  NAND2X0 P1_add_468_U131 ( .IN1(P1_N3871), .IN2(P1_add_468_n126), 
        .QN(P1_add_468_n125) );
  NAND2X0 P1_add_468_U130 ( .IN1(P1_add_468_n124), .IN2(P1_add_468_n125), 
        .QN(P1_add_468_n117) );
  OR2X1 P1_add_468_U128 ( .IN2(P1_N3872), .IN1(n7090), .Q(P1_add_468_n121) );
  NAND2X0 P1_add_468_U127 ( .IN1(P1_N3872), .IN2(n7090), .QN(P1_add_468_n122)
         );
  NAND2X0 P1_add_468_U126 ( .IN1(P1_add_468_n121), .IN2(P1_add_468_n122), 
        .QN(P1_add_468_n120) );
  NOR2X0 P1_add_468_U125 ( .QN(P1_add_468_n118), .IN1(P1_add_468_n117), 
        .IN2(P1_add_468_n120) );
  AND2X1 P1_add_468_U124 ( .IN1(P1_add_468_n117), .IN2(P1_add_468_n120), 
        .Q(P1_add_468_n119) );
  NOR2X0 P1_add_468_U123 ( .QN(P1_N4114), .IN1(P1_add_468_n118), 
        .IN2(P1_add_468_n119) );
  NAND2X0 P1_add_468_U122 ( .IN1(n7089), .IN2(P1_add_468_n117), 
        .QN(P1_add_468_n114) );
  OR2X1 P1_add_468_U121 ( .IN2(n7089), .IN1(P1_add_468_n117), 
        .Q(P1_add_468_n116) );
  NAND2X0 P1_add_468_U120 ( .IN1(P1_N3872), .IN2(P1_add_468_n116), 
        .QN(P1_add_468_n115) );
  NAND2X0 P1_add_468_U119 ( .IN1(P1_add_468_n114), .IN2(P1_add_468_n115), 
        .QN(P1_add_468_n107) );
  OR2X1 P1_add_468_U117 ( .IN2(P1_N3873), .IN1(n7144), .Q(P1_add_468_n111) );
  NAND2X0 P1_add_468_U116 ( .IN1(P1_N3873), .IN2(n7144), .QN(P1_add_468_n112)
         );
  NAND2X0 P1_add_468_U115 ( .IN1(P1_add_468_n111), .IN2(P1_add_468_n112), 
        .QN(P1_add_468_n110) );
  NOR2X0 P1_add_468_U114 ( .QN(P1_add_468_n108), .IN1(P1_add_468_n107), 
        .IN2(P1_add_468_n110) );
  AND2X1 P1_add_468_U113 ( .IN1(P1_add_468_n107), .IN2(P1_add_468_n110), 
        .Q(P1_add_468_n109) );
  NOR2X0 P1_add_468_U112 ( .QN(P1_N4115), .IN1(P1_add_468_n108), 
        .IN2(P1_add_468_n109) );
  NAND2X0 P1_add_468_U111 ( .IN1(n7141), .IN2(P1_add_468_n107), 
        .QN(P1_add_468_n104) );
  OR2X1 P1_add_468_U110 ( .IN2(n7141), .IN1(P1_add_468_n107), 
        .Q(P1_add_468_n106) );
  NAND2X0 P1_add_468_U109 ( .IN1(P1_N3873), .IN2(P1_add_468_n106), 
        .QN(P1_add_468_n105) );
  NAND2X0 P1_add_468_U108 ( .IN1(P1_add_468_n104), .IN2(P1_add_468_n105), 
        .QN(P1_add_468_n97) );
  OR2X1 P1_add_468_U106 ( .IN2(P1_N3874), .IN1(n7136), .Q(P1_add_468_n101) );
  NAND2X0 P1_add_468_U105 ( .IN1(P1_N3874), .IN2(n7136), .QN(P1_add_468_n102)
         );
  NAND2X0 P1_add_468_U104 ( .IN1(P1_add_468_n101), .IN2(P1_add_468_n102), 
        .QN(P1_add_468_n100) );
  NOR2X0 P1_add_468_U103 ( .QN(P1_add_468_n98), .IN1(P1_add_468_n97), 
        .IN2(P1_add_468_n100) );
  AND2X1 P1_add_468_U102 ( .IN1(P1_add_468_n97), .IN2(P1_add_468_n100), 
        .Q(P1_add_468_n99) );
  NOR2X0 P1_add_468_U101 ( .QN(P1_N4116), .IN1(P1_add_468_n98), 
        .IN2(P1_add_468_n99) );
  NAND2X0 P1_add_468_U100 ( .IN1(P1_N5173), .IN2(P1_add_468_n97), 
        .QN(P1_add_468_n94) );
  OR2X1 P1_add_468_U99 ( .IN2(P1_N5173), .IN1(P1_add_468_n97), 
        .Q(P1_add_468_n96) );
  NAND2X0 P1_add_468_U98 ( .IN1(P1_N3874), .IN2(P1_add_468_n96), 
        .QN(P1_add_468_n95) );
  NAND2X0 P1_add_468_U97 ( .IN1(P1_add_468_n94), .IN2(P1_add_468_n95), 
        .QN(P1_add_468_n87) );
  OR2X1 P1_add_468_U95 ( .IN2(P1_N3875), .IN1(n7130), .Q(P1_add_468_n91) );
  NAND2X0 P1_add_468_U94 ( .IN1(P1_N3875), .IN2(n7130), .QN(P1_add_468_n92) );
  NAND2X0 P1_add_468_U93 ( .IN1(P1_add_468_n91), .IN2(P1_add_468_n92), 
        .QN(P1_add_468_n90) );
  NOR2X0 P1_add_468_U92 ( .QN(P1_add_468_n88), .IN1(P1_add_468_n87), 
        .IN2(P1_add_468_n90) );
  AND2X1 P1_add_468_U91 ( .IN1(P1_add_468_n87), .IN2(P1_add_468_n90), 
        .Q(P1_add_468_n89) );
  NOR2X0 P1_add_468_U90 ( .QN(P1_N4117), .IN1(P1_add_468_n88), 
        .IN2(P1_add_468_n89) );
  NAND2X0 P1_add_468_U89 ( .IN1(n7129), .IN2(P1_add_468_n87), 
        .QN(P1_add_468_n84) );
  OR2X1 P1_add_468_U88 ( .IN2(n7129), .IN1(P1_add_468_n87), .Q(P1_add_468_n86)
         );
  NAND2X0 P1_add_468_U87 ( .IN1(P1_N3875), .IN2(P1_add_468_n86), 
        .QN(P1_add_468_n85) );
  NAND2X0 P1_add_468_U86 ( .IN1(P1_add_468_n84), .IN2(P1_add_468_n85), 
        .QN(P1_add_468_n77) );
  OR2X1 P1_add_468_U84 ( .IN2(P1_N3876), .IN1(n7125), .Q(P1_add_468_n81) );
  NAND2X0 P1_add_468_U83 ( .IN1(P1_N3876), .IN2(n7125), .QN(P1_add_468_n82) );
  NAND2X0 P1_add_468_U82 ( .IN1(P1_add_468_n81), .IN2(P1_add_468_n82), 
        .QN(P1_add_468_n80) );
  NOR2X0 P1_add_468_U81 ( .QN(P1_add_468_n78), .IN1(P1_add_468_n77), 
        .IN2(P1_add_468_n80) );
  AND2X1 P1_add_468_U80 ( .IN1(P1_add_468_n77), .IN2(P1_add_468_n80), 
        .Q(P1_add_468_n79) );
  NOR2X0 P1_add_468_U79 ( .QN(P1_N4118), .IN1(P1_add_468_n78), 
        .IN2(P1_add_468_n79) );
  NAND2X0 P1_add_468_U78 ( .IN1(P1_N5175), .IN2(P1_add_468_n77), 
        .QN(P1_add_468_n74) );
  OR2X1 P1_add_468_U77 ( .IN2(P1_N5175), .IN1(P1_add_468_n77), 
        .Q(P1_add_468_n76) );
  NAND2X0 P1_add_468_U76 ( .IN1(P1_N3876), .IN2(P1_add_468_n76), 
        .QN(P1_add_468_n75) );
  NAND2X0 P1_add_468_U75 ( .IN1(P1_add_468_n74), .IN2(P1_add_468_n75), 
        .QN(P1_add_468_n64) );
  OR2X1 P1_add_468_U73 ( .IN2(P1_N3877), .IN1(n7119), .Q(P1_add_468_n71) );
  NAND2X0 P1_add_468_U72 ( .IN1(P1_N3877), .IN2(n7119), .QN(P1_add_468_n72) );
  NAND2X0 P1_add_468_U71 ( .IN1(P1_add_468_n71), .IN2(P1_add_468_n72), 
        .QN(P1_add_468_n70) );
  NOR2X0 P1_add_468_U70 ( .QN(P1_add_468_n68), .IN1(P1_add_468_n64), 
        .IN2(P1_add_468_n70) );
  AND2X1 P1_add_468_U69 ( .IN1(P1_add_468_n64), .IN2(P1_add_468_n70), 
        .Q(P1_add_468_n69) );
  NOR2X0 P1_add_468_U68 ( .QN(P1_N4119), .IN1(P1_add_468_n68), 
        .IN2(P1_add_468_n69) );
  OR2X1 P1_add_468_U66 ( .IN2(P1_N3878), .IN1(n7117), .Q(P1_add_468_n65) );
  NAND2X0 P1_add_468_U65 ( .IN1(P1_N3878), .IN2(n7117), .QN(P1_add_468_n66) );
  NAND2X0 P1_add_468_U64 ( .IN1(P1_add_468_n65), .IN2(P1_add_468_n66), 
        .QN(P1_add_468_n60) );
  NAND2X0 P1_add_468_U63 ( .IN1(P1_N5176), .IN2(P1_add_468_n64), 
        .QN(P1_add_468_n61) );
  OR2X1 P1_add_468_U62 ( .IN2(P1_N5176), .IN1(P1_add_468_n64), 
        .Q(P1_add_468_n63) );
  NAND2X0 P1_add_468_U61 ( .IN1(P1_N3877), .IN2(P1_add_468_n63), 
        .QN(P1_add_468_n62) );
  NAND2X0 P1_add_468_U60 ( .IN1(P1_add_468_n61), .IN2(P1_add_468_n62), 
        .QN(P1_add_468_n59) );
  NOR2X0 P1_add_468_U59 ( .QN(P1_add_468_n57), .IN1(P1_add_468_n60), 
        .IN2(P1_add_468_n59) );
  AND2X1 P1_add_468_U58 ( .IN1(P1_add_468_n59), .IN2(P1_add_468_n60), 
        .Q(P1_add_468_n58) );
  NOR2X0 P1_add_468_U57 ( .QN(P1_N4120), .IN1(P1_add_468_n57), 
        .IN2(P1_add_468_n58) );
  NAND2X0 P1_add_468_U242 ( .IN1(P1_add_468_n228), .IN2(P1_add_468_n229), 
        .QN(P1_add_468_n227) );
  NOR2X0 P1_add_468_U241 ( .QN(P1_add_468_n225), .IN1(P1_add_468_n224), 
        .IN2(P1_add_468_n227) );
  AND2X1 P1_add_468_U240 ( .IN1(P1_add_468_n224), .IN2(P1_add_468_n227), 
        .Q(P1_add_468_n226) );
  NOR2X0 P1_add_468_U239 ( .QN(P1_N4104), .IN1(P1_add_468_n225), 
        .IN2(P1_add_468_n226) );
  NAND2X0 P1_add_468_U238 ( .IN1(P1_N5161), .IN2(P1_add_468_n224), 
        .QN(P1_add_468_n221) );
  OR2X1 P1_add_468_U237 ( .IN2(P1_N5161), .IN1(P1_add_468_n224), 
        .Q(P1_add_468_n223) );
  NAND2X0 P1_add_468_U236 ( .IN1(P1_N3862), .IN2(P1_add_468_n223), 
        .QN(P1_add_468_n222) );
  NAND2X0 P1_add_468_U235 ( .IN1(P1_add_468_n221), .IN2(P1_add_468_n222), 
        .QN(P1_add_468_n214) );
  OR2X1 P1_add_468_U233 ( .IN2(P1_N3863), .IN1(n7056), .Q(P1_add_468_n218) );
  NAND2X0 P1_add_468_U232 ( .IN1(P1_N3863), .IN2(n7056), .QN(P1_add_468_n219)
         );
  NAND2X0 P1_add_468_U231 ( .IN1(P1_add_468_n218), .IN2(P1_add_468_n219), 
        .QN(P1_add_468_n217) );
  NOR2X0 P1_add_468_U230 ( .QN(P1_add_468_n215), .IN1(P1_add_468_n214), 
        .IN2(P1_add_468_n217) );
  AND2X1 P1_add_468_U229 ( .IN1(P1_add_468_n214), .IN2(P1_add_468_n217), 
        .Q(P1_add_468_n216) );
  NOR2X0 P1_add_468_U228 ( .QN(P1_N4105), .IN1(P1_add_468_n215), 
        .IN2(P1_add_468_n216) );
  NAND2X0 P1_add_468_U227 ( .IN1(P1_N5162), .IN2(P1_add_468_n214), 
        .QN(P1_add_468_n211) );
  OR2X1 P1_add_468_U226 ( .IN2(P1_N5162), .IN1(P1_add_468_n214), 
        .Q(P1_add_468_n213) );
  NAND2X0 P1_add_468_U225 ( .IN1(P1_N3863), .IN2(P1_add_468_n213), 
        .QN(P1_add_468_n212) );
  NAND2X0 P1_add_468_U224 ( .IN1(P1_add_468_n211), .IN2(P1_add_468_n212), 
        .QN(P1_add_468_n204) );
  OR2X1 P1_add_468_U222 ( .IN2(P1_N3864), .IN1(n7115), .Q(P1_add_468_n208) );
  NAND2X0 P1_add_468_U221 ( .IN1(P1_N3864), .IN2(n7115), .QN(P1_add_468_n209)
         );
  NAND2X0 P1_add_468_U220 ( .IN1(P1_add_468_n208), .IN2(P1_add_468_n209), 
        .QN(P1_add_468_n207) );
  NOR2X0 P1_add_468_U219 ( .QN(P1_add_468_n205), .IN1(P1_add_468_n204), 
        .IN2(P1_add_468_n207) );
  AND2X1 P1_add_468_U218 ( .IN1(P1_add_468_n204), .IN2(P1_add_468_n207), 
        .Q(P1_add_468_n206) );
  NOR2X0 P1_add_468_U217 ( .QN(P1_N4106), .IN1(P1_add_468_n205), 
        .IN2(P1_add_468_n206) );
  NAND2X0 P1_add_468_U216 ( .IN1(P1_N5163), .IN2(P1_add_468_n204), 
        .QN(P1_add_468_n201) );
  OR2X1 P1_add_468_U215 ( .IN2(P1_N5163), .IN1(P1_add_468_n204), 
        .Q(P1_add_468_n203) );
  NAND2X0 P1_add_468_U214 ( .IN1(P1_N3864), .IN2(P1_add_468_n203), 
        .QN(P1_add_468_n202) );
  NAND2X0 P1_add_468_U213 ( .IN1(P1_add_468_n201), .IN2(P1_add_468_n202), 
        .QN(P1_add_468_n194) );
  OR2X1 P1_add_468_U211 ( .IN2(P1_N3865), .IN1(n7112), .Q(P1_add_468_n198) );
  NAND2X0 P1_add_468_U210 ( .IN1(P1_N3865), .IN2(n7112), .QN(P1_add_468_n199)
         );
  NAND2X0 P1_add_468_U209 ( .IN1(P1_add_468_n198), .IN2(P1_add_468_n199), 
        .QN(P1_add_468_n197) );
  NOR2X0 P1_add_468_U208 ( .QN(P1_add_468_n195), .IN1(P1_add_468_n194), 
        .IN2(P1_add_468_n197) );
  AND2X1 P1_add_468_U207 ( .IN1(P1_add_468_n194), .IN2(P1_add_468_n197), 
        .Q(P1_add_468_n196) );
  NOR2X0 P1_add_468_U206 ( .QN(P1_N4107), .IN1(P1_add_468_n195), 
        .IN2(P1_add_468_n196) );
  NAND2X0 P1_add_468_U205 ( .IN1(P1_N5164), .IN2(P1_add_468_n194), 
        .QN(P1_add_468_n191) );
  OR2X1 P1_add_468_U204 ( .IN2(P1_N5164), .IN1(P1_add_468_n194), 
        .Q(P1_add_468_n193) );
  NAND2X0 P1_add_468_U203 ( .IN1(P1_N3865), .IN2(P1_add_468_n193), 
        .QN(P1_add_468_n192) );
  NAND2X0 P1_add_468_U202 ( .IN1(P1_add_468_n191), .IN2(P1_add_468_n192), 
        .QN(P1_add_468_n184) );
  OR2X1 P1_add_468_U200 ( .IN2(P1_N3866), .IN1(n7109), .Q(P1_add_468_n188) );
  NAND2X0 P1_add_468_U199 ( .IN1(P1_N3866), .IN2(n7109), .QN(P1_add_468_n189)
         );
  NAND2X0 P1_add_468_U198 ( .IN1(P1_add_468_n188), .IN2(P1_add_468_n189), 
        .QN(P1_add_468_n187) );
  NOR2X0 P1_add_468_U197 ( .QN(P1_add_468_n185), .IN1(P1_add_468_n184), 
        .IN2(P1_add_468_n187) );
  AND2X1 P1_add_468_U196 ( .IN1(P1_add_468_n184), .IN2(P1_add_468_n187), 
        .Q(P1_add_468_n186) );
  NOR2X0 P1_add_468_U195 ( .QN(P1_N4108), .IN1(P1_add_468_n185), 
        .IN2(P1_add_468_n186) );
  NAND2X0 P1_add_468_U194 ( .IN1(n7110), .IN2(P1_add_468_n184), 
        .QN(P1_add_468_n181) );
  OR2X1 P1_add_468_U193 ( .IN2(n7110), .IN1(P1_add_468_n184), 
        .Q(P1_add_468_n183) );
  NAND2X0 P1_add_468_U192 ( .IN1(P1_N3866), .IN2(P1_add_468_n183), 
        .QN(P1_add_468_n182) );
  NAND2X0 P1_add_468_U191 ( .IN1(P1_add_468_n181), .IN2(P1_add_468_n182), 
        .QN(P1_add_468_n174) );
  OR2X1 P1_add_468_U189 ( .IN2(P1_N3867), .IN1(n7105), .Q(P1_add_468_n178) );
  NAND2X0 P1_add_468_U188 ( .IN1(P1_N3867), .IN2(n7105), .QN(P1_add_468_n179)
         );
  NAND2X0 P1_add_468_U187 ( .IN1(P1_add_468_n178), .IN2(P1_add_468_n179), 
        .QN(P1_add_468_n177) );
  NOR2X0 P1_add_468_U186 ( .QN(P1_add_468_n175), .IN1(P1_add_468_n174), 
        .IN2(P1_add_468_n177) );
  AND2X1 P1_add_468_U185 ( .IN1(P1_add_468_n174), .IN2(P1_add_468_n177), 
        .Q(P1_add_468_n176) );
  NOR2X0 P1_add_468_U184 ( .QN(P1_N4109), .IN1(P1_add_468_n175), 
        .IN2(P1_add_468_n176) );
  NAND2X0 P1_add_468_U183 ( .IN1(P1_N5166), .IN2(P1_add_468_n174), 
        .QN(P1_add_468_n171) );
  OR2X1 P1_add_468_U182 ( .IN2(P1_N5166), .IN1(P1_add_468_n174), 
        .Q(P1_add_468_n173) );
  NAND2X0 P1_add_468_U181 ( .IN1(P1_N3867), .IN2(P1_add_468_n173), 
        .QN(P1_add_468_n172) );
  NAND2X0 P1_add_468_U180 ( .IN1(P1_add_468_n171), .IN2(P1_add_468_n172), 
        .QN(P1_add_468_n164) );
  OR2X1 P1_add_468_U178 ( .IN2(P1_N3868), .IN1(n7102), .Q(P1_add_468_n168) );
  NAND2X0 P1_add_468_U177 ( .IN1(P1_N3868), .IN2(n7102), .QN(P1_add_468_n169)
         );
  NAND2X0 P1_add_468_U176 ( .IN1(P1_add_468_n168), .IN2(P1_add_468_n169), 
        .QN(P1_add_468_n167) );
  NOR2X0 P1_add_468_U175 ( .QN(P1_add_468_n165), .IN1(P1_add_468_n164), 
        .IN2(P1_add_468_n167) );
  AND2X1 P1_add_468_U174 ( .IN1(P1_add_468_n164), .IN2(P1_add_468_n167), 
        .Q(P1_add_468_n166) );
  NOR2X0 P1_add_468_U173 ( .QN(P1_N4110), .IN1(P1_add_468_n165), 
        .IN2(P1_add_468_n166) );
  NAND2X0 P1_add_468_U172 ( .IN1(n7103), .IN2(P1_add_468_n164), 
        .QN(P1_add_468_n161) );
  OR2X1 P1_add_468_U171 ( .IN2(n7103), .IN1(P1_add_468_n164), 
        .Q(P1_add_468_n163) );
  NAND2X0 P1_add_468_U170 ( .IN1(P1_N3868), .IN2(P1_add_468_n163), 
        .QN(P1_add_468_n162) );
  NAND2X0 P1_add_468_U169 ( .IN1(P1_add_468_n161), .IN2(P1_add_468_n162), 
        .QN(P1_add_468_n147) );
  OR2X1 P1_add_468_U167 ( .IN2(P1_N3869), .IN1(n7098), .Q(P1_add_468_n158) );
  NAND2X0 P1_add_468_U166 ( .IN1(P1_N3869), .IN2(n7098), .QN(P1_add_468_n159)
         );
  NAND2X0 P1_add_468_U165 ( .IN1(P1_add_468_n158), .IN2(P1_add_468_n159), 
        .QN(P1_add_468_n157) );
  NOR2X0 P1_add_468_U164 ( .QN(P1_add_468_n155), .IN1(P1_add_468_n147), 
        .IN2(P1_add_468_n157) );
  AND2X1 P1_add_468_U163 ( .IN1(P1_add_468_n147), .IN2(P1_add_468_n157), 
        .Q(P1_add_468_n156) );
  NOR2X0 P1_add_468_U162 ( .QN(P1_N4111), .IN1(P1_add_468_n155), 
        .IN2(P1_add_468_n156) );
  OR2X1 P1_add_468_U161 ( .IN2(P1_N3851), .IN1(n7051), .Q(P1_add_468_n152) );
  NAND2X0 P1_add_468_U160 ( .IN1(P1_N3851), .IN2(n7051), .QN(P1_add_468_n153)
         );
  NAND2X0 P1_add_468_U159 ( .IN1(P1_add_468_n152), .IN2(P1_add_468_n153), 
        .QN(P1_add_468_n150) );
  NAND2X0 P1_add_468_U158 ( .IN1(P1_add_468_n150), .IN2(P1_add_468_n151), 
        .QN(P1_add_468_n148) );
  OR2X1 P1_add_468_U157 ( .IN2(P1_add_468_n151), .IN1(P1_add_468_n150), 
        .Q(P1_add_468_n149) );
  NAND2X0 P1_add_468_U156 ( .IN1(P1_add_468_n148), .IN2(P1_add_468_n149), 
        .QN(P1_N4093) );
  NAND2X0 P1_add_468_U155 ( .IN1(n7099), .IN2(P1_add_468_n147), 
        .QN(P1_add_468_n144) );
  OR2X1 P1_add_468_U154 ( .IN2(n7099), .IN1(P1_add_468_n147), 
        .Q(P1_add_468_n146) );
  NAND2X0 P1_add_468_U153 ( .IN1(P1_N3869), .IN2(P1_add_468_n146), 
        .QN(P1_add_468_n145) );
  NAND2X0 P1_add_468_U152 ( .IN1(P1_add_468_n144), .IN2(P1_add_468_n145), 
        .QN(P1_add_468_n137) );
  OR2X1 P1_add_468_U150 ( .IN2(P1_N3870), .IN1(n7095), .Q(P1_add_468_n141) );
  OR2X1 P1_add_468_U308 ( .IN2(P1_N3850), .IN1(n4803), .Q(P1_add_468_n278) );
  NAND2X0 P1_add_468_U307 ( .IN1(P1_N3850), .IN2(n4803), .QN(P1_add_468_n279)
         );
  NAND2X0 P1_add_468_U306 ( .IN1(P1_add_468_n278), .IN2(P1_add_468_n279), 
        .QN(P1_N4092) );
  NAND2X0 P1_add_468_U304 ( .IN1(P1_N3850), .IN2(n7034), .QN(P1_add_468_n151)
         );
  OR2X1 P1_add_468_U303 ( .IN2(P1_add_468_n151), .IN1(n7051), 
        .Q(P1_add_468_n275) );
  NAND2X0 P1_add_468_U302 ( .IN1(n7051), .IN2(P1_add_468_n151), 
        .QN(P1_add_468_n277) );
  NAND2X0 P1_add_468_U301 ( .IN1(P1_N3851), .IN2(P1_add_468_n277), 
        .QN(P1_add_468_n276) );
  NAND2X0 P1_add_468_U300 ( .IN1(P1_add_468_n275), .IN2(P1_add_468_n276), 
        .QN(P1_add_468_n52) );
  NAND2X0 P1_add_468_U299 ( .IN1(P1_N5151), .IN2(P1_add_468_n52), 
        .QN(P1_add_468_n272) );
  OR2X1 P1_add_468_U298 ( .IN2(P1_N5151), .IN1(P1_add_468_n52), 
        .Q(P1_add_468_n274) );
  NAND2X0 P1_add_468_U297 ( .IN1(P1_N3852), .IN2(P1_add_468_n274), 
        .QN(P1_add_468_n273) );
  NAND2X0 P1_add_468_U296 ( .IN1(P1_add_468_n272), .IN2(P1_add_468_n273), 
        .QN(P1_add_468_n45) );
  NAND2X0 P1_add_468_U295 ( .IN1(n7041), .IN2(P1_add_468_n45), 
        .QN(P1_add_468_n269) );
  OR2X1 P1_add_468_U294 ( .IN2(n7041), .IN1(P1_add_468_n45), 
        .Q(P1_add_468_n271) );
  NAND2X0 P1_add_468_U293 ( .IN1(P1_N3853), .IN2(P1_add_468_n271), 
        .QN(P1_add_468_n270) );
  NAND2X0 P1_add_468_U292 ( .IN1(P1_add_468_n269), .IN2(P1_add_468_n270), 
        .QN(P1_add_468_n38) );
  NAND2X0 P1_add_468_U291 ( .IN1(n7036), .IN2(P1_add_468_n38), 
        .QN(P1_add_468_n266) );
  OR2X1 P1_add_468_U290 ( .IN2(n7036), .IN1(P1_add_468_n38), 
        .Q(P1_add_468_n268) );
  NAND2X0 P1_add_468_U289 ( .IN1(P1_N3854), .IN2(P1_add_468_n268), 
        .QN(P1_add_468_n267) );
  NAND2X0 P1_add_468_U288 ( .IN1(P1_add_468_n266), .IN2(P1_add_468_n267), 
        .QN(P1_add_468_n31) );
  NAND2X0 P1_add_468_U287 ( .IN1(n7081), .IN2(P1_add_468_n31), 
        .QN(P1_add_468_n263) );
  OR2X1 P1_add_468_U286 ( .IN2(n7081), .IN1(P1_add_468_n31), 
        .Q(P1_add_468_n265) );
  NAND2X0 P1_add_468_U285 ( .IN1(P1_N3855), .IN2(P1_add_468_n265), 
        .QN(P1_add_468_n264) );
  NAND2X0 P1_add_468_U284 ( .IN1(P1_add_468_n263), .IN2(P1_add_468_n264), 
        .QN(P1_add_468_n24) );
  NAND2X0 P1_add_468_U283 ( .IN1(n7080), .IN2(P1_add_468_n24), 
        .QN(P1_add_468_n260) );
  OR2X1 P1_add_468_U282 ( .IN2(P1_N5155), .IN1(P1_add_468_n24), 
        .Q(P1_add_468_n262) );
  NAND2X0 P1_add_468_U281 ( .IN1(P1_N3856), .IN2(P1_add_468_n262), 
        .QN(P1_add_468_n261) );
  NAND2X0 P1_add_468_U280 ( .IN1(P1_add_468_n260), .IN2(P1_add_468_n261), 
        .QN(P1_add_468_n17) );
  NAND2X0 P1_add_468_U279 ( .IN1(n7075), .IN2(P1_add_468_n17), 
        .QN(P1_add_468_n257) );
  OR2X1 P1_add_468_U278 ( .IN2(n7075), .IN1(P1_add_468_n17), 
        .Q(P1_add_468_n259) );
  NAND2X0 P1_add_468_U277 ( .IN1(P1_N3857), .IN2(P1_add_468_n259), 
        .QN(P1_add_468_n258) );
  NAND2X0 P1_add_468_U276 ( .IN1(P1_add_468_n257), .IN2(P1_add_468_n258), 
        .QN(P1_add_468_n10) );
  NAND2X0 P1_add_468_U275 ( .IN1(n7072), .IN2(P1_add_468_n10), 
        .QN(P1_add_468_n254) );
  OR2X1 P1_add_468_U274 ( .IN2(n7072), .IN1(P1_add_468_n10), 
        .Q(P1_add_468_n256) );
  NAND2X0 P1_add_468_U273 ( .IN1(P1_N3858), .IN2(P1_add_468_n256), 
        .QN(P1_add_468_n255) );
  NAND2X0 P1_add_468_U272 ( .IN1(P1_add_468_n254), .IN2(P1_add_468_n255), 
        .QN(P1_add_468_n3) );
  NAND2X0 P1_add_468_U271 ( .IN1(P1_N5158), .IN2(P1_add_468_n3), 
        .QN(P1_add_468_n251) );
  OR2X1 P1_add_468_U270 ( .IN2(P1_N5158), .IN1(P1_add_468_n3), 
        .Q(P1_add_468_n253) );
  NAND2X0 P1_add_468_U269 ( .IN1(P1_N3859), .IN2(P1_add_468_n253), 
        .QN(P1_add_468_n252) );
  NAND2X0 P1_add_468_U268 ( .IN1(P1_add_468_n251), .IN2(P1_add_468_n252), 
        .QN(P1_add_468_n244) );
  OR2X1 P1_add_468_U266 ( .IN2(P1_N3860), .IN1(n7067), .Q(P1_add_468_n248) );
  NAND2X0 P1_add_468_U265 ( .IN1(P1_N3860), .IN2(n7067), .QN(P1_add_468_n249)
         );
  NAND2X0 P1_add_468_U264 ( .IN1(P1_add_468_n248), .IN2(P1_add_468_n249), 
        .QN(P1_add_468_n247) );
  NOR2X0 P1_add_468_U263 ( .QN(P1_add_468_n245), .IN1(P1_add_468_n244), 
        .IN2(P1_add_468_n247) );
  AND2X1 P1_add_468_U262 ( .IN1(P1_add_468_n244), .IN2(P1_add_468_n247), 
        .Q(P1_add_468_n246) );
  NOR2X0 P1_add_468_U261 ( .QN(P1_N4102), .IN1(P1_add_468_n245), 
        .IN2(P1_add_468_n246) );
  NAND2X0 P1_add_468_U260 ( .IN1(P1_N5159), .IN2(P1_add_468_n244), 
        .QN(P1_add_468_n241) );
  OR2X1 P1_add_468_U259 ( .IN2(P1_N5159), .IN1(P1_add_468_n244), 
        .Q(P1_add_468_n243) );
  NAND2X0 P1_add_468_U258 ( .IN1(P1_N3860), .IN2(P1_add_468_n243), 
        .QN(P1_add_468_n242) );
  NAND2X0 P1_add_468_U257 ( .IN1(P1_add_468_n241), .IN2(P1_add_468_n242), 
        .QN(P1_add_468_n234) );
  OR2X1 P1_add_468_U255 ( .IN2(P1_N3861), .IN1(n7063), .Q(P1_add_468_n238) );
  NAND2X0 P1_add_468_U254 ( .IN1(P1_N3861), .IN2(n7063), .QN(P1_add_468_n239)
         );
  NAND2X0 P1_add_468_U253 ( .IN1(P1_add_468_n238), .IN2(P1_add_468_n239), 
        .QN(P1_add_468_n237) );
  NOR2X0 P1_add_468_U252 ( .QN(P1_add_468_n235), .IN1(P1_add_468_n234), 
        .IN2(P1_add_468_n237) );
  AND2X1 P1_add_468_U251 ( .IN1(P1_add_468_n234), .IN2(P1_add_468_n237), 
        .Q(P1_add_468_n236) );
  NOR2X0 P1_add_468_U250 ( .QN(P1_N4103), .IN1(P1_add_468_n235), 
        .IN2(P1_add_468_n236) );
  NAND2X0 P1_add_468_U249 ( .IN1(P1_N5160), .IN2(P1_add_468_n234), 
        .QN(P1_add_468_n231) );
  OR2X1 P1_add_468_U248 ( .IN2(P1_N5160), .IN1(P1_add_468_n234), 
        .Q(P1_add_468_n233) );
  NAND2X0 P1_add_468_U247 ( .IN1(P1_N3861), .IN2(P1_add_468_n233), 
        .QN(P1_add_468_n232) );
  NAND2X0 P1_add_468_U246 ( .IN1(P1_add_468_n231), .IN2(P1_add_468_n232), 
        .QN(P1_add_468_n224) );
  OR2X1 P1_add_468_U244 ( .IN2(P1_N3862), .IN1(n7058), .Q(P1_add_468_n228) );
  NAND2X0 P1_add_468_U243 ( .IN1(P1_N3862), .IN2(n7058), .QN(P1_add_468_n229)
         );
  OR2X1 r845_U27 ( .IN2(P2_N2611), .IN1(n7164), .Q(r845_n26) );
  NAND2X0 r845_U26 ( .IN1(P2_N2611), .IN2(n7164), .QN(r845_n27) );
  NAND2X0 r845_U25 ( .IN1(r845_n26), .IN2(r845_n27), .QN(r845_n25) );
  NOR2X0 r845_U24 ( .QN(r845_n22), .IN1(r845_n24), .IN2(r845_n25) );
  AND2X1 r845_U23 ( .IN1(r845_n24), .IN2(r845_n25), .Q(r845_n23) );
  NOR2X0 r845_U22 ( .QN(P2_N2763), .IN1(r845_n22), .IN2(r845_n23) );
  OR2X1 r845_U20 ( .IN2(P2_N2612), .IN1(n7157), .Q(r845_n19) );
  NAND2X0 r845_U19 ( .IN1(P2_N2612), .IN2(n7157), .QN(r845_n20) );
  NAND2X0 r845_U18 ( .IN1(r845_n19), .IN2(r845_n20), .QN(r845_n18) );
  NOR2X0 r845_U17 ( .QN(r845_n15), .IN1(r845_n17), .IN2(r845_n18) );
  AND2X1 r845_U16 ( .IN1(r845_n17), .IN2(r845_n18), .Q(r845_n16) );
  NOR2X0 r845_U15 ( .QN(P2_N2764), .IN1(r845_n15), .IN2(r845_n16) );
  OR2X1 r845_U13 ( .IN2(P2_N2613), .IN1(n7153), .Q(r845_n12) );
  NAND2X0 r845_U12 ( .IN1(P2_N2613), .IN2(n7153), .QN(r845_n13) );
  NAND2X0 r845_U11 ( .IN1(r845_n12), .IN2(r845_n13), .QN(r845_n11) );
  NOR2X0 r845_U10 ( .QN(r845_n8), .IN1(r845_n10), .IN2(r845_n11) );
  AND2X1 r845_U9 ( .IN1(r845_n10), .IN2(r845_n11), .Q(r845_n9) );
  NOR2X0 r845_U8 ( .QN(P2_N2765), .IN1(r845_n8), .IN2(r845_n9) );
  OR2X1 r845_U6 ( .IN2(P2_N2614), .IN1(n7149), .Q(r845_n5) );
  NAND2X0 r845_U5 ( .IN1(P2_N2614), .IN2(n7149), .QN(r845_n6) );
  NAND2X0 r845_U4 ( .IN1(r845_n5), .IN2(r845_n6), .QN(r845_n4) );
  NOR2X0 r845_U3 ( .QN(r845_n1), .IN1(r845_n3), .IN2(r845_n4) );
  AND2X1 r845_U2 ( .IN1(r845_n3), .IN2(r845_n4), .Q(r845_n2) );
  NOR2X0 r845_U1 ( .QN(P2_N2766), .IN1(r845_n1), .IN2(r845_n2) );
  NAND2X0 r845_U120 ( .IN1(P2_N2628), .IN2(r845_n116), .QN(r845_n115) );
  NAND2X0 r845_U119 ( .IN1(r845_n114), .IN2(r845_n115), .QN(r845_n107) );
  OR2X1 r845_U117 ( .IN2(P2_N2629), .IN1(n7239), .Q(r845_n111) );
  NAND2X0 r845_U116 ( .IN1(P2_N2629), .IN2(n7239), .QN(r845_n112) );
  NAND2X0 r845_U115 ( .IN1(r845_n111), .IN2(r845_n112), .QN(r845_n110) );
  NOR2X0 r845_U114 ( .QN(r845_n108), .IN1(r845_n107), .IN2(r845_n110) );
  AND2X1 r845_U113 ( .IN1(r845_n107), .IN2(r845_n110), .Q(r845_n109) );
  NOR2X0 r845_U112 ( .QN(P2_N2781), .IN1(r845_n108), .IN2(r845_n109) );
  NAND2X0 r845_U111 ( .IN1(n7238), .IN2(r845_n107), .QN(r845_n104) );
  OR2X1 r845_U110 ( .IN2(n7238), .IN1(r845_n107), .Q(r845_n106) );
  NAND2X0 r845_U109 ( .IN1(P2_N2629), .IN2(r845_n106), .QN(r845_n105) );
  NAND2X0 r845_U108 ( .IN1(r845_n104), .IN2(r845_n105), .QN(r845_n97) );
  OR2X1 r845_U106 ( .IN2(P2_N2630), .IN1(n7234), .Q(r845_n101) );
  NAND2X0 r845_U105 ( .IN1(P2_N2630), .IN2(n7234), .QN(r845_n102) );
  NAND2X0 r845_U104 ( .IN1(r845_n101), .IN2(r845_n102), .QN(r845_n100) );
  NOR2X0 r845_U103 ( .QN(r845_n98), .IN1(r845_n97), .IN2(r845_n100) );
  AND2X1 r845_U102 ( .IN1(r845_n97), .IN2(r845_n100), .Q(r845_n99) );
  NOR2X0 r845_U101 ( .QN(P2_N2782), .IN1(r845_n98), .IN2(r845_n99) );
  NAND2X0 r845_U100 ( .IN1(P2_N5096), .IN2(r845_n97), .QN(r845_n94) );
  OR2X1 r845_U99 ( .IN2(P2_N5096), .IN1(r845_n97), .Q(r845_n96) );
  NAND2X0 r845_U98 ( .IN1(P2_N2630), .IN2(r845_n96), .QN(r845_n95) );
  NAND2X0 r845_U97 ( .IN1(r845_n94), .IN2(r845_n95), .QN(r845_n87) );
  OR2X1 r845_U95 ( .IN2(P2_N2631), .IN1(n7229), .Q(r845_n91) );
  NAND2X0 r845_U94 ( .IN1(P2_N2631), .IN2(n7229), .QN(r845_n92) );
  NAND2X0 r845_U93 ( .IN1(r845_n91), .IN2(r845_n92), .QN(r845_n90) );
  NOR2X0 r845_U92 ( .QN(r845_n88), .IN1(r845_n87), .IN2(r845_n90) );
  AND2X1 r845_U91 ( .IN1(r845_n87), .IN2(r845_n90), .Q(r845_n89) );
  NOR2X0 r845_U90 ( .QN(P2_N2783), .IN1(r845_n88), .IN2(r845_n89) );
  NAND2X0 r845_U89 ( .IN1(P2_N5097), .IN2(r845_n87), .QN(r845_n84) );
  OR2X1 r845_U88 ( .IN2(P2_N5097), .IN1(r845_n87), .Q(r845_n86) );
  NAND2X0 r845_U87 ( .IN1(P2_N2631), .IN2(r845_n86), .QN(r845_n85) );
  NAND2X0 r845_U86 ( .IN1(r845_n84), .IN2(r845_n85), .QN(r845_n77) );
  OR2X1 r845_U84 ( .IN2(P2_N2632), .IN1(n7224), .Q(r845_n81) );
  NAND2X0 r845_U83 ( .IN1(P2_N2632), .IN2(n7224), .QN(r845_n82) );
  NAND2X0 r845_U82 ( .IN1(r845_n81), .IN2(r845_n82), .QN(r845_n80) );
  NOR2X0 r845_U81 ( .QN(r845_n78), .IN1(r845_n77), .IN2(r845_n80) );
  AND2X1 r845_U80 ( .IN1(r845_n77), .IN2(r845_n80), .Q(r845_n79) );
  NOR2X0 r845_U79 ( .QN(P2_N2784), .IN1(r845_n78), .IN2(r845_n79) );
  NAND2X0 r845_U78 ( .IN1(n7227), .IN2(r845_n77), .QN(r845_n74) );
  OR2X1 r845_U77 ( .IN2(P2_N5098), .IN1(r845_n77), .Q(r845_n76) );
  NAND2X0 r845_U76 ( .IN1(P2_N2632), .IN2(r845_n76), .QN(r845_n75) );
  NAND2X0 r845_U75 ( .IN1(r845_n74), .IN2(r845_n75), .QN(r845_n64) );
  OR2X1 r845_U73 ( .IN2(P2_N2633), .IN1(n7222), .Q(r845_n71) );
  NAND2X0 r845_U72 ( .IN1(P2_N2633), .IN2(n7222), .QN(r845_n72) );
  NAND2X0 r845_U71 ( .IN1(r845_n71), .IN2(r845_n72), .QN(r845_n70) );
  NOR2X0 r845_U70 ( .QN(r845_n68), .IN1(r845_n64), .IN2(r845_n70) );
  AND2X1 r845_U69 ( .IN1(r845_n64), .IN2(r845_n70), .Q(r845_n69) );
  NOR2X0 r845_U68 ( .QN(P2_N2785), .IN1(r845_n68), .IN2(r845_n69) );
  OR2X1 r845_U66 ( .IN2(P2_N2634), .IN1(n7266), .Q(r845_n65) );
  NAND2X0 r845_U65 ( .IN1(P2_N2634), .IN2(n7266), .QN(r845_n66) );
  NAND2X0 r845_U64 ( .IN1(r845_n65), .IN2(r845_n66), .QN(r845_n60) );
  NAND2X0 r845_U63 ( .IN1(P2_N5099), .IN2(r845_n64), .QN(r845_n61) );
  OR2X1 r845_U62 ( .IN2(P2_N5099), .IN1(r845_n64), .Q(r845_n63) );
  NAND2X0 r845_U61 ( .IN1(P2_N2633), .IN2(r845_n63), .QN(r845_n62) );
  NAND2X0 r845_U60 ( .IN1(r845_n61), .IN2(r845_n62), .QN(r845_n59) );
  NOR2X0 r845_U59 ( .QN(r845_n57), .IN1(r845_n60), .IN2(r845_n59) );
  AND2X1 r845_U58 ( .IN1(r845_n59), .IN2(r845_n60), .Q(r845_n58) );
  NOR2X0 r845_U57 ( .QN(P2_N2786), .IN1(r845_n57), .IN2(r845_n58) );
  OR2X1 r845_U55 ( .IN2(P2_N2607), .IN1(n7182), .Q(r845_n54) );
  NAND2X0 r845_U54 ( .IN1(P2_N2607), .IN2(n7182), .QN(r845_n55) );
  NAND2X0 r845_U53 ( .IN1(r845_n54), .IN2(r845_n55), .QN(r845_n53) );
  NOR2X0 r845_U52 ( .QN(r845_n50), .IN1(r845_n52), .IN2(r845_n53) );
  AND2X1 r845_U51 ( .IN1(r845_n52), .IN2(r845_n53), .Q(r845_n51) );
  NOR2X0 r845_U50 ( .QN(P2_N2759), .IN1(r845_n50), .IN2(r845_n51) );
  OR2X1 r845_U48 ( .IN2(P2_N2608), .IN1(n7178), .Q(r845_n47) );
  NAND2X0 r845_U47 ( .IN1(P2_N2608), .IN2(n7178), .QN(r845_n48) );
  NAND2X0 r845_U46 ( .IN1(r845_n47), .IN2(r845_n48), .QN(r845_n46) );
  NOR2X0 r845_U45 ( .QN(r845_n43), .IN1(r845_n45), .IN2(r845_n46) );
  AND2X1 r845_U44 ( .IN1(r845_n45), .IN2(r845_n46), .Q(r845_n44) );
  NOR2X0 r845_U43 ( .QN(P2_N2760), .IN1(r845_n43), .IN2(r845_n44) );
  OR2X1 r845_U41 ( .IN2(P2_N2609), .IN1(n7174), .Q(r845_n40) );
  NAND2X0 r845_U40 ( .IN1(P2_N2609), .IN2(n7174), .QN(r845_n41) );
  NAND2X0 r845_U39 ( .IN1(r845_n40), .IN2(r845_n41), .QN(r845_n39) );
  NOR2X0 r845_U38 ( .QN(r845_n36), .IN1(r845_n38), .IN2(r845_n39) );
  AND2X1 r845_U37 ( .IN1(r845_n38), .IN2(r845_n39), .Q(r845_n37) );
  NOR2X0 r845_U36 ( .QN(P2_N2761), .IN1(r845_n36), .IN2(r845_n37) );
  OR2X1 r845_U34 ( .IN2(P2_N2610), .IN1(n7166), .Q(r845_n33) );
  NAND2X0 r845_U33 ( .IN1(P2_N2610), .IN2(n7166), .QN(r845_n34) );
  NAND2X0 r845_U32 ( .IN1(r845_n33), .IN2(r845_n34), .QN(r845_n32) );
  NOR2X0 r845_U31 ( .QN(r845_n29), .IN1(r845_n31), .IN2(r845_n32) );
  AND2X1 r845_U30 ( .IN1(r845_n31), .IN2(r845_n32), .Q(r845_n30) );
  NOR2X0 r845_U29 ( .QN(P2_N2762), .IN1(r845_n29), .IN2(r845_n30) );
  NAND2X0 r845_U213 ( .IN1(r845_n201), .IN2(r845_n202), .QN(r845_n194) );
  OR2X1 r845_U211 ( .IN2(P2_N2621), .IN1(n7197), .Q(r845_n198) );
  NAND2X0 r845_U210 ( .IN1(P2_N2621), .IN2(n7197), .QN(r845_n199) );
  NAND2X0 r845_U209 ( .IN1(r845_n198), .IN2(r845_n199), .QN(r845_n197) );
  NOR2X0 r845_U208 ( .QN(r845_n195), .IN1(r845_n194), .IN2(r845_n197) );
  AND2X1 r845_U207 ( .IN1(r845_n194), .IN2(r845_n197), .Q(r845_n196) );
  NOR2X0 r845_U206 ( .QN(P2_N2773), .IN1(r845_n195), .IN2(r845_n196) );
  NAND2X0 r845_U205 ( .IN1(P2_N5087), .IN2(r845_n194), .QN(r845_n191) );
  OR2X1 r845_U204 ( .IN2(P2_N5087), .IN1(r845_n194), .Q(r845_n193) );
  NAND2X0 r845_U203 ( .IN1(P2_N2621), .IN2(r845_n193), .QN(r845_n192) );
  NAND2X0 r845_U202 ( .IN1(r845_n191), .IN2(r845_n192), .QN(r845_n184) );
  OR2X1 r845_U200 ( .IN2(P2_N2622), .IN1(n7195), .Q(r845_n188) );
  NAND2X0 r845_U199 ( .IN1(P2_N2622), .IN2(n7195), .QN(r845_n189) );
  NAND2X0 r845_U198 ( .IN1(r845_n188), .IN2(r845_n189), .QN(r845_n187) );
  NOR2X0 r845_U197 ( .QN(r845_n185), .IN1(r845_n184), .IN2(r845_n187) );
  AND2X1 r845_U196 ( .IN1(r845_n184), .IN2(r845_n187), .Q(r845_n186) );
  NOR2X0 r845_U195 ( .QN(P2_N2774), .IN1(r845_n185), .IN2(r845_n186) );
  NAND2X0 r845_U194 ( .IN1(n7194), .IN2(r845_n184), .QN(r845_n181) );
  OR2X1 r845_U193 ( .IN2(n7194), .IN1(r845_n184), .Q(r845_n183) );
  NAND2X0 r845_U192 ( .IN1(P2_N2622), .IN2(r845_n183), .QN(r845_n182) );
  NAND2X0 r845_U191 ( .IN1(r845_n181), .IN2(r845_n182), .QN(r845_n174) );
  OR2X1 r845_U189 ( .IN2(P2_N2623), .IN1(n7188), .Q(r845_n178) );
  NAND2X0 r845_U188 ( .IN1(P2_N2623), .IN2(n7188), .QN(r845_n179) );
  NAND2X0 r845_U187 ( .IN1(r845_n178), .IN2(r845_n179), .QN(r845_n177) );
  NOR2X0 r845_U186 ( .QN(r845_n175), .IN1(r845_n174), .IN2(r845_n177) );
  AND2X1 r845_U185 ( .IN1(r845_n174), .IN2(r845_n177), .Q(r845_n176) );
  NOR2X0 r845_U184 ( .QN(P2_N2775), .IN1(r845_n175), .IN2(r845_n176) );
  NAND2X0 r845_U183 ( .IN1(n7187), .IN2(r845_n174), .QN(r845_n171) );
  OR2X1 r845_U182 ( .IN2(n7187), .IN1(r845_n174), .Q(r845_n173) );
  NAND2X0 r845_U181 ( .IN1(P2_N2623), .IN2(r845_n173), .QN(r845_n172) );
  NAND2X0 r845_U180 ( .IN1(r845_n171), .IN2(r845_n172), .QN(r845_n157) );
  OR2X1 r845_U178 ( .IN2(P2_N2624), .IN1(n7264), .Q(r845_n168) );
  NAND2X0 r845_U177 ( .IN1(P2_N2624), .IN2(n7264), .QN(r845_n169) );
  NAND2X0 r845_U176 ( .IN1(r845_n168), .IN2(r845_n169), .QN(r845_n167) );
  NOR2X0 r845_U175 ( .QN(r845_n165), .IN1(r845_n157), .IN2(r845_n167) );
  AND2X1 r845_U174 ( .IN1(r845_n157), .IN2(r845_n167), .Q(r845_n166) );
  NOR2X0 r845_U173 ( .QN(P2_N2776), .IN1(r845_n165), .IN2(r845_n166) );
  OR2X1 r845_U172 ( .IN2(P2_N2606), .IN1(n7186), .Q(r845_n162) );
  NAND2X0 r845_U171 ( .IN1(P2_N2606), .IN2(n7186), .QN(r845_n163) );
  NAND2X0 r845_U170 ( .IN1(r845_n162), .IN2(r845_n163), .QN(r845_n160) );
  NAND2X0 r845_U169 ( .IN1(r845_n160), .IN2(r845_n161), .QN(r845_n158) );
  OR2X1 r845_U168 ( .IN2(r845_n161), .IN1(r845_n160), .Q(r845_n159) );
  NAND2X0 r845_U167 ( .IN1(r845_n158), .IN2(r845_n159), .QN(P2_N2758) );
  NAND2X0 r845_U166 ( .IN1(n7263), .IN2(r845_n157), .QN(r845_n154) );
  OR2X1 r845_U165 ( .IN2(n7263), .IN1(r845_n157), .Q(r845_n156) );
  NAND2X0 r845_U164 ( .IN1(P2_N2624), .IN2(r845_n156), .QN(r845_n155) );
  NAND2X0 r845_U163 ( .IN1(r845_n154), .IN2(r845_n155), .QN(r845_n147) );
  OR2X1 r845_U161 ( .IN2(P2_N2625), .IN1(n7260), .Q(r845_n151) );
  NAND2X0 r845_U160 ( .IN1(P2_N2625), .IN2(n7260), .QN(r845_n152) );
  NAND2X0 r845_U159 ( .IN1(r845_n151), .IN2(r845_n152), .QN(r845_n150) );
  NOR2X0 r845_U158 ( .QN(r845_n148), .IN1(r845_n147), .IN2(r845_n150) );
  AND2X1 r845_U157 ( .IN1(r845_n147), .IN2(r845_n150), .Q(r845_n149) );
  NOR2X0 r845_U156 ( .QN(P2_N2777), .IN1(r845_n148), .IN2(r845_n149) );
  NAND2X0 r845_U155 ( .IN1(n7259), .IN2(r845_n147), .QN(r845_n144) );
  OR2X1 r845_U154 ( .IN2(n7259), .IN1(r845_n147), .Q(r845_n146) );
  NAND2X0 r845_U153 ( .IN1(P2_N2625), .IN2(r845_n146), .QN(r845_n145) );
  NAND2X0 r845_U152 ( .IN1(r845_n144), .IN2(r845_n145), .QN(r845_n137) );
  OR2X1 r845_U150 ( .IN2(P2_N2626), .IN1(n7253), .Q(r845_n141) );
  NAND2X0 r845_U149 ( .IN1(P2_N2626), .IN2(n7253), .QN(r845_n142) );
  NAND2X0 r845_U148 ( .IN1(r845_n141), .IN2(r845_n142), .QN(r845_n140) );
  NOR2X0 r845_U147 ( .QN(r845_n138), .IN1(r845_n137), .IN2(r845_n140) );
  AND2X1 r845_U146 ( .IN1(r845_n137), .IN2(r845_n140), .Q(r845_n139) );
  NOR2X0 r845_U145 ( .QN(P2_N2778), .IN1(r845_n138), .IN2(r845_n139) );
  NAND2X0 r845_U144 ( .IN1(n7252), .IN2(r845_n137), .QN(r845_n134) );
  OR2X1 r845_U143 ( .IN2(n7252), .IN1(r845_n137), .Q(r845_n136) );
  NAND2X0 r845_U142 ( .IN1(P2_N2626), .IN2(r845_n136), .QN(r845_n135) );
  NAND2X0 r845_U141 ( .IN1(r845_n134), .IN2(r845_n135), .QN(r845_n127) );
  OR2X1 r845_U139 ( .IN2(P2_N2627), .IN1(n7248), .Q(r845_n131) );
  NAND2X0 r845_U138 ( .IN1(P2_N2627), .IN2(n7248), .QN(r845_n132) );
  NAND2X0 r845_U137 ( .IN1(r845_n131), .IN2(r845_n132), .QN(r845_n130) );
  NOR2X0 r845_U136 ( .QN(r845_n128), .IN1(r845_n127), .IN2(r845_n130) );
  AND2X1 r845_U135 ( .IN1(r845_n127), .IN2(r845_n130), .Q(r845_n129) );
  NOR2X0 r845_U134 ( .QN(P2_N2779), .IN1(r845_n128), .IN2(r845_n129) );
  NAND2X0 r845_U133 ( .IN1(P2_N5093), .IN2(r845_n127), .QN(r845_n124) );
  OR2X1 r845_U132 ( .IN2(P2_N5093), .IN1(r845_n127), .Q(r845_n126) );
  NAND2X0 r845_U131 ( .IN1(P2_N2627), .IN2(r845_n126), .QN(r845_n125) );
  NAND2X0 r845_U130 ( .IN1(r845_n124), .IN2(r845_n125), .QN(r845_n117) );
  OR2X1 r845_U128 ( .IN2(P2_N2628), .IN1(n7243), .Q(r845_n121) );
  NAND2X0 r845_U127 ( .IN1(P2_N2628), .IN2(n7243), .QN(r845_n122) );
  NAND2X0 r845_U126 ( .IN1(r845_n121), .IN2(r845_n122), .QN(r845_n120) );
  NOR2X0 r845_U125 ( .QN(r845_n118), .IN1(r845_n117), .IN2(r845_n120) );
  AND2X1 r845_U124 ( .IN1(r845_n117), .IN2(r845_n120), .Q(r845_n119) );
  NOR2X0 r845_U123 ( .QN(P2_N2780), .IN1(r845_n118), .IN2(r845_n119) );
  NAND2X0 r845_U122 ( .IN1(n7242), .IN2(r845_n117), .QN(r845_n114) );
  OR2X1 r845_U121 ( .IN2(n7242), .IN1(r845_n117), .Q(r845_n116) );
  NAND2X0 r845_U306 ( .IN1(n7177), .IN2(r845_n45), .QN(r845_n279) );
  OR2X1 r845_U305 ( .IN2(n7177), .IN1(r845_n45), .Q(r845_n281) );
  NAND2X0 r845_U304 ( .IN1(P2_N2608), .IN2(r845_n281), .QN(r845_n280) );
  NAND2X0 r845_U303 ( .IN1(r845_n279), .IN2(r845_n280), .QN(r845_n38) );
  NAND2X0 r845_U302 ( .IN1(n7173), .IN2(r845_n38), .QN(r845_n276) );
  OR2X1 r845_U301 ( .IN2(n7173), .IN1(r845_n38), .Q(r845_n278) );
  NAND2X0 r845_U300 ( .IN1(P2_N2609), .IN2(r845_n278), .QN(r845_n277) );
  NAND2X0 r845_U299 ( .IN1(r845_n276), .IN2(r845_n277), .QN(r845_n31) );
  NAND2X0 r845_U298 ( .IN1(n7165), .IN2(r845_n31), .QN(r845_n273) );
  OR2X1 r845_U297 ( .IN2(n7165), .IN1(r845_n31), .Q(r845_n275) );
  NAND2X0 r845_U296 ( .IN1(P2_N2610), .IN2(r845_n275), .QN(r845_n274) );
  NAND2X0 r845_U295 ( .IN1(r845_n273), .IN2(r845_n274), .QN(r845_n24) );
  NAND2X0 r845_U294 ( .IN1(P2_N5077), .IN2(r845_n24), .QN(r845_n270) );
  OR2X1 r845_U293 ( .IN2(P2_N5077), .IN1(r845_n24), .Q(r845_n272) );
  NAND2X0 r845_U292 ( .IN1(P2_N2611), .IN2(r845_n272), .QN(r845_n271) );
  NAND2X0 r845_U291 ( .IN1(r845_n270), .IN2(r845_n271), .QN(r845_n17) );
  NAND2X0 r845_U290 ( .IN1(P2_N5078), .IN2(r845_n17), .QN(r845_n267) );
  OR2X1 r845_U289 ( .IN2(P2_N5078), .IN1(r845_n17), .Q(r845_n269) );
  NAND2X0 r845_U288 ( .IN1(P2_N2612), .IN2(r845_n269), .QN(r845_n268) );
  NAND2X0 r845_U287 ( .IN1(r845_n267), .IN2(r845_n268), .QN(r845_n10) );
  NAND2X0 r845_U286 ( .IN1(P2_N5079), .IN2(r845_n10), .QN(r845_n264) );
  OR2X1 r845_U285 ( .IN2(P2_N5079), .IN1(r845_n10), .Q(r845_n266) );
  NAND2X0 r845_U284 ( .IN1(P2_N2613), .IN2(r845_n266), .QN(r845_n265) );
  NAND2X0 r845_U283 ( .IN1(r845_n264), .IN2(r845_n265), .QN(r845_n3) );
  NAND2X0 r845_U282 ( .IN1(P2_N5080), .IN2(r845_n3), .QN(r845_n261) );
  OR2X1 r845_U281 ( .IN2(P2_N5080), .IN1(r845_n3), .Q(r845_n263) );
  NAND2X0 r845_U280 ( .IN1(P2_N2614), .IN2(r845_n263), .QN(r845_n262) );
  NAND2X0 r845_U279 ( .IN1(r845_n261), .IN2(r845_n262), .QN(r845_n254) );
  OR2X1 r845_U277 ( .IN2(P2_N2615), .IN1(n7219), .Q(r845_n258) );
  NAND2X0 r845_U276 ( .IN1(P2_N2615), .IN2(n7219), .QN(r845_n259) );
  NAND2X0 r845_U275 ( .IN1(r845_n258), .IN2(r845_n259), .QN(r845_n257) );
  NOR2X0 r845_U274 ( .QN(r845_n255), .IN1(r845_n254), .IN2(r845_n257) );
  AND2X1 r845_U273 ( .IN1(r845_n254), .IN2(r845_n257), .Q(r845_n256) );
  NOR2X0 r845_U272 ( .QN(P2_N2767), .IN1(r845_n255), .IN2(r845_n256) );
  NAND2X0 r845_U271 ( .IN1(P2_N5081), .IN2(r845_n254), .QN(r845_n251) );
  OR2X1 r845_U270 ( .IN2(P2_N5081), .IN1(r845_n254), .Q(r845_n253) );
  NAND2X0 r845_U269 ( .IN1(P2_N2615), .IN2(r845_n253), .QN(r845_n252) );
  NAND2X0 r845_U268 ( .IN1(r845_n251), .IN2(r845_n252), .QN(r845_n244) );
  OR2X1 r845_U266 ( .IN2(P2_N2616), .IN1(n7214), .Q(r845_n248) );
  NAND2X0 r845_U265 ( .IN1(P2_N2616), .IN2(n7214), .QN(r845_n249) );
  NAND2X0 r845_U264 ( .IN1(r845_n248), .IN2(r845_n249), .QN(r845_n247) );
  NOR2X0 r845_U263 ( .QN(r845_n245), .IN1(r845_n244), .IN2(r845_n247) );
  AND2X1 r845_U262 ( .IN1(r845_n244), .IN2(r845_n247), .Q(r845_n246) );
  NOR2X0 r845_U261 ( .QN(P2_N2768), .IN1(r845_n245), .IN2(r845_n246) );
  NAND2X0 r845_U260 ( .IN1(n7216), .IN2(r845_n244), .QN(r845_n241) );
  OR2X1 r845_U259 ( .IN2(n7216), .IN1(r845_n244), .Q(r845_n243) );
  NAND2X0 r845_U258 ( .IN1(P2_N2616), .IN2(r845_n243), .QN(r845_n242) );
  NAND2X0 r845_U257 ( .IN1(r845_n241), .IN2(r845_n242), .QN(r845_n234) );
  OR2X1 r845_U255 ( .IN2(P2_N2617), .IN1(n7211), .Q(r845_n238) );
  NAND2X0 r845_U254 ( .IN1(P2_N2617), .IN2(n7211), .QN(r845_n239) );
  NAND2X0 r845_U253 ( .IN1(r845_n238), .IN2(r845_n239), .QN(r845_n237) );
  NOR2X0 r845_U252 ( .QN(r845_n235), .IN1(r845_n234), .IN2(r845_n237) );
  AND2X1 r845_U251 ( .IN1(r845_n234), .IN2(r845_n237), .Q(r845_n236) );
  NOR2X0 r845_U250 ( .QN(P2_N2769), .IN1(r845_n235), .IN2(r845_n236) );
  NAND2X0 r845_U249 ( .IN1(n7210), .IN2(r845_n234), .QN(r845_n231) );
  OR2X1 r845_U248 ( .IN2(n7210), .IN1(r845_n234), .Q(r845_n233) );
  NAND2X0 r845_U247 ( .IN1(P2_N2617), .IN2(r845_n233), .QN(r845_n232) );
  NAND2X0 r845_U246 ( .IN1(r845_n231), .IN2(r845_n232), .QN(r845_n224) );
  OR2X1 r845_U244 ( .IN2(P2_N2618), .IN1(n7208), .Q(r845_n228) );
  NAND2X0 r845_U243 ( .IN1(P2_N2618), .IN2(n7208), .QN(r845_n229) );
  NAND2X0 r845_U242 ( .IN1(r845_n228), .IN2(r845_n229), .QN(r845_n227) );
  NOR2X0 r845_U241 ( .QN(r845_n225), .IN1(r845_n224), .IN2(r845_n227) );
  AND2X1 r845_U240 ( .IN1(r845_n224), .IN2(r845_n227), .Q(r845_n226) );
  NOR2X0 r845_U239 ( .QN(P2_N2770), .IN1(r845_n225), .IN2(r845_n226) );
  NAND2X0 r845_U238 ( .IN1(P2_N5084), .IN2(r845_n224), .QN(r845_n221) );
  OR2X1 r845_U237 ( .IN2(P2_N5084), .IN1(r845_n224), .Q(r845_n223) );
  NAND2X0 r845_U236 ( .IN1(P2_N2618), .IN2(r845_n223), .QN(r845_n222) );
  NAND2X0 r845_U235 ( .IN1(r845_n221), .IN2(r845_n222), .QN(r845_n214) );
  OR2X1 r845_U233 ( .IN2(P2_N2619), .IN1(n7205), .Q(r845_n218) );
  NAND2X0 r845_U232 ( .IN1(P2_N2619), .IN2(n7205), .QN(r845_n219) );
  NAND2X0 r845_U231 ( .IN1(r845_n218), .IN2(r845_n219), .QN(r845_n217) );
  NOR2X0 r845_U230 ( .QN(r845_n215), .IN1(r845_n214), .IN2(r845_n217) );
  AND2X1 r845_U229 ( .IN1(r845_n214), .IN2(r845_n217), .Q(r845_n216) );
  NOR2X0 r845_U228 ( .QN(P2_N2771), .IN1(r845_n215), .IN2(r845_n216) );
  NAND2X0 r845_U227 ( .IN1(P2_N5085), .IN2(r845_n214), .QN(r845_n211) );
  OR2X1 r845_U226 ( .IN2(P2_N5085), .IN1(r845_n214), .Q(r845_n213) );
  NAND2X0 r845_U225 ( .IN1(P2_N2619), .IN2(r845_n213), .QN(r845_n212) );
  NAND2X0 r845_U224 ( .IN1(r845_n211), .IN2(r845_n212), .QN(r845_n204) );
  OR2X1 r845_U222 ( .IN2(P2_N2620), .IN1(n7201), .Q(r845_n208) );
  NAND2X0 r845_U221 ( .IN1(P2_N2620), .IN2(n7201), .QN(r845_n209) );
  NAND2X0 r845_U220 ( .IN1(r845_n208), .IN2(r845_n209), .QN(r845_n207) );
  NOR2X0 r845_U219 ( .QN(r845_n205), .IN1(r845_n204), .IN2(r845_n207) );
  AND2X1 r845_U218 ( .IN1(r845_n204), .IN2(r845_n207), .Q(r845_n206) );
  NOR2X0 r845_U217 ( .QN(P2_N2772), .IN1(r845_n205), .IN2(r845_n206) );
  NAND2X0 r845_U216 ( .IN1(P2_N5086), .IN2(r845_n204), .QN(r845_n201) );
  OR2X1 r845_U215 ( .IN2(P2_N5086), .IN1(r845_n204), .Q(r845_n203) );
  NAND2X0 r845_U214 ( .IN1(P2_N2620), .IN2(r845_n203), .QN(r845_n202) );
  OR2X1 r845_U319 ( .IN2(P2_N2605), .IN1(n2919), .Q(r845_n288) );
  NAND2X0 r845_U318 ( .IN1(P2_N2605), .IN2(n2919), .QN(r845_n289) );
  NAND2X0 r845_U317 ( .IN1(r845_n288), .IN2(r845_n289), .QN(P2_N2757) );
  NAND2X0 r845_U315 ( .IN1(P2_N2605), .IN2(n7035), .QN(r845_n161) );
  OR2X1 r845_U314 ( .IN2(r845_n161), .IN1(n7186), .Q(r845_n285) );
  NAND2X0 r845_U313 ( .IN1(n7186), .IN2(r845_n161), .QN(r845_n287) );
  NAND2X0 r845_U312 ( .IN1(P2_N2606), .IN2(r845_n287), .QN(r845_n286) );
  NAND2X0 r845_U311 ( .IN1(r845_n285), .IN2(r845_n286), .QN(r845_n52) );
  NAND2X0 r845_U310 ( .IN1(n7181), .IN2(r845_n52), .QN(r845_n282) );
  OR2X1 r845_U309 ( .IN2(n7181), .IN1(r845_n52), .Q(r845_n284) );
  NAND2X0 r845_U308 ( .IN1(P2_N2607), .IN2(r845_n284), .QN(r845_n283) );
  NAND2X0 r845_U307 ( .IN1(r845_n282), .IN2(r845_n283), .QN(r845_n45) );
  NAND2X0 r847_U69 ( .IN1(P2_N5099), .IN2(r847_n64), .QN(r847_n77) );
  OR2X1 r847_U68 ( .IN2(P2_N5099), .IN1(r847_n64), .Q(r847_n78) );
  NAND2X0 r847_U67 ( .IN1(r847_n77), .IN2(r847_n78), .QN(r847_n71) );
  NAND2X0 r847_U66 ( .IN1(n7227), .IN2(r847_n76), .QN(r847_n72) );
  OR2X1 r847_U65 ( .IN2(n7227), .IN1(r847_n76), .Q(r847_n74) );
  NAND2X0 r847_U64 ( .IN1(r847_n74), .IN2(r847_n75), .QN(r847_n73) );
  NAND2X0 r847_U63 ( .IN1(r847_n72), .IN2(r847_n73), .QN(r847_n65) );
  NAND2X0 r847_U62 ( .IN1(r847_n71), .IN2(r847_n65), .QN(r847_n69) );
  OR2X1 r847_U61 ( .IN2(r847_n65), .IN1(r847_n71), .Q(r847_n70) );
  NAND2X0 r847_U60 ( .IN1(r847_n69), .IN2(r847_n70), .QN(P2_N3158) );
  OR2X1 r847_U58 ( .IN2(P2_N3007), .IN1(n7266), .Q(r847_n66) );
  NAND2X0 r847_U57 ( .IN1(P2_N3007), .IN2(n7266), .QN(r847_n67) );
  NAND2X0 r847_U56 ( .IN1(r847_n66), .IN2(r847_n67), .QN(r847_n60) );
  NAND2X0 r847_U55 ( .IN1(P2_N5099), .IN2(r847_n65), .QN(r847_n61) );
  OR2X1 r847_U54 ( .IN2(P2_N5099), .IN1(r847_n65), .Q(r847_n63) );
  NAND2X0 r847_U53 ( .IN1(r847_n63), .IN2(r847_n64), .QN(r847_n62) );
  NAND2X0 r847_U52 ( .IN1(r847_n61), .IN2(r847_n62), .QN(r847_n59) );
  NAND2X0 r847_U51 ( .IN1(r847_n60), .IN2(r847_n59), .QN(r847_n57) );
  OR2X1 r847_U50 ( .IN2(r847_n60), .IN1(r847_n59), .Q(r847_n58) );
  NAND2X0 r847_U49 ( .IN1(r847_n57), .IN2(r847_n58), .QN(P2_N3159) );
  NAND2X0 r847_U48 ( .IN1(n7181), .IN2(r847_n56), .QN(r847_n54) );
  OR2X1 r847_U47 ( .IN2(n7181), .IN1(r847_n56), .Q(r847_n55) );
  NAND2X0 r847_U46 ( .IN1(r847_n54), .IN2(r847_n55), .QN(r847_n52) );
  NAND2X0 r847_U45 ( .IN1(r847_n52), .IN2(r847_n53), .QN(r847_n50) );
  OR2X1 r847_U44 ( .IN2(r847_n53), .IN1(r847_n52), .Q(r847_n51) );
  NAND2X0 r847_U43 ( .IN1(r847_n50), .IN2(r847_n51), .QN(P2_N3132) );
  NAND2X0 r847_U42 ( .IN1(P2_N5074), .IN2(r847_n49), .QN(r847_n47) );
  OR2X1 r847_U41 ( .IN2(P2_N5074), .IN1(r847_n49), .Q(r847_n48) );
  NAND2X0 r847_U40 ( .IN1(r847_n47), .IN2(r847_n48), .QN(r847_n45) );
  NAND2X0 r847_U39 ( .IN1(r847_n45), .IN2(r847_n46), .QN(r847_n43) );
  OR2X1 r847_U38 ( .IN2(r847_n46), .IN1(r847_n45), .Q(r847_n44) );
  NAND2X0 r847_U37 ( .IN1(r847_n43), .IN2(r847_n44), .QN(P2_N3133) );
  NAND2X0 r847_U36 ( .IN1(P2_N5075), .IN2(r847_n42), .QN(r847_n40) );
  OR2X1 r847_U35 ( .IN2(P2_N5075), .IN1(r847_n42), .Q(r847_n41) );
  NAND2X0 r847_U34 ( .IN1(r847_n40), .IN2(r847_n41), .QN(r847_n38) );
  NAND2X0 r847_U33 ( .IN1(r847_n38), .IN2(r847_n39), .QN(r847_n36) );
  OR2X1 r847_U32 ( .IN2(r847_n39), .IN1(r847_n38), .Q(r847_n37) );
  NAND2X0 r847_U31 ( .IN1(r847_n36), .IN2(r847_n37), .QN(P2_N3134) );
  NAND2X0 r847_U30 ( .IN1(n7165), .IN2(r847_n35), .QN(r847_n33) );
  OR2X1 r847_U29 ( .IN2(n7165), .IN1(r847_n35), .Q(r847_n34) );
  NAND2X0 r847_U28 ( .IN1(r847_n33), .IN2(r847_n34), .QN(r847_n31) );
  NAND2X0 r847_U27 ( .IN1(r847_n31), .IN2(r847_n32), .QN(r847_n29) );
  OR2X1 r847_U26 ( .IN2(r847_n32), .IN1(r847_n31), .Q(r847_n30) );
  NAND2X0 r847_U25 ( .IN1(r847_n29), .IN2(r847_n30), .QN(P2_N3135) );
  NAND2X0 r847_U24 ( .IN1(n7162), .IN2(r847_n28), .QN(r847_n26) );
  OR2X1 r847_U23 ( .IN2(n7162), .IN1(r847_n28), .Q(r847_n27) );
  NAND2X0 r847_U22 ( .IN1(r847_n26), .IN2(r847_n27), .QN(r847_n24) );
  NAND2X0 r847_U21 ( .IN1(r847_n24), .IN2(r847_n25), .QN(r847_n22) );
  OR2X1 r847_U20 ( .IN2(r847_n25), .IN1(r847_n24), .Q(r847_n23) );
  NAND2X0 r847_U19 ( .IN1(r847_n22), .IN2(r847_n23), .QN(P2_N3136) );
  NAND2X0 r847_U18 ( .IN1(n7158), .IN2(r847_n21), .QN(r847_n19) );
  OR2X1 r847_U17 ( .IN2(n7158), .IN1(r847_n21), .Q(r847_n20) );
  NAND2X0 r847_U16 ( .IN1(r847_n19), .IN2(r847_n20), .QN(r847_n17) );
  NAND2X0 r847_U15 ( .IN1(r847_n17), .IN2(r847_n18), .QN(r847_n15) );
  OR2X1 r847_U14 ( .IN2(r847_n18), .IN1(r847_n17), .Q(r847_n16) );
  NAND2X0 r847_U13 ( .IN1(r847_n15), .IN2(r847_n16), .QN(P2_N3137) );
  NAND2X0 r847_U12 ( .IN1(P2_N5079), .IN2(r847_n14), .QN(r847_n12) );
  OR2X1 r847_U11 ( .IN2(P2_N5079), .IN1(r847_n14), .Q(r847_n13) );
  NAND2X0 r847_U10 ( .IN1(r847_n12), .IN2(r847_n13), .QN(r847_n10) );
  NAND2X0 r847_U9 ( .IN1(r847_n10), .IN2(r847_n11), .QN(r847_n8) );
  OR2X1 r847_U8 ( .IN2(r847_n11), .IN1(r847_n10), .Q(r847_n9) );
  NAND2X0 r847_U7 ( .IN1(r847_n8), .IN2(r847_n9), .QN(P2_N3138) );
  NAND2X0 r847_U6 ( .IN1(n7151), .IN2(r847_n7), .QN(r847_n5) );
  OR2X1 r847_U5 ( .IN2(n7151), .IN1(r847_n7), .Q(r847_n6) );
  NAND2X0 r847_U4 ( .IN1(r847_n5), .IN2(r847_n6), .QN(r847_n3) );
  NAND2X0 r847_U3 ( .IN1(r847_n3), .IN2(r847_n4), .QN(r847_n1) );
  OR2X1 r847_U2 ( .IN2(r847_n4), .IN1(r847_n3), .Q(r847_n2) );
  NAND2X0 r847_U1 ( .IN1(r847_n1), .IN2(r847_n2), .QN(P2_N3139) );
  NAND2X0 r847_U162 ( .IN1(r847_n163), .IN2(r847_n164), .QN(r847_n161) );
  NAND2X0 r847_U161 ( .IN1(r847_n161), .IN2(r847_n162), .QN(r847_n159) );
  OR2X1 r847_U160 ( .IN2(r847_n162), .IN1(r847_n161), .Q(r847_n160) );
  NAND2X0 r847_U159 ( .IN1(r847_n159), .IN2(r847_n160), .QN(P2_N3131) );
  INVX0 r847_U158 ( .ZN(r847_n145), .INP(P2_N2998) );
  NAND2X0 r847_U157 ( .IN1(P2_N5091), .IN2(r847_n145), .QN(r847_n157) );
  OR2X1 r847_U156 ( .IN2(P2_N5091), .IN1(r847_n145), .Q(r847_n158) );
  NAND2X0 r847_U155 ( .IN1(r847_n157), .IN2(r847_n158), .QN(r847_n151) );
  NAND2X0 r847_U154 ( .IN1(P2_N5090), .IN2(r847_n156), .QN(r847_n152) );
  OR2X1 r847_U153 ( .IN2(P2_N5090), .IN1(r847_n156), .Q(r847_n154) );
  NAND2X0 r847_U152 ( .IN1(r847_n154), .IN2(r847_n155), .QN(r847_n153) );
  NAND2X0 r847_U151 ( .IN1(r847_n152), .IN2(r847_n153), .QN(r847_n146) );
  NAND2X0 r847_U150 ( .IN1(r847_n151), .IN2(r847_n146), .QN(r847_n149) );
  OR2X1 r847_U149 ( .IN2(r847_n146), .IN1(r847_n151), .Q(r847_n150) );
  NAND2X0 r847_U148 ( .IN1(r847_n149), .IN2(r847_n150), .QN(P2_N3150) );
  INVX0 r847_U147 ( .ZN(r847_n135), .INP(P2_N2999) );
  NAND2X0 r847_U146 ( .IN1(n7252), .IN2(r847_n135), .QN(r847_n147) );
  OR2X1 r847_U145 ( .IN2(n7252), .IN1(r847_n135), .Q(r847_n148) );
  NAND2X0 r847_U144 ( .IN1(r847_n147), .IN2(r847_n148), .QN(r847_n141) );
  NAND2X0 r847_U143 ( .IN1(P2_N5091), .IN2(r847_n146), .QN(r847_n142) );
  OR2X1 r847_U142 ( .IN2(P2_N5091), .IN1(r847_n146), .Q(r847_n144) );
  NAND2X0 r847_U141 ( .IN1(r847_n144), .IN2(r847_n145), .QN(r847_n143) );
  NAND2X0 r847_U140 ( .IN1(r847_n142), .IN2(r847_n143), .QN(r847_n136) );
  NAND2X0 r847_U139 ( .IN1(r847_n141), .IN2(r847_n136), .QN(r847_n139) );
  OR2X1 r847_U138 ( .IN2(r847_n136), .IN1(r847_n141), .Q(r847_n140) );
  NAND2X0 r847_U137 ( .IN1(r847_n139), .IN2(r847_n140), .QN(P2_N3151) );
  INVX0 r847_U136 ( .ZN(r847_n125), .INP(P2_N3000) );
  NAND2X0 r847_U135 ( .IN1(P2_N5093), .IN2(r847_n125), .QN(r847_n137) );
  OR2X1 r847_U134 ( .IN2(P2_N5093), .IN1(r847_n125), .Q(r847_n138) );
  NAND2X0 r847_U133 ( .IN1(r847_n137), .IN2(r847_n138), .QN(r847_n131) );
  NAND2X0 r847_U132 ( .IN1(n7252), .IN2(r847_n136), .QN(r847_n132) );
  OR2X1 r847_U131 ( .IN2(n7252), .IN1(r847_n136), .Q(r847_n134) );
  NAND2X0 r847_U130 ( .IN1(r847_n134), .IN2(r847_n135), .QN(r847_n133) );
  NAND2X0 r847_U129 ( .IN1(r847_n132), .IN2(r847_n133), .QN(r847_n126) );
  NAND2X0 r847_U128 ( .IN1(r847_n131), .IN2(r847_n126), .QN(r847_n129) );
  OR2X1 r847_U127 ( .IN2(r847_n126), .IN1(r847_n131), .Q(r847_n130) );
  NAND2X0 r847_U126 ( .IN1(r847_n129), .IN2(r847_n130), .QN(P2_N3152) );
  INVX0 r847_U125 ( .ZN(r847_n115), .INP(P2_N3001) );
  NAND2X0 r847_U124 ( .IN1(n7242), .IN2(r847_n115), .QN(r847_n127) );
  OR2X1 r847_U123 ( .IN2(n7242), .IN1(r847_n115), .Q(r847_n128) );
  NAND2X0 r847_U122 ( .IN1(r847_n127), .IN2(r847_n128), .QN(r847_n121) );
  NAND2X0 r847_U121 ( .IN1(P2_N5093), .IN2(r847_n126), .QN(r847_n122) );
  OR2X1 r847_U120 ( .IN2(P2_N5093), .IN1(r847_n126), .Q(r847_n124) );
  NAND2X0 r847_U119 ( .IN1(r847_n124), .IN2(r847_n125), .QN(r847_n123) );
  NAND2X0 r847_U118 ( .IN1(r847_n122), .IN2(r847_n123), .QN(r847_n116) );
  NAND2X0 r847_U117 ( .IN1(r847_n121), .IN2(r847_n116), .QN(r847_n119) );
  OR2X1 r847_U116 ( .IN2(r847_n116), .IN1(r847_n121), .Q(r847_n120) );
  NAND2X0 r847_U115 ( .IN1(r847_n119), .IN2(r847_n120), .QN(P2_N3153) );
  INVX0 r847_U114 ( .ZN(r847_n105), .INP(P2_N3002) );
  NAND2X0 r847_U113 ( .IN1(n7238), .IN2(r847_n105), .QN(r847_n117) );
  OR2X1 r847_U112 ( .IN2(n7238), .IN1(r847_n105), .Q(r847_n118) );
  NAND2X0 r847_U111 ( .IN1(r847_n117), .IN2(r847_n118), .QN(r847_n111) );
  NAND2X0 r847_U110 ( .IN1(n7242), .IN2(r847_n116), .QN(r847_n112) );
  OR2X1 r847_U109 ( .IN2(n7242), .IN1(r847_n116), .Q(r847_n114) );
  NAND2X0 r847_U108 ( .IN1(r847_n114), .IN2(r847_n115), .QN(r847_n113) );
  NAND2X0 r847_U107 ( .IN1(r847_n112), .IN2(r847_n113), .QN(r847_n106) );
  NAND2X0 r847_U106 ( .IN1(r847_n111), .IN2(r847_n106), .QN(r847_n109) );
  OR2X1 r847_U105 ( .IN2(r847_n106), .IN1(r847_n111), .Q(r847_n110) );
  NAND2X0 r847_U104 ( .IN1(r847_n109), .IN2(r847_n110), .QN(P2_N3154) );
  INVX0 r847_U103 ( .ZN(r847_n95), .INP(P2_N3003) );
  NAND2X0 r847_U102 ( .IN1(P2_N5096), .IN2(r847_n95), .QN(r847_n107) );
  OR2X1 r847_U101 ( .IN2(P2_N5096), .IN1(r847_n95), .Q(r847_n108) );
  NAND2X0 r847_U100 ( .IN1(r847_n107), .IN2(r847_n108), .QN(r847_n101) );
  NAND2X0 r847_U99 ( .IN1(n7238), .IN2(r847_n106), .QN(r847_n102) );
  OR2X1 r847_U98 ( .IN2(n7238), .IN1(r847_n106), .Q(r847_n104) );
  NAND2X0 r847_U97 ( .IN1(r847_n104), .IN2(r847_n105), .QN(r847_n103) );
  NAND2X0 r847_U96 ( .IN1(r847_n102), .IN2(r847_n103), .QN(r847_n96) );
  NAND2X0 r847_U95 ( .IN1(r847_n101), .IN2(r847_n96), .QN(r847_n99) );
  OR2X1 r847_U94 ( .IN2(r847_n96), .IN1(r847_n101), .Q(r847_n100) );
  NAND2X0 r847_U93 ( .IN1(r847_n99), .IN2(r847_n100), .QN(P2_N3155) );
  INVX0 r847_U92 ( .ZN(r847_n85), .INP(P2_N3004) );
  NAND2X0 r847_U91 ( .IN1(P2_N5097), .IN2(r847_n85), .QN(r847_n97) );
  OR2X1 r847_U90 ( .IN2(P2_N5097), .IN1(r847_n85), .Q(r847_n98) );
  NAND2X0 r847_U89 ( .IN1(r847_n97), .IN2(r847_n98), .QN(r847_n91) );
  NAND2X0 r847_U88 ( .IN1(P2_N5096), .IN2(r847_n96), .QN(r847_n92) );
  OR2X1 r847_U87 ( .IN2(P2_N5096), .IN1(r847_n96), .Q(r847_n94) );
  NAND2X0 r847_U86 ( .IN1(r847_n94), .IN2(r847_n95), .QN(r847_n93) );
  NAND2X0 r847_U85 ( .IN1(r847_n92), .IN2(r847_n93), .QN(r847_n86) );
  NAND2X0 r847_U84 ( .IN1(r847_n91), .IN2(r847_n86), .QN(r847_n89) );
  OR2X1 r847_U83 ( .IN2(r847_n86), .IN1(r847_n91), .Q(r847_n90) );
  NAND2X0 r847_U82 ( .IN1(r847_n89), .IN2(r847_n90), .QN(P2_N3156) );
  INVX0 r847_U81 ( .ZN(r847_n75), .INP(P2_N3005) );
  NAND2X0 r847_U80 ( .IN1(n7227), .IN2(r847_n75), .QN(r847_n87) );
  OR2X1 r847_U79 ( .IN2(n7227), .IN1(r847_n75), .Q(r847_n88) );
  NAND2X0 r847_U78 ( .IN1(r847_n87), .IN2(r847_n88), .QN(r847_n81) );
  NAND2X0 r847_U77 ( .IN1(P2_N5097), .IN2(r847_n86), .QN(r847_n82) );
  OR2X1 r847_U76 ( .IN2(P2_N5097), .IN1(r847_n86), .Q(r847_n84) );
  NAND2X0 r847_U75 ( .IN1(r847_n84), .IN2(r847_n85), .QN(r847_n83) );
  NAND2X0 r847_U74 ( .IN1(r847_n82), .IN2(r847_n83), .QN(r847_n76) );
  NAND2X0 r847_U73 ( .IN1(r847_n81), .IN2(r847_n76), .QN(r847_n79) );
  OR2X1 r847_U72 ( .IN2(r847_n76), .IN1(r847_n81), .Q(r847_n80) );
  NAND2X0 r847_U71 ( .IN1(r847_n79), .IN2(r847_n80), .QN(P2_N3157) );
  INVX0 r847_U70 ( .ZN(r847_n64), .INP(P2_N3006) );
  NAND2X0 r847_U255 ( .IN1(r847_n249), .IN2(r847_n244), .QN(r847_n247) );
  OR2X1 r847_U254 ( .IN2(r847_n244), .IN1(r847_n249), .Q(r847_n248) );
  NAND2X0 r847_U253 ( .IN1(r847_n247), .IN2(r847_n248), .QN(P2_N3141) );
  INVX0 r847_U252 ( .ZN(r847_n233), .INP(P2_N2990) );
  NAND2X0 r847_U251 ( .IN1(P2_N5083), .IN2(r847_n233), .QN(r847_n245) );
  OR2X1 r847_U250 ( .IN2(P2_N5083), .IN1(r847_n233), .Q(r847_n246) );
  NAND2X0 r847_U249 ( .IN1(r847_n245), .IN2(r847_n246), .QN(r847_n239) );
  NAND2X0 r847_U248 ( .IN1(P2_N5082), .IN2(r847_n244), .QN(r847_n240) );
  OR2X1 r847_U247 ( .IN2(P2_N5082), .IN1(r847_n244), .Q(r847_n242) );
  NAND2X0 r847_U246 ( .IN1(r847_n242), .IN2(r847_n243), .QN(r847_n241) );
  NAND2X0 r847_U245 ( .IN1(r847_n240), .IN2(r847_n241), .QN(r847_n234) );
  NAND2X0 r847_U244 ( .IN1(r847_n239), .IN2(r847_n234), .QN(r847_n237) );
  OR2X1 r847_U243 ( .IN2(r847_n234), .IN1(r847_n239), .Q(r847_n238) );
  NAND2X0 r847_U242 ( .IN1(r847_n237), .IN2(r847_n238), .QN(P2_N3142) );
  INVX0 r847_U241 ( .ZN(r847_n223), .INP(P2_N2991) );
  NAND2X0 r847_U240 ( .IN1(n7209), .IN2(r847_n223), .QN(r847_n235) );
  OR2X1 r847_U239 ( .IN2(n7209), .IN1(r847_n223), .Q(r847_n236) );
  NAND2X0 r847_U238 ( .IN1(r847_n235), .IN2(r847_n236), .QN(r847_n229) );
  NAND2X0 r847_U237 ( .IN1(P2_N5083), .IN2(r847_n234), .QN(r847_n230) );
  OR2X1 r847_U236 ( .IN2(P2_N5083), .IN1(r847_n234), .Q(r847_n232) );
  NAND2X0 r847_U235 ( .IN1(r847_n232), .IN2(r847_n233), .QN(r847_n231) );
  NAND2X0 r847_U234 ( .IN1(r847_n230), .IN2(r847_n231), .QN(r847_n224) );
  NAND2X0 r847_U233 ( .IN1(r847_n229), .IN2(r847_n224), .QN(r847_n227) );
  OR2X1 r847_U232 ( .IN2(r847_n224), .IN1(r847_n229), .Q(r847_n228) );
  NAND2X0 r847_U231 ( .IN1(r847_n227), .IN2(r847_n228), .QN(P2_N3143) );
  INVX0 r847_U230 ( .ZN(r847_n213), .INP(P2_N2992) );
  NAND2X0 r847_U229 ( .IN1(n7206), .IN2(r847_n213), .QN(r847_n225) );
  OR2X1 r847_U228 ( .IN2(n7206), .IN1(r847_n213), .Q(r847_n226) );
  NAND2X0 r847_U227 ( .IN1(r847_n225), .IN2(r847_n226), .QN(r847_n219) );
  NAND2X0 r847_U226 ( .IN1(n7209), .IN2(r847_n224), .QN(r847_n220) );
  OR2X1 r847_U225 ( .IN2(n7209), .IN1(r847_n224), .Q(r847_n222) );
  NAND2X0 r847_U224 ( .IN1(r847_n222), .IN2(r847_n223), .QN(r847_n221) );
  NAND2X0 r847_U223 ( .IN1(r847_n220), .IN2(r847_n221), .QN(r847_n214) );
  NAND2X0 r847_U222 ( .IN1(r847_n219), .IN2(r847_n214), .QN(r847_n217) );
  OR2X1 r847_U221 ( .IN2(r847_n214), .IN1(r847_n219), .Q(r847_n218) );
  NAND2X0 r847_U220 ( .IN1(r847_n217), .IN2(r847_n218), .QN(P2_N3144) );
  INVX0 r847_U219 ( .ZN(r847_n203), .INP(P2_N2993) );
  NAND2X0 r847_U218 ( .IN1(P2_N5086), .IN2(r847_n203), .QN(r847_n215) );
  OR2X1 r847_U217 ( .IN2(P2_N5086), .IN1(r847_n203), .Q(r847_n216) );
  NAND2X0 r847_U216 ( .IN1(r847_n215), .IN2(r847_n216), .QN(r847_n209) );
  NAND2X0 r847_U215 ( .IN1(n7206), .IN2(r847_n214), .QN(r847_n210) );
  OR2X1 r847_U214 ( .IN2(n7206), .IN1(r847_n214), .Q(r847_n212) );
  NAND2X0 r847_U213 ( .IN1(r847_n212), .IN2(r847_n213), .QN(r847_n211) );
  NAND2X0 r847_U212 ( .IN1(r847_n210), .IN2(r847_n211), .QN(r847_n204) );
  NAND2X0 r847_U211 ( .IN1(r847_n209), .IN2(r847_n204), .QN(r847_n207) );
  OR2X1 r847_U210 ( .IN2(r847_n204), .IN1(r847_n209), .Q(r847_n208) );
  NAND2X0 r847_U209 ( .IN1(r847_n207), .IN2(r847_n208), .QN(P2_N3145) );
  INVX0 r847_U208 ( .ZN(r847_n193), .INP(P2_N2994) );
  NAND2X0 r847_U207 ( .IN1(P2_N5087), .IN2(r847_n193), .QN(r847_n205) );
  OR2X1 r847_U206 ( .IN2(P2_N5087), .IN1(r847_n193), .Q(r847_n206) );
  NAND2X0 r847_U205 ( .IN1(r847_n205), .IN2(r847_n206), .QN(r847_n199) );
  NAND2X0 r847_U204 ( .IN1(P2_N5086), .IN2(r847_n204), .QN(r847_n200) );
  OR2X1 r847_U203 ( .IN2(P2_N5086), .IN1(r847_n204), .Q(r847_n202) );
  NAND2X0 r847_U202 ( .IN1(r847_n202), .IN2(r847_n203), .QN(r847_n201) );
  NAND2X0 r847_U201 ( .IN1(r847_n200), .IN2(r847_n201), .QN(r847_n194) );
  NAND2X0 r847_U200 ( .IN1(r847_n199), .IN2(r847_n194), .QN(r847_n197) );
  OR2X1 r847_U199 ( .IN2(r847_n194), .IN1(r847_n199), .Q(r847_n198) );
  NAND2X0 r847_U198 ( .IN1(r847_n197), .IN2(r847_n198), .QN(P2_N3146) );
  INVX0 r847_U197 ( .ZN(r847_n183), .INP(P2_N2995) );
  NAND2X0 r847_U196 ( .IN1(P2_N5088), .IN2(r847_n183), .QN(r847_n195) );
  OR2X1 r847_U195 ( .IN2(P2_N5088), .IN1(r847_n183), .Q(r847_n196) );
  NAND2X0 r847_U194 ( .IN1(r847_n195), .IN2(r847_n196), .QN(r847_n189) );
  NAND2X0 r847_U193 ( .IN1(P2_N5087), .IN2(r847_n194), .QN(r847_n190) );
  OR2X1 r847_U192 ( .IN2(P2_N5087), .IN1(r847_n194), .Q(r847_n192) );
  NAND2X0 r847_U191 ( .IN1(r847_n192), .IN2(r847_n193), .QN(r847_n191) );
  NAND2X0 r847_U190 ( .IN1(r847_n190), .IN2(r847_n191), .QN(r847_n184) );
  NAND2X0 r847_U189 ( .IN1(r847_n189), .IN2(r847_n184), .QN(r847_n187) );
  OR2X1 r847_U188 ( .IN2(r847_n184), .IN1(r847_n189), .Q(r847_n188) );
  NAND2X0 r847_U187 ( .IN1(r847_n187), .IN2(r847_n188), .QN(P2_N3147) );
  INVX0 r847_U186 ( .ZN(r847_n173), .INP(P2_N2996) );
  NAND2X0 r847_U185 ( .IN1(n7187), .IN2(r847_n173), .QN(r847_n185) );
  OR2X1 r847_U184 ( .IN2(n7187), .IN1(r847_n173), .Q(r847_n186) );
  NAND2X0 r847_U183 ( .IN1(r847_n185), .IN2(r847_n186), .QN(r847_n179) );
  NAND2X0 r847_U182 ( .IN1(P2_N5088), .IN2(r847_n184), .QN(r847_n180) );
  OR2X1 r847_U181 ( .IN2(P2_N5088), .IN1(r847_n184), .Q(r847_n182) );
  NAND2X0 r847_U180 ( .IN1(r847_n182), .IN2(r847_n183), .QN(r847_n181) );
  NAND2X0 r847_U179 ( .IN1(r847_n180), .IN2(r847_n181), .QN(r847_n174) );
  NAND2X0 r847_U178 ( .IN1(r847_n179), .IN2(r847_n174), .QN(r847_n177) );
  OR2X1 r847_U177 ( .IN2(r847_n174), .IN1(r847_n179), .Q(r847_n178) );
  NAND2X0 r847_U176 ( .IN1(r847_n177), .IN2(r847_n178), .QN(P2_N3148) );
  INVX0 r847_U175 ( .ZN(r847_n155), .INP(P2_N2997) );
  NAND2X0 r847_U174 ( .IN1(P2_N5090), .IN2(r847_n155), .QN(r847_n175) );
  OR2X1 r847_U173 ( .IN2(P2_N5090), .IN1(r847_n155), .Q(r847_n176) );
  NAND2X0 r847_U172 ( .IN1(r847_n175), .IN2(r847_n176), .QN(r847_n169) );
  NAND2X0 r847_U171 ( .IN1(n7187), .IN2(r847_n174), .QN(r847_n170) );
  OR2X1 r847_U170 ( .IN2(n7187), .IN1(r847_n174), .Q(r847_n172) );
  NAND2X0 r847_U169 ( .IN1(r847_n172), .IN2(r847_n173), .QN(r847_n171) );
  NAND2X0 r847_U168 ( .IN1(r847_n170), .IN2(r847_n171), .QN(r847_n156) );
  NAND2X0 r847_U167 ( .IN1(r847_n169), .IN2(r847_n156), .QN(r847_n167) );
  OR2X1 r847_U166 ( .IN2(r847_n156), .IN1(r847_n169), .Q(r847_n168) );
  NAND2X0 r847_U165 ( .IN1(r847_n167), .IN2(r847_n168), .QN(P2_N3149) );
  NAND2X0 r847_U164 ( .IN1(P2_N5072), .IN2(r847_n166), .QN(r847_n163) );
  NAND2X0 r847_U163 ( .IN1(P2_N2979), .IN2(n7184), .QN(r847_n164) );
  INVX0 r847_U321 ( .ZN(r847_n291), .INP(P2_N2978) );
  NOR2X0 r847_U320 ( .QN(r847_n287), .IN1(r847_n291), .IN2(n7035) );
  INVX0 r847_U319 ( .ZN(r847_n162), .INP(r847_n287) );
  NAND2X0 r847_U318 ( .IN1(n7035), .IN2(r847_n291), .QN(r847_n290) );
  NAND2X0 r847_U317 ( .IN1(r847_n162), .IN2(r847_n290), .QN(P2_N3130) );
  INVX0 r847_U316 ( .ZN(r847_n253), .INP(P2_N2988) );
  NAND2X0 r847_U315 ( .IN1(n7220), .IN2(r847_n253), .QN(r847_n288) );
  OR2X1 r847_U314 ( .IN2(n7220), .IN1(r847_n253), .Q(r847_n289) );
  NAND2X0 r847_U313 ( .IN1(r847_n288), .IN2(r847_n289), .QN(r847_n259) );
  NAND2X0 r847_U312 ( .IN1(P2_N5072), .IN2(r847_n162), .QN(r847_n284) );
  NAND2X0 r847_U310 ( .IN1(r847_n287), .IN2(n7184), .QN(r847_n286) );
  INVX0 r847_U309 ( .ZN(r847_n166), .INP(P2_N2979) );
  NAND2X0 r847_U308 ( .IN1(r847_n286), .IN2(r847_n166), .QN(r847_n285) );
  NAND2X0 r847_U307 ( .IN1(r847_n284), .IN2(r847_n285), .QN(r847_n53) );
  NAND2X0 r847_U306 ( .IN1(n7181), .IN2(r847_n53), .QN(r847_n281) );
  OR2X1 r847_U305 ( .IN2(n7181), .IN1(r847_n53), .Q(r847_n283) );
  INVX0 r847_U304 ( .ZN(r847_n56), .INP(P2_N2980) );
  NAND2X0 r847_U303 ( .IN1(r847_n283), .IN2(r847_n56), .QN(r847_n282) );
  NAND2X0 r847_U302 ( .IN1(r847_n281), .IN2(r847_n282), .QN(r847_n46) );
  NAND2X0 r847_U301 ( .IN1(P2_N5074), .IN2(r847_n46), .QN(r847_n278) );
  OR2X1 r847_U300 ( .IN2(P2_N5074), .IN1(r847_n46), .Q(r847_n280) );
  INVX0 r847_U299 ( .ZN(r847_n49), .INP(P2_N2981) );
  NAND2X0 r847_U298 ( .IN1(r847_n280), .IN2(r847_n49), .QN(r847_n279) );
  NAND2X0 r847_U297 ( .IN1(r847_n278), .IN2(r847_n279), .QN(r847_n39) );
  NAND2X0 r847_U296 ( .IN1(P2_N5075), .IN2(r847_n39), .QN(r847_n275) );
  OR2X1 r847_U295 ( .IN2(P2_N5075), .IN1(r847_n39), .Q(r847_n277) );
  INVX0 r847_U294 ( .ZN(r847_n42), .INP(P2_N2982) );
  NAND2X0 r847_U293 ( .IN1(r847_n277), .IN2(r847_n42), .QN(r847_n276) );
  NAND2X0 r847_U292 ( .IN1(r847_n275), .IN2(r847_n276), .QN(r847_n32) );
  NAND2X0 r847_U291 ( .IN1(n7165), .IN2(r847_n32), .QN(r847_n272) );
  OR2X1 r847_U290 ( .IN2(n7165), .IN1(r847_n32), .Q(r847_n274) );
  INVX0 r847_U289 ( .ZN(r847_n35), .INP(P2_N2983) );
  NAND2X0 r847_U288 ( .IN1(r847_n274), .IN2(r847_n35), .QN(r847_n273) );
  NAND2X0 r847_U287 ( .IN1(r847_n272), .IN2(r847_n273), .QN(r847_n25) );
  NAND2X0 r847_U286 ( .IN1(n7162), .IN2(r847_n25), .QN(r847_n269) );
  OR2X1 r847_U285 ( .IN2(n7162), .IN1(r847_n25), .Q(r847_n271) );
  INVX0 r847_U284 ( .ZN(r847_n28), .INP(P2_N2984) );
  NAND2X0 r847_U283 ( .IN1(r847_n271), .IN2(r847_n28), .QN(r847_n270) );
  NAND2X0 r847_U282 ( .IN1(r847_n269), .IN2(r847_n270), .QN(r847_n18) );
  NAND2X0 r847_U281 ( .IN1(n7158), .IN2(r847_n18), .QN(r847_n266) );
  OR2X1 r847_U280 ( .IN2(n7158), .IN1(r847_n18), .Q(r847_n268) );
  INVX0 r847_U279 ( .ZN(r847_n21), .INP(P2_N2985) );
  NAND2X0 r847_U278 ( .IN1(r847_n268), .IN2(r847_n21), .QN(r847_n267) );
  NAND2X0 r847_U277 ( .IN1(r847_n266), .IN2(r847_n267), .QN(r847_n11) );
  NAND2X0 r847_U276 ( .IN1(P2_N5079), .IN2(r847_n11), .QN(r847_n263) );
  OR2X1 r847_U275 ( .IN2(P2_N5079), .IN1(r847_n11), .Q(r847_n265) );
  INVX0 r847_U274 ( .ZN(r847_n14), .INP(P2_N2986) );
  NAND2X0 r847_U273 ( .IN1(r847_n265), .IN2(r847_n14), .QN(r847_n264) );
  NAND2X0 r847_U272 ( .IN1(r847_n263), .IN2(r847_n264), .QN(r847_n4) );
  NAND2X0 r847_U271 ( .IN1(n7151), .IN2(r847_n4), .QN(r847_n260) );
  OR2X1 r847_U270 ( .IN2(n7151), .IN1(r847_n4), .Q(r847_n262) );
  INVX0 r847_U269 ( .ZN(r847_n7), .INP(P2_N2987) );
  NAND2X0 r847_U268 ( .IN1(r847_n262), .IN2(r847_n7), .QN(r847_n261) );
  NAND2X0 r847_U267 ( .IN1(r847_n260), .IN2(r847_n261), .QN(r847_n254) );
  NAND2X0 r847_U266 ( .IN1(r847_n259), .IN2(r847_n254), .QN(r847_n257) );
  OR2X1 r847_U265 ( .IN2(r847_n254), .IN1(r847_n259), .Q(r847_n258) );
  NAND2X0 r847_U264 ( .IN1(r847_n257), .IN2(r847_n258), .QN(P2_N3140) );
  INVX0 r847_U263 ( .ZN(r847_n243), .INP(P2_N2989) );
  NAND2X0 r847_U262 ( .IN1(P2_N5082), .IN2(r847_n243), .QN(r847_n255) );
  OR2X1 r847_U261 ( .IN2(P2_N5082), .IN1(r847_n243), .Q(r847_n256) );
  NAND2X0 r847_U260 ( .IN1(r847_n255), .IN2(r847_n256), .QN(r847_n249) );
  NAND2X0 r847_U259 ( .IN1(n7220), .IN2(r847_n254), .QN(r847_n250) );
  OR2X1 r847_U258 ( .IN2(n7220), .IN1(r847_n254), .Q(r847_n252) );
  NAND2X0 r847_U257 ( .IN1(r847_n252), .IN2(r847_n253), .QN(r847_n251) );
  NAND2X0 r847_U256 ( .IN1(r847_n250), .IN2(r847_n251), .QN(r847_n244) );
  NOR2X0 r849_U17 ( .QN(r849_n15), .IN1(r849_n17), .IN2(r849_n18) );
  AND2X1 r849_U16 ( .IN1(r849_n17), .IN2(r849_n18), .Q(r849_n16) );
  NOR2X0 r849_U15 ( .QN(P2_N3510), .IN1(r849_n15), .IN2(r849_n16) );
  OR2X1 r849_U13 ( .IN2(P2_N3359), .IN1(n7153), .Q(r849_n12) );
  NAND2X0 r849_U12 ( .IN1(P2_N3359), .IN2(n7153), .QN(r849_n13) );
  NAND2X0 r849_U11 ( .IN1(r849_n12), .IN2(r849_n13), .QN(r849_n11) );
  NOR2X0 r849_U10 ( .QN(r849_n8), .IN1(r849_n10), .IN2(r849_n11) );
  AND2X1 r849_U9 ( .IN1(r849_n10), .IN2(r849_n11), .Q(r849_n9) );
  NOR2X0 r849_U8 ( .QN(P2_N3511), .IN1(r849_n8), .IN2(r849_n9) );
  OR2X1 r849_U6 ( .IN2(P2_N3360), .IN1(n7149), .Q(r849_n5) );
  NAND2X0 r849_U5 ( .IN1(P2_N3360), .IN2(n7149), .QN(r849_n6) );
  NAND2X0 r849_U4 ( .IN1(r849_n5), .IN2(r849_n6), .QN(r849_n4) );
  NOR2X0 r849_U3 ( .QN(r849_n1), .IN1(r849_n3), .IN2(r849_n4) );
  AND2X1 r849_U2 ( .IN1(r849_n3), .IN2(r849_n4), .Q(r849_n2) );
  NOR2X0 r849_U1 ( .QN(P2_N3512), .IN1(r849_n1), .IN2(r849_n2) );
  OR2X1 r849_U110 ( .IN2(n7238), .IN1(r849_n107), .Q(r849_n106) );
  NAND2X0 r849_U109 ( .IN1(P2_N3375), .IN2(r849_n106), .QN(r849_n105) );
  NAND2X0 r849_U108 ( .IN1(r849_n104), .IN2(r849_n105), .QN(r849_n97) );
  OR2X1 r849_U106 ( .IN2(P2_N3376), .IN1(n7234), .Q(r849_n101) );
  NAND2X0 r849_U105 ( .IN1(P2_N3376), .IN2(n7234), .QN(r849_n102) );
  NAND2X0 r849_U104 ( .IN1(r849_n101), .IN2(r849_n102), .QN(r849_n100) );
  NOR2X0 r849_U103 ( .QN(r849_n98), .IN1(r849_n97), .IN2(r849_n100) );
  AND2X1 r849_U102 ( .IN1(r849_n97), .IN2(r849_n100), .Q(r849_n99) );
  NOR2X0 r849_U101 ( .QN(P2_N3528), .IN1(r849_n98), .IN2(r849_n99) );
  NAND2X0 r849_U100 ( .IN1(n7237), .IN2(r849_n97), .QN(r849_n94) );
  OR2X1 r849_U99 ( .IN2(n7237), .IN1(r849_n97), .Q(r849_n96) );
  NAND2X0 r849_U98 ( .IN1(P2_N3376), .IN2(r849_n96), .QN(r849_n95) );
  NAND2X0 r849_U97 ( .IN1(r849_n94), .IN2(r849_n95), .QN(r849_n87) );
  OR2X1 r849_U95 ( .IN2(P2_N3377), .IN1(n7229), .Q(r849_n91) );
  NAND2X0 r849_U94 ( .IN1(P2_N3377), .IN2(n7229), .QN(r849_n92) );
  NAND2X0 r849_U93 ( .IN1(r849_n91), .IN2(r849_n92), .QN(r849_n90) );
  NOR2X0 r849_U92 ( .QN(r849_n88), .IN1(r849_n87), .IN2(r849_n90) );
  AND2X1 r849_U91 ( .IN1(r849_n87), .IN2(r849_n90), .Q(r849_n89) );
  NOR2X0 r849_U90 ( .QN(P2_N3529), .IN1(r849_n88), .IN2(r849_n89) );
  NAND2X0 r849_U89 ( .IN1(P2_N5097), .IN2(r849_n87), .QN(r849_n84) );
  OR2X1 r849_U88 ( .IN2(P2_N5097), .IN1(r849_n87), .Q(r849_n86) );
  NAND2X0 r849_U87 ( .IN1(P2_N3377), .IN2(r849_n86), .QN(r849_n85) );
  NAND2X0 r849_U86 ( .IN1(r849_n84), .IN2(r849_n85), .QN(r849_n77) );
  OR2X1 r849_U84 ( .IN2(P2_N3378), .IN1(n7224), .Q(r849_n81) );
  NAND2X0 r849_U83 ( .IN1(P2_N3378), .IN2(n7224), .QN(r849_n82) );
  NAND2X0 r849_U82 ( .IN1(r849_n81), .IN2(r849_n82), .QN(r849_n80) );
  NOR2X0 r849_U81 ( .QN(r849_n78), .IN1(r849_n77), .IN2(r849_n80) );
  AND2X1 r849_U80 ( .IN1(r849_n77), .IN2(r849_n80), .Q(r849_n79) );
  NOR2X0 r849_U79 ( .QN(P2_N3530), .IN1(r849_n78), .IN2(r849_n79) );
  NAND2X0 r849_U78 ( .IN1(P2_N5098), .IN2(r849_n77), .QN(r849_n74) );
  OR2X1 r849_U77 ( .IN2(P2_N5098), .IN1(r849_n77), .Q(r849_n76) );
  NAND2X0 r849_U76 ( .IN1(P2_N3378), .IN2(r849_n76), .QN(r849_n75) );
  NAND2X0 r849_U75 ( .IN1(r849_n74), .IN2(r849_n75), .QN(r849_n64) );
  OR2X1 r849_U73 ( .IN2(P2_N3379), .IN1(n7222), .Q(r849_n71) );
  NAND2X0 r849_U72 ( .IN1(P2_N3379), .IN2(n7222), .QN(r849_n72) );
  NAND2X0 r849_U71 ( .IN1(r849_n71), .IN2(r849_n72), .QN(r849_n70) );
  NOR2X0 r849_U70 ( .QN(r849_n68), .IN1(r849_n64), .IN2(r849_n70) );
  AND2X1 r849_U69 ( .IN1(r849_n64), .IN2(r849_n70), .Q(r849_n69) );
  NOR2X0 r849_U68 ( .QN(P2_N3531), .IN1(r849_n68), .IN2(r849_n69) );
  OR2X1 r849_U66 ( .IN2(P2_N3380), .IN1(n7266), .Q(r849_n65) );
  NAND2X0 r849_U65 ( .IN1(P2_N3380), .IN2(n7266), .QN(r849_n66) );
  NAND2X0 r849_U64 ( .IN1(r849_n65), .IN2(r849_n66), .QN(r849_n60) );
  NAND2X0 r849_U63 ( .IN1(P2_N5099), .IN2(r849_n64), .QN(r849_n61) );
  OR2X1 r849_U62 ( .IN2(P2_N5099), .IN1(r849_n64), .Q(r849_n63) );
  NAND2X0 r849_U61 ( .IN1(P2_N3379), .IN2(r849_n63), .QN(r849_n62) );
  NAND2X0 r849_U60 ( .IN1(r849_n61), .IN2(r849_n62), .QN(r849_n59) );
  NOR2X0 r849_U59 ( .QN(r849_n57), .IN1(r849_n60), .IN2(r849_n59) );
  AND2X1 r849_U58 ( .IN1(r849_n59), .IN2(r849_n60), .Q(r849_n58) );
  NOR2X0 r849_U57 ( .QN(P2_N3532), .IN1(r849_n57), .IN2(r849_n58) );
  OR2X1 r849_U55 ( .IN2(P2_N3353), .IN1(n7182), .Q(r849_n54) );
  NAND2X0 r849_U54 ( .IN1(P2_N3353), .IN2(n7182), .QN(r849_n55) );
  NAND2X0 r849_U53 ( .IN1(r849_n54), .IN2(r849_n55), .QN(r849_n53) );
  NOR2X0 r849_U52 ( .QN(r849_n50), .IN1(r849_n52), .IN2(r849_n53) );
  AND2X1 r849_U51 ( .IN1(r849_n52), .IN2(r849_n53), .Q(r849_n51) );
  NOR2X0 r849_U50 ( .QN(P2_N3505), .IN1(r849_n50), .IN2(r849_n51) );
  OR2X1 r849_U48 ( .IN2(P2_N3354), .IN1(n7178), .Q(r849_n47) );
  NAND2X0 r849_U47 ( .IN1(P2_N3354), .IN2(n7178), .QN(r849_n48) );
  NAND2X0 r849_U46 ( .IN1(r849_n47), .IN2(r849_n48), .QN(r849_n46) );
  NOR2X0 r849_U45 ( .QN(r849_n43), .IN1(r849_n45), .IN2(r849_n46) );
  AND2X1 r849_U44 ( .IN1(r849_n45), .IN2(r849_n46), .Q(r849_n44) );
  NOR2X0 r849_U43 ( .QN(P2_N3506), .IN1(r849_n43), .IN2(r849_n44) );
  OR2X1 r849_U41 ( .IN2(P2_N3355), .IN1(n7174), .Q(r849_n40) );
  NAND2X0 r849_U40 ( .IN1(P2_N3355), .IN2(n7174), .QN(r849_n41) );
  NAND2X0 r849_U39 ( .IN1(r849_n40), .IN2(r849_n41), .QN(r849_n39) );
  NOR2X0 r849_U38 ( .QN(r849_n36), .IN1(r849_n38), .IN2(r849_n39) );
  AND2X1 r849_U37 ( .IN1(r849_n38), .IN2(r849_n39), .Q(r849_n37) );
  NOR2X0 r849_U36 ( .QN(P2_N3507), .IN1(r849_n36), .IN2(r849_n37) );
  OR2X1 r849_U34 ( .IN2(P2_N3356), .IN1(n7166), .Q(r849_n33) );
  NAND2X0 r849_U33 ( .IN1(P2_N3356), .IN2(n7166), .QN(r849_n34) );
  NAND2X0 r849_U32 ( .IN1(r849_n33), .IN2(r849_n34), .QN(r849_n32) );
  NOR2X0 r849_U31 ( .QN(r849_n29), .IN1(r849_n31), .IN2(r849_n32) );
  AND2X1 r849_U30 ( .IN1(r849_n31), .IN2(r849_n32), .Q(r849_n30) );
  NOR2X0 r849_U29 ( .QN(P2_N3508), .IN1(r849_n29), .IN2(r849_n30) );
  OR2X1 r849_U27 ( .IN2(P2_N3357), .IN1(n7164), .Q(r849_n26) );
  NAND2X0 r849_U26 ( .IN1(P2_N3357), .IN2(n7164), .QN(r849_n27) );
  NAND2X0 r849_U25 ( .IN1(r849_n26), .IN2(r849_n27), .QN(r849_n25) );
  NOR2X0 r849_U24 ( .QN(r849_n22), .IN1(r849_n24), .IN2(r849_n25) );
  AND2X1 r849_U23 ( .IN1(r849_n24), .IN2(r849_n25), .Q(r849_n23) );
  NOR2X0 r849_U22 ( .QN(P2_N3509), .IN1(r849_n22), .IN2(r849_n23) );
  OR2X1 r849_U20 ( .IN2(P2_N3358), .IN1(n7157), .Q(r849_n19) );
  NAND2X0 r849_U19 ( .IN1(P2_N3358), .IN2(n7157), .QN(r849_n20) );
  NAND2X0 r849_U18 ( .IN1(r849_n19), .IN2(r849_n20), .QN(r849_n18) );
  NAND2X0 r849_U203 ( .IN1(P2_N3367), .IN2(r849_n193), .QN(r849_n192) );
  NAND2X0 r849_U202 ( .IN1(r849_n191), .IN2(r849_n192), .QN(r849_n184) );
  OR2X1 r849_U200 ( .IN2(P2_N3368), .IN1(n7195), .Q(r849_n188) );
  NAND2X0 r849_U199 ( .IN1(P2_N3368), .IN2(n7195), .QN(r849_n189) );
  NAND2X0 r849_U198 ( .IN1(r849_n188), .IN2(r849_n189), .QN(r849_n187) );
  NOR2X0 r849_U197 ( .QN(r849_n185), .IN1(r849_n184), .IN2(r849_n187) );
  AND2X1 r849_U196 ( .IN1(r849_n184), .IN2(r849_n187), .Q(r849_n186) );
  NOR2X0 r849_U195 ( .QN(P2_N3520), .IN1(r849_n185), .IN2(r849_n186) );
  NAND2X0 r849_U194 ( .IN1(n7194), .IN2(r849_n184), .QN(r849_n181) );
  OR2X1 r849_U193 ( .IN2(n7194), .IN1(r849_n184), .Q(r849_n183) );
  NAND2X0 r849_U192 ( .IN1(P2_N3368), .IN2(r849_n183), .QN(r849_n182) );
  NAND2X0 r849_U191 ( .IN1(r849_n181), .IN2(r849_n182), .QN(r849_n174) );
  OR2X1 r849_U189 ( .IN2(P2_N3369), .IN1(n7188), .Q(r849_n178) );
  NAND2X0 r849_U188 ( .IN1(P2_N3369), .IN2(n7188), .QN(r849_n179) );
  NAND2X0 r849_U187 ( .IN1(r849_n178), .IN2(r849_n179), .QN(r849_n177) );
  NOR2X0 r849_U186 ( .QN(r849_n175), .IN1(r849_n174), .IN2(r849_n177) );
  AND2X1 r849_U185 ( .IN1(r849_n174), .IN2(r849_n177), .Q(r849_n176) );
  NOR2X0 r849_U184 ( .QN(P2_N3521), .IN1(r849_n175), .IN2(r849_n176) );
  NAND2X0 r849_U183 ( .IN1(P2_N5089), .IN2(r849_n174), .QN(r849_n171) );
  OR2X1 r849_U182 ( .IN2(P2_N5089), .IN1(r849_n174), .Q(r849_n173) );
  NAND2X0 r849_U181 ( .IN1(P2_N3369), .IN2(r849_n173), .QN(r849_n172) );
  NAND2X0 r849_U180 ( .IN1(r849_n171), .IN2(r849_n172), .QN(r849_n157) );
  OR2X1 r849_U178 ( .IN2(P2_N3370), .IN1(n7264), .Q(r849_n168) );
  NAND2X0 r849_U177 ( .IN1(P2_N3370), .IN2(n7264), .QN(r849_n169) );
  NAND2X0 r849_U176 ( .IN1(r849_n168), .IN2(r849_n169), .QN(r849_n167) );
  NOR2X0 r849_U175 ( .QN(r849_n165), .IN1(r849_n157), .IN2(r849_n167) );
  AND2X1 r849_U174 ( .IN1(r849_n157), .IN2(r849_n167), .Q(r849_n166) );
  NOR2X0 r849_U173 ( .QN(P2_N3522), .IN1(r849_n165), .IN2(r849_n166) );
  OR2X1 r849_U172 ( .IN2(P2_N3352), .IN1(n7184), .Q(r849_n162) );
  NAND2X0 r849_U171 ( .IN1(P2_N3352), .IN2(n7184), .QN(r849_n163) );
  NAND2X0 r849_U170 ( .IN1(r849_n162), .IN2(r849_n163), .QN(r849_n160) );
  NAND2X0 r849_U169 ( .IN1(r849_n160), .IN2(r849_n161), .QN(r849_n158) );
  OR2X1 r849_U168 ( .IN2(r849_n161), .IN1(r849_n160), .Q(r849_n159) );
  NAND2X0 r849_U167 ( .IN1(r849_n158), .IN2(r849_n159), .QN(P2_N3504) );
  NAND2X0 r849_U166 ( .IN1(P2_N5090), .IN2(r849_n157), .QN(r849_n154) );
  OR2X1 r849_U165 ( .IN2(P2_N5090), .IN1(r849_n157), .Q(r849_n156) );
  NAND2X0 r849_U164 ( .IN1(P2_N3370), .IN2(r849_n156), .QN(r849_n155) );
  NAND2X0 r849_U163 ( .IN1(r849_n154), .IN2(r849_n155), .QN(r849_n147) );
  OR2X1 r849_U161 ( .IN2(P2_N3371), .IN1(n7260), .Q(r849_n151) );
  NAND2X0 r849_U160 ( .IN1(P2_N3371), .IN2(n7260), .QN(r849_n152) );
  NAND2X0 r849_U159 ( .IN1(r849_n151), .IN2(r849_n152), .QN(r849_n150) );
  NOR2X0 r849_U158 ( .QN(r849_n148), .IN1(r849_n147), .IN2(r849_n150) );
  AND2X1 r849_U157 ( .IN1(r849_n147), .IN2(r849_n150), .Q(r849_n149) );
  NOR2X0 r849_U156 ( .QN(P2_N3523), .IN1(r849_n148), .IN2(r849_n149) );
  NAND2X0 r849_U155 ( .IN1(P2_N5091), .IN2(r849_n147), .QN(r849_n144) );
  OR2X1 r849_U154 ( .IN2(P2_N5091), .IN1(r849_n147), .Q(r849_n146) );
  NAND2X0 r849_U153 ( .IN1(P2_N3371), .IN2(r849_n146), .QN(r849_n145) );
  NAND2X0 r849_U152 ( .IN1(r849_n144), .IN2(r849_n145), .QN(r849_n137) );
  OR2X1 r849_U150 ( .IN2(P2_N3372), .IN1(n7253), .Q(r849_n141) );
  NAND2X0 r849_U149 ( .IN1(P2_N3372), .IN2(n7253), .QN(r849_n142) );
  NAND2X0 r849_U148 ( .IN1(r849_n141), .IN2(r849_n142), .QN(r849_n140) );
  NOR2X0 r849_U147 ( .QN(r849_n138), .IN1(r849_n137), .IN2(r849_n140) );
  AND2X1 r849_U146 ( .IN1(r849_n137), .IN2(r849_n140), .Q(r849_n139) );
  NOR2X0 r849_U145 ( .QN(P2_N3524), .IN1(r849_n138), .IN2(r849_n139) );
  NAND2X0 r849_U144 ( .IN1(n7252), .IN2(r849_n137), .QN(r849_n134) );
  OR2X1 r849_U143 ( .IN2(n7252), .IN1(r849_n137), .Q(r849_n136) );
  NAND2X0 r849_U142 ( .IN1(P2_N3372), .IN2(r849_n136), .QN(r849_n135) );
  NAND2X0 r849_U141 ( .IN1(r849_n134), .IN2(r849_n135), .QN(r849_n127) );
  OR2X1 r849_U139 ( .IN2(P2_N3373), .IN1(n7248), .Q(r849_n131) );
  NAND2X0 r849_U138 ( .IN1(P2_N3373), .IN2(n7248), .QN(r849_n132) );
  NAND2X0 r849_U137 ( .IN1(r849_n131), .IN2(r849_n132), .QN(r849_n130) );
  NOR2X0 r849_U136 ( .QN(r849_n128), .IN1(r849_n127), .IN2(r849_n130) );
  AND2X1 r849_U135 ( .IN1(r849_n127), .IN2(r849_n130), .Q(r849_n129) );
  NOR2X0 r849_U134 ( .QN(P2_N3525), .IN1(r849_n128), .IN2(r849_n129) );
  NAND2X0 r849_U133 ( .IN1(n7247), .IN2(r849_n127), .QN(r849_n124) );
  OR2X1 r849_U132 ( .IN2(n7247), .IN1(r849_n127), .Q(r849_n126) );
  NAND2X0 r849_U131 ( .IN1(P2_N3373), .IN2(r849_n126), .QN(r849_n125) );
  NAND2X0 r849_U130 ( .IN1(r849_n124), .IN2(r849_n125), .QN(r849_n117) );
  OR2X1 r849_U128 ( .IN2(P2_N3374), .IN1(n7243), .Q(r849_n121) );
  NAND2X0 r849_U127 ( .IN1(P2_N3374), .IN2(n7243), .QN(r849_n122) );
  NAND2X0 r849_U126 ( .IN1(r849_n121), .IN2(r849_n122), .QN(r849_n120) );
  NOR2X0 r849_U125 ( .QN(r849_n118), .IN1(r849_n117), .IN2(r849_n120) );
  AND2X1 r849_U124 ( .IN1(r849_n117), .IN2(r849_n120), .Q(r849_n119) );
  NOR2X0 r849_U123 ( .QN(P2_N3526), .IN1(r849_n118), .IN2(r849_n119) );
  NAND2X0 r849_U122 ( .IN1(n7242), .IN2(r849_n117), .QN(r849_n114) );
  OR2X1 r849_U121 ( .IN2(n7242), .IN1(r849_n117), .Q(r849_n116) );
  NAND2X0 r849_U120 ( .IN1(P2_N3374), .IN2(r849_n116), .QN(r849_n115) );
  NAND2X0 r849_U119 ( .IN1(r849_n114), .IN2(r849_n115), .QN(r849_n107) );
  OR2X1 r849_U117 ( .IN2(P2_N3375), .IN1(n7239), .Q(r849_n111) );
  NAND2X0 r849_U116 ( .IN1(P2_N3375), .IN2(n7239), .QN(r849_n112) );
  NAND2X0 r849_U115 ( .IN1(r849_n111), .IN2(r849_n112), .QN(r849_n110) );
  NOR2X0 r849_U114 ( .QN(r849_n108), .IN1(r849_n107), .IN2(r849_n110) );
  AND2X1 r849_U113 ( .IN1(r849_n107), .IN2(r849_n110), .Q(r849_n109) );
  NOR2X0 r849_U112 ( .QN(P2_N3527), .IN1(r849_n108), .IN2(r849_n109) );
  NAND2X0 r849_U111 ( .IN1(n7238), .IN2(r849_n107), .QN(r849_n104) );
  NAND2X0 r849_U296 ( .IN1(P2_N3356), .IN2(r849_n275), .QN(r849_n274) );
  NAND2X0 r849_U295 ( .IN1(r849_n273), .IN2(r849_n274), .QN(r849_n24) );
  NAND2X0 r849_U294 ( .IN1(n7162), .IN2(r849_n24), .QN(r849_n270) );
  OR2X1 r849_U293 ( .IN2(n7162), .IN1(r849_n24), .Q(r849_n272) );
  NAND2X0 r849_U292 ( .IN1(P2_N3357), .IN2(r849_n272), .QN(r849_n271) );
  NAND2X0 r849_U291 ( .IN1(r849_n270), .IN2(r849_n271), .QN(r849_n17) );
  NAND2X0 r849_U290 ( .IN1(P2_N5078), .IN2(r849_n17), .QN(r849_n267) );
  OR2X1 r849_U289 ( .IN2(P2_N5078), .IN1(r849_n17), .Q(r849_n269) );
  NAND2X0 r849_U288 ( .IN1(P2_N3358), .IN2(r849_n269), .QN(r849_n268) );
  NAND2X0 r849_U287 ( .IN1(r849_n267), .IN2(r849_n268), .QN(r849_n10) );
  NAND2X0 r849_U286 ( .IN1(P2_N5079), .IN2(r849_n10), .QN(r849_n264) );
  OR2X1 r849_U285 ( .IN2(P2_N5079), .IN1(r849_n10), .Q(r849_n266) );
  NAND2X0 r849_U284 ( .IN1(P2_N3359), .IN2(r849_n266), .QN(r849_n265) );
  NAND2X0 r849_U283 ( .IN1(r849_n264), .IN2(r849_n265), .QN(r849_n3) );
  NAND2X0 r849_U282 ( .IN1(P2_N5080), .IN2(r849_n3), .QN(r849_n261) );
  OR2X1 r849_U281 ( .IN2(P2_N5080), .IN1(r849_n3), .Q(r849_n263) );
  NAND2X0 r849_U280 ( .IN1(P2_N3360), .IN2(r849_n263), .QN(r849_n262) );
  NAND2X0 r849_U279 ( .IN1(r849_n261), .IN2(r849_n262), .QN(r849_n254) );
  OR2X1 r849_U277 ( .IN2(P2_N3361), .IN1(n7219), .Q(r849_n258) );
  NAND2X0 r849_U276 ( .IN1(P2_N3361), .IN2(n7219), .QN(r849_n259) );
  NAND2X0 r849_U275 ( .IN1(r849_n258), .IN2(r849_n259), .QN(r849_n257) );
  NOR2X0 r849_U274 ( .QN(r849_n255), .IN1(r849_n254), .IN2(r849_n257) );
  AND2X1 r849_U273 ( .IN1(r849_n254), .IN2(r849_n257), .Q(r849_n256) );
  NOR2X0 r849_U272 ( .QN(P2_N3513), .IN1(r849_n255), .IN2(r849_n256) );
  NAND2X0 r849_U271 ( .IN1(n7220), .IN2(r849_n254), .QN(r849_n251) );
  OR2X1 r849_U270 ( .IN2(n7220), .IN1(r849_n254), .Q(r849_n253) );
  NAND2X0 r849_U269 ( .IN1(P2_N3361), .IN2(r849_n253), .QN(r849_n252) );
  NAND2X0 r849_U268 ( .IN1(r849_n251), .IN2(r849_n252), .QN(r849_n244) );
  OR2X1 r849_U266 ( .IN2(P2_N3362), .IN1(n7214), .Q(r849_n248) );
  NAND2X0 r849_U265 ( .IN1(P2_N3362), .IN2(n7214), .QN(r849_n249) );
  NAND2X0 r849_U264 ( .IN1(r849_n248), .IN2(r849_n249), .QN(r849_n247) );
  NOR2X0 r849_U263 ( .QN(r849_n245), .IN1(r849_n244), .IN2(r849_n247) );
  AND2X1 r849_U262 ( .IN1(r849_n244), .IN2(r849_n247), .Q(r849_n246) );
  NOR2X0 r849_U261 ( .QN(P2_N3514), .IN1(r849_n245), .IN2(r849_n246) );
  NAND2X0 r849_U260 ( .IN1(n7216), .IN2(r849_n244), .QN(r849_n241) );
  OR2X1 r849_U259 ( .IN2(n7216), .IN1(r849_n244), .Q(r849_n243) );
  NAND2X0 r849_U258 ( .IN1(P2_N3362), .IN2(r849_n243), .QN(r849_n242) );
  NAND2X0 r849_U257 ( .IN1(r849_n241), .IN2(r849_n242), .QN(r849_n234) );
  OR2X1 r849_U255 ( .IN2(P2_N3363), .IN1(n7211), .Q(r849_n238) );
  NAND2X0 r849_U254 ( .IN1(P2_N3363), .IN2(n7211), .QN(r849_n239) );
  NAND2X0 r849_U253 ( .IN1(r849_n238), .IN2(r849_n239), .QN(r849_n237) );
  NOR2X0 r849_U252 ( .QN(r849_n235), .IN1(r849_n234), .IN2(r849_n237) );
  AND2X1 r849_U251 ( .IN1(r849_n234), .IN2(r849_n237), .Q(r849_n236) );
  NOR2X0 r849_U250 ( .QN(P2_N3515), .IN1(r849_n235), .IN2(r849_n236) );
  NAND2X0 r849_U249 ( .IN1(n7210), .IN2(r849_n234), .QN(r849_n231) );
  OR2X1 r849_U248 ( .IN2(n7210), .IN1(r849_n234), .Q(r849_n233) );
  NAND2X0 r849_U247 ( .IN1(P2_N3363), .IN2(r849_n233), .QN(r849_n232) );
  NAND2X0 r849_U246 ( .IN1(r849_n231), .IN2(r849_n232), .QN(r849_n224) );
  OR2X1 r849_U244 ( .IN2(P2_N3364), .IN1(n7208), .Q(r849_n228) );
  NAND2X0 r849_U243 ( .IN1(P2_N3364), .IN2(n7208), .QN(r849_n229) );
  NAND2X0 r849_U242 ( .IN1(r849_n228), .IN2(r849_n229), .QN(r849_n227) );
  NOR2X0 r849_U241 ( .QN(r849_n225), .IN1(r849_n224), .IN2(r849_n227) );
  AND2X1 r849_U240 ( .IN1(r849_n224), .IN2(r849_n227), .Q(r849_n226) );
  NOR2X0 r849_U239 ( .QN(P2_N3516), .IN1(r849_n225), .IN2(r849_n226) );
  NAND2X0 r849_U238 ( .IN1(P2_N5084), .IN2(r849_n224), .QN(r849_n221) );
  OR2X1 r849_U237 ( .IN2(P2_N5084), .IN1(r849_n224), .Q(r849_n223) );
  NAND2X0 r849_U236 ( .IN1(P2_N3364), .IN2(r849_n223), .QN(r849_n222) );
  NAND2X0 r849_U235 ( .IN1(r849_n221), .IN2(r849_n222), .QN(r849_n214) );
  OR2X1 r849_U233 ( .IN2(P2_N3365), .IN1(n7205), .Q(r849_n218) );
  NAND2X0 r849_U232 ( .IN1(P2_N3365), .IN2(n7205), .QN(r849_n219) );
  NAND2X0 r849_U231 ( .IN1(r849_n218), .IN2(r849_n219), .QN(r849_n217) );
  NOR2X0 r849_U230 ( .QN(r849_n215), .IN1(r849_n214), .IN2(r849_n217) );
  AND2X1 r849_U229 ( .IN1(r849_n214), .IN2(r849_n217), .Q(r849_n216) );
  NOR2X0 r849_U228 ( .QN(P2_N3517), .IN1(r849_n215), .IN2(r849_n216) );
  NAND2X0 r849_U227 ( .IN1(P2_N5085), .IN2(r849_n214), .QN(r849_n211) );
  OR2X1 r849_U226 ( .IN2(P2_N5085), .IN1(r849_n214), .Q(r849_n213) );
  NAND2X0 r849_U225 ( .IN1(P2_N3365), .IN2(r849_n213), .QN(r849_n212) );
  NAND2X0 r849_U224 ( .IN1(r849_n211), .IN2(r849_n212), .QN(r849_n204) );
  OR2X1 r849_U222 ( .IN2(P2_N3366), .IN1(n7201), .Q(r849_n208) );
  NAND2X0 r849_U221 ( .IN1(P2_N3366), .IN2(n7201), .QN(r849_n209) );
  NAND2X0 r849_U220 ( .IN1(r849_n208), .IN2(r849_n209), .QN(r849_n207) );
  NOR2X0 r849_U219 ( .QN(r849_n205), .IN1(r849_n204), .IN2(r849_n207) );
  AND2X1 r849_U218 ( .IN1(r849_n204), .IN2(r849_n207), .Q(r849_n206) );
  NOR2X0 r849_U217 ( .QN(P2_N3518), .IN1(r849_n205), .IN2(r849_n206) );
  NAND2X0 r849_U216 ( .IN1(P2_N5086), .IN2(r849_n204), .QN(r849_n201) );
  OR2X1 r849_U215 ( .IN2(P2_N5086), .IN1(r849_n204), .Q(r849_n203) );
  NAND2X0 r849_U214 ( .IN1(P2_N3366), .IN2(r849_n203), .QN(r849_n202) );
  NAND2X0 r849_U213 ( .IN1(r849_n201), .IN2(r849_n202), .QN(r849_n194) );
  OR2X1 r849_U211 ( .IN2(P2_N3367), .IN1(n7197), .Q(r849_n198) );
  NAND2X0 r849_U210 ( .IN1(P2_N3367), .IN2(n7197), .QN(r849_n199) );
  NAND2X0 r849_U209 ( .IN1(r849_n198), .IN2(r849_n199), .QN(r849_n197) );
  NOR2X0 r849_U208 ( .QN(r849_n195), .IN1(r849_n194), .IN2(r849_n197) );
  AND2X1 r849_U207 ( .IN1(r849_n194), .IN2(r849_n197), .Q(r849_n196) );
  NOR2X0 r849_U206 ( .QN(P2_N3519), .IN1(r849_n195), .IN2(r849_n196) );
  NAND2X0 r849_U205 ( .IN1(P2_N5087), .IN2(r849_n194), .QN(r849_n191) );
  OR2X1 r849_U204 ( .IN2(P2_N5087), .IN1(r849_n194), .Q(r849_n193) );
  OR2X1 r849_U319 ( .IN2(P2_N3351), .IN1(n2919), .Q(r849_n288) );
  NAND2X0 r849_U318 ( .IN1(P2_N3351), .IN2(n2919), .QN(r849_n289) );
  NAND2X0 r849_U317 ( .IN1(r849_n288), .IN2(r849_n289), .QN(P2_N3503) );
  NAND2X0 r849_U315 ( .IN1(P2_N3351), .IN2(n7035), .QN(r849_n161) );
  OR2X1 r849_U314 ( .IN2(r849_n161), .IN1(n7184), .Q(r849_n285) );
  NAND2X0 r849_U313 ( .IN1(n7184), .IN2(r849_n161), .QN(r849_n287) );
  NAND2X0 r849_U312 ( .IN1(P2_N3352), .IN2(r849_n287), .QN(r849_n286) );
  NAND2X0 r849_U311 ( .IN1(r849_n285), .IN2(r849_n286), .QN(r849_n52) );
  NAND2X0 r849_U310 ( .IN1(n7181), .IN2(r849_n52), .QN(r849_n282) );
  OR2X1 r849_U309 ( .IN2(n7181), .IN1(r849_n52), .Q(r849_n284) );
  NAND2X0 r849_U308 ( .IN1(P2_N3353), .IN2(r849_n284), .QN(r849_n283) );
  NAND2X0 r849_U307 ( .IN1(r849_n282), .IN2(r849_n283), .QN(r849_n45) );
  NAND2X0 r849_U306 ( .IN1(n7177), .IN2(r849_n45), .QN(r849_n279) );
  OR2X1 r849_U305 ( .IN2(n7177), .IN1(r849_n45), .Q(r849_n281) );
  NAND2X0 r849_U304 ( .IN1(P2_N3354), .IN2(r849_n281), .QN(r849_n280) );
  NAND2X0 r849_U303 ( .IN1(r849_n279), .IN2(r849_n280), .QN(r849_n38) );
  NAND2X0 r849_U302 ( .IN1(n7173), .IN2(r849_n38), .QN(r849_n276) );
  OR2X1 r849_U301 ( .IN2(n7173), .IN1(r849_n38), .Q(r849_n278) );
  NAND2X0 r849_U300 ( .IN1(P2_N3355), .IN2(r849_n278), .QN(r849_n277) );
  NAND2X0 r849_U299 ( .IN1(r849_n276), .IN2(r849_n277), .QN(r849_n31) );
  NAND2X0 r849_U298 ( .IN1(n7165), .IN2(r849_n31), .QN(r849_n273) );
  OR2X1 r849_U297 ( .IN2(n7165), .IN1(r849_n31), .Q(r849_n275) );
  OR2X1 r851_U58 ( .IN2(P2_N3753), .IN1(n7266), .Q(r851_n66) );
  NAND2X0 r851_U57 ( .IN1(P2_N3753), .IN2(n7266), .QN(r851_n67) );
  NAND2X0 r851_U56 ( .IN1(r851_n66), .IN2(r851_n67), .QN(r851_n60) );
  NAND2X0 r851_U55 ( .IN1(P2_N5099), .IN2(r851_n65), .QN(r851_n61) );
  OR2X1 r851_U54 ( .IN2(P2_N5099), .IN1(r851_n65), .Q(r851_n63) );
  NAND2X0 r851_U53 ( .IN1(r851_n63), .IN2(r851_n64), .QN(r851_n62) );
  NAND2X0 r851_U52 ( .IN1(r851_n61), .IN2(r851_n62), .QN(r851_n59) );
  NAND2X0 r851_U51 ( .IN1(r851_n60), .IN2(r851_n59), .QN(r851_n57) );
  OR2X1 r851_U50 ( .IN2(r851_n60), .IN1(r851_n59), .Q(r851_n58) );
  NAND2X0 r851_U49 ( .IN1(r851_n57), .IN2(r851_n58), .QN(P2_N3905) );
  NAND2X0 r851_U48 ( .IN1(P2_N5073), .IN2(r851_n56), .QN(r851_n54) );
  OR2X1 r851_U47 ( .IN2(P2_N5073), .IN1(r851_n56), .Q(r851_n55) );
  NAND2X0 r851_U46 ( .IN1(r851_n54), .IN2(r851_n55), .QN(r851_n52) );
  NAND2X0 r851_U45 ( .IN1(r851_n52), .IN2(r851_n53), .QN(r851_n50) );
  OR2X1 r851_U44 ( .IN2(r851_n53), .IN1(r851_n52), .Q(r851_n51) );
  NAND2X0 r851_U43 ( .IN1(r851_n50), .IN2(r851_n51), .QN(P2_N3878) );
  NAND2X0 r851_U42 ( .IN1(n7177), .IN2(r851_n49), .QN(r851_n47) );
  OR2X1 r851_U41 ( .IN2(n7177), .IN1(r851_n49), .Q(r851_n48) );
  NAND2X0 r851_U40 ( .IN1(r851_n47), .IN2(r851_n48), .QN(r851_n45) );
  NAND2X0 r851_U39 ( .IN1(r851_n45), .IN2(r851_n46), .QN(r851_n43) );
  OR2X1 r851_U38 ( .IN2(r851_n46), .IN1(r851_n45), .Q(r851_n44) );
  NAND2X0 r851_U37 ( .IN1(r851_n43), .IN2(r851_n44), .QN(P2_N3879) );
  NAND2X0 r851_U36 ( .IN1(n7173), .IN2(r851_n42), .QN(r851_n40) );
  OR2X1 r851_U35 ( .IN2(n7173), .IN1(r851_n42), .Q(r851_n41) );
  NAND2X0 r851_U34 ( .IN1(r851_n40), .IN2(r851_n41), .QN(r851_n38) );
  NAND2X0 r851_U33 ( .IN1(r851_n38), .IN2(r851_n39), .QN(r851_n36) );
  OR2X1 r851_U32 ( .IN2(r851_n39), .IN1(r851_n38), .Q(r851_n37) );
  NAND2X0 r851_U31 ( .IN1(r851_n36), .IN2(r851_n37), .QN(P2_N3880) );
  NAND2X0 r851_U30 ( .IN1(P2_N5076), .IN2(r851_n35), .QN(r851_n33) );
  OR2X1 r851_U29 ( .IN2(P2_N5076), .IN1(r851_n35), .Q(r851_n34) );
  NAND2X0 r851_U28 ( .IN1(r851_n33), .IN2(r851_n34), .QN(r851_n31) );
  NAND2X0 r851_U27 ( .IN1(r851_n31), .IN2(r851_n32), .QN(r851_n29) );
  OR2X1 r851_U26 ( .IN2(r851_n32), .IN1(r851_n31), .Q(r851_n30) );
  NAND2X0 r851_U25 ( .IN1(r851_n29), .IN2(r851_n30), .QN(P2_N3881) );
  NAND2X0 r851_U24 ( .IN1(n7162), .IN2(r851_n28), .QN(r851_n26) );
  OR2X1 r851_U23 ( .IN2(n7162), .IN1(r851_n28), .Q(r851_n27) );
  NAND2X0 r851_U22 ( .IN1(r851_n26), .IN2(r851_n27), .QN(r851_n24) );
  NAND2X0 r851_U21 ( .IN1(r851_n24), .IN2(r851_n25), .QN(r851_n22) );
  OR2X1 r851_U20 ( .IN2(r851_n25), .IN1(r851_n24), .Q(r851_n23) );
  NAND2X0 r851_U19 ( .IN1(r851_n22), .IN2(r851_n23), .QN(P2_N3882) );
  NAND2X0 r851_U18 ( .IN1(P2_N5078), .IN2(r851_n21), .QN(r851_n19) );
  OR2X1 r851_U17 ( .IN2(P2_N5078), .IN1(r851_n21), .Q(r851_n20) );
  NAND2X0 r851_U16 ( .IN1(r851_n19), .IN2(r851_n20), .QN(r851_n17) );
  NAND2X0 r851_U15 ( .IN1(r851_n17), .IN2(r851_n18), .QN(r851_n15) );
  OR2X1 r851_U14 ( .IN2(r851_n18), .IN1(r851_n17), .Q(r851_n16) );
  NAND2X0 r851_U13 ( .IN1(r851_n15), .IN2(r851_n16), .QN(P2_N3883) );
  NAND2X0 r851_U12 ( .IN1(n7154), .IN2(r851_n14), .QN(r851_n12) );
  OR2X1 r851_U11 ( .IN2(n7154), .IN1(r851_n14), .Q(r851_n13) );
  NAND2X0 r851_U10 ( .IN1(r851_n12), .IN2(r851_n13), .QN(r851_n10) );
  NAND2X0 r851_U9 ( .IN1(r851_n10), .IN2(r851_n11), .QN(r851_n8) );
  OR2X1 r851_U8 ( .IN2(r851_n11), .IN1(r851_n10), .Q(r851_n9) );
  NAND2X0 r851_U7 ( .IN1(r851_n8), .IN2(r851_n9), .QN(P2_N3884) );
  NAND2X0 r851_U6 ( .IN1(n7151), .IN2(r851_n7), .QN(r851_n5) );
  OR2X1 r851_U5 ( .IN2(n7151), .IN1(r851_n7), .Q(r851_n6) );
  NAND2X0 r851_U4 ( .IN1(r851_n5), .IN2(r851_n6), .QN(r851_n3) );
  NAND2X0 r851_U3 ( .IN1(r851_n3), .IN2(r851_n4), .QN(r851_n1) );
  OR2X1 r851_U2 ( .IN2(r851_n4), .IN1(r851_n3), .Q(r851_n2) );
  NAND2X0 r851_U1 ( .IN1(r851_n1), .IN2(r851_n2), .QN(P2_N3885) );
  NAND2X0 r851_U152 ( .IN1(r851_n154), .IN2(r851_n155), .QN(r851_n153) );
  NAND2X0 r851_U151 ( .IN1(r851_n152), .IN2(r851_n153), .QN(r851_n146) );
  NAND2X0 r851_U150 ( .IN1(r851_n151), .IN2(r851_n146), .QN(r851_n149) );
  OR2X1 r851_U149 ( .IN2(r851_n146), .IN1(r851_n151), .Q(r851_n150) );
  NAND2X0 r851_U148 ( .IN1(r851_n149), .IN2(r851_n150), .QN(P2_N3896) );
  INVX0 r851_U147 ( .ZN(r851_n135), .INP(P2_N3745) );
  NAND2X0 r851_U146 ( .IN1(n7252), .IN2(r851_n135), .QN(r851_n147) );
  OR2X1 r851_U145 ( .IN2(n7252), .IN1(r851_n135), .Q(r851_n148) );
  NAND2X0 r851_U144 ( .IN1(r851_n147), .IN2(r851_n148), .QN(r851_n141) );
  NAND2X0 r851_U143 ( .IN1(P2_N5091), .IN2(r851_n146), .QN(r851_n142) );
  OR2X1 r851_U142 ( .IN2(P2_N5091), .IN1(r851_n146), .Q(r851_n144) );
  NAND2X0 r851_U141 ( .IN1(r851_n144), .IN2(r851_n145), .QN(r851_n143) );
  NAND2X0 r851_U140 ( .IN1(r851_n142), .IN2(r851_n143), .QN(r851_n136) );
  NAND2X0 r851_U139 ( .IN1(r851_n141), .IN2(r851_n136), .QN(r851_n139) );
  OR2X1 r851_U138 ( .IN2(r851_n136), .IN1(r851_n141), .Q(r851_n140) );
  NAND2X0 r851_U137 ( .IN1(r851_n139), .IN2(r851_n140), .QN(P2_N3897) );
  INVX0 r851_U136 ( .ZN(r851_n125), .INP(P2_N3746) );
  NAND2X0 r851_U135 ( .IN1(P2_N5093), .IN2(r851_n125), .QN(r851_n137) );
  OR2X1 r851_U134 ( .IN2(P2_N5093), .IN1(r851_n125), .Q(r851_n138) );
  NAND2X0 r851_U133 ( .IN1(r851_n137), .IN2(r851_n138), .QN(r851_n131) );
  NAND2X0 r851_U132 ( .IN1(n7252), .IN2(r851_n136), .QN(r851_n132) );
  OR2X1 r851_U131 ( .IN2(n7252), .IN1(r851_n136), .Q(r851_n134) );
  NAND2X0 r851_U130 ( .IN1(r851_n134), .IN2(r851_n135), .QN(r851_n133) );
  NAND2X0 r851_U129 ( .IN1(r851_n132), .IN2(r851_n133), .QN(r851_n126) );
  NAND2X0 r851_U128 ( .IN1(r851_n131), .IN2(r851_n126), .QN(r851_n129) );
  OR2X1 r851_U127 ( .IN2(r851_n126), .IN1(r851_n131), .Q(r851_n130) );
  NAND2X0 r851_U126 ( .IN1(r851_n129), .IN2(r851_n130), .QN(P2_N3898) );
  INVX0 r851_U125 ( .ZN(r851_n115), .INP(P2_N3747) );
  NAND2X0 r851_U124 ( .IN1(n7242), .IN2(r851_n115), .QN(r851_n127) );
  OR2X1 r851_U123 ( .IN2(n7242), .IN1(r851_n115), .Q(r851_n128) );
  NAND2X0 r851_U122 ( .IN1(r851_n127), .IN2(r851_n128), .QN(r851_n121) );
  NAND2X0 r851_U121 ( .IN1(P2_N5093), .IN2(r851_n126), .QN(r851_n122) );
  OR2X1 r851_U120 ( .IN2(P2_N5093), .IN1(r851_n126), .Q(r851_n124) );
  NAND2X0 r851_U119 ( .IN1(r851_n124), .IN2(r851_n125), .QN(r851_n123) );
  NAND2X0 r851_U118 ( .IN1(r851_n122), .IN2(r851_n123), .QN(r851_n116) );
  NAND2X0 r851_U117 ( .IN1(r851_n121), .IN2(r851_n116), .QN(r851_n119) );
  OR2X1 r851_U116 ( .IN2(r851_n116), .IN1(r851_n121), .Q(r851_n120) );
  NAND2X0 r851_U115 ( .IN1(r851_n119), .IN2(r851_n120), .QN(P2_N3899) );
  INVX0 r851_U114 ( .ZN(r851_n105), .INP(P2_N3748) );
  NAND2X0 r851_U113 ( .IN1(n7238), .IN2(r851_n105), .QN(r851_n117) );
  OR2X1 r851_U112 ( .IN2(n7238), .IN1(r851_n105), .Q(r851_n118) );
  NAND2X0 r851_U111 ( .IN1(r851_n117), .IN2(r851_n118), .QN(r851_n111) );
  NAND2X0 r851_U110 ( .IN1(n7242), .IN2(r851_n116), .QN(r851_n112) );
  OR2X1 r851_U109 ( .IN2(n7242), .IN1(r851_n116), .Q(r851_n114) );
  NAND2X0 r851_U108 ( .IN1(r851_n114), .IN2(r851_n115), .QN(r851_n113) );
  NAND2X0 r851_U107 ( .IN1(r851_n112), .IN2(r851_n113), .QN(r851_n106) );
  NAND2X0 r851_U106 ( .IN1(r851_n111), .IN2(r851_n106), .QN(r851_n109) );
  OR2X1 r851_U105 ( .IN2(r851_n106), .IN1(r851_n111), .Q(r851_n110) );
  NAND2X0 r851_U104 ( .IN1(r851_n109), .IN2(r851_n110), .QN(P2_N3900) );
  INVX0 r851_U103 ( .ZN(r851_n95), .INP(P2_N3749) );
  NAND2X0 r851_U102 ( .IN1(P2_N5096), .IN2(r851_n95), .QN(r851_n107) );
  OR2X1 r851_U101 ( .IN2(P2_N5096), .IN1(r851_n95), .Q(r851_n108) );
  NAND2X0 r851_U100 ( .IN1(r851_n107), .IN2(r851_n108), .QN(r851_n101) );
  NAND2X0 r851_U99 ( .IN1(n7238), .IN2(r851_n106), .QN(r851_n102) );
  OR2X1 r851_U98 ( .IN2(n7238), .IN1(r851_n106), .Q(r851_n104) );
  NAND2X0 r851_U97 ( .IN1(r851_n104), .IN2(r851_n105), .QN(r851_n103) );
  NAND2X0 r851_U96 ( .IN1(r851_n102), .IN2(r851_n103), .QN(r851_n96) );
  NAND2X0 r851_U95 ( .IN1(r851_n101), .IN2(r851_n96), .QN(r851_n99) );
  OR2X1 r851_U94 ( .IN2(r851_n96), .IN1(r851_n101), .Q(r851_n100) );
  NAND2X0 r851_U93 ( .IN1(r851_n99), .IN2(r851_n100), .QN(P2_N3901) );
  INVX0 r851_U92 ( .ZN(r851_n85), .INP(P2_N3750) );
  NAND2X0 r851_U91 ( .IN1(P2_N5097), .IN2(r851_n85), .QN(r851_n97) );
  OR2X1 r851_U90 ( .IN2(P2_N5097), .IN1(r851_n85), .Q(r851_n98) );
  NAND2X0 r851_U89 ( .IN1(r851_n97), .IN2(r851_n98), .QN(r851_n91) );
  NAND2X0 r851_U88 ( .IN1(P2_N5096), .IN2(r851_n96), .QN(r851_n92) );
  OR2X1 r851_U87 ( .IN2(P2_N5096), .IN1(r851_n96), .Q(r851_n94) );
  NAND2X0 r851_U86 ( .IN1(r851_n94), .IN2(r851_n95), .QN(r851_n93) );
  NAND2X0 r851_U85 ( .IN1(r851_n92), .IN2(r851_n93), .QN(r851_n86) );
  NAND2X0 r851_U84 ( .IN1(r851_n91), .IN2(r851_n86), .QN(r851_n89) );
  OR2X1 r851_U83 ( .IN2(r851_n86), .IN1(r851_n91), .Q(r851_n90) );
  NAND2X0 r851_U82 ( .IN1(r851_n89), .IN2(r851_n90), .QN(P2_N3902) );
  INVX0 r851_U81 ( .ZN(r851_n75), .INP(P2_N3751) );
  NAND2X0 r851_U80 ( .IN1(n7227), .IN2(r851_n75), .QN(r851_n87) );
  OR2X1 r851_U79 ( .IN2(n7227), .IN1(r851_n75), .Q(r851_n88) );
  NAND2X0 r851_U78 ( .IN1(r851_n87), .IN2(r851_n88), .QN(r851_n81) );
  NAND2X0 r851_U77 ( .IN1(P2_N5097), .IN2(r851_n86), .QN(r851_n82) );
  OR2X1 r851_U76 ( .IN2(P2_N5097), .IN1(r851_n86), .Q(r851_n84) );
  NAND2X0 r851_U75 ( .IN1(r851_n84), .IN2(r851_n85), .QN(r851_n83) );
  NAND2X0 r851_U74 ( .IN1(r851_n82), .IN2(r851_n83), .QN(r851_n76) );
  NAND2X0 r851_U73 ( .IN1(r851_n81), .IN2(r851_n76), .QN(r851_n79) );
  OR2X1 r851_U72 ( .IN2(r851_n76), .IN1(r851_n81), .Q(r851_n80) );
  NAND2X0 r851_U71 ( .IN1(r851_n79), .IN2(r851_n80), .QN(P2_N3903) );
  INVX0 r851_U70 ( .ZN(r851_n64), .INP(P2_N3752) );
  NAND2X0 r851_U69 ( .IN1(P2_N5099), .IN2(r851_n64), .QN(r851_n77) );
  OR2X1 r851_U68 ( .IN2(P2_N5099), .IN1(r851_n64), .Q(r851_n78) );
  NAND2X0 r851_U67 ( .IN1(r851_n77), .IN2(r851_n78), .QN(r851_n71) );
  NAND2X0 r851_U66 ( .IN1(n7227), .IN2(r851_n76), .QN(r851_n72) );
  OR2X1 r851_U65 ( .IN2(n7227), .IN1(r851_n76), .Q(r851_n74) );
  NAND2X0 r851_U64 ( .IN1(r851_n74), .IN2(r851_n75), .QN(r851_n73) );
  NAND2X0 r851_U63 ( .IN1(r851_n72), .IN2(r851_n73), .QN(r851_n65) );
  NAND2X0 r851_U62 ( .IN1(r851_n71), .IN2(r851_n65), .QN(r851_n69) );
  OR2X1 r851_U61 ( .IN2(r851_n65), .IN1(r851_n71), .Q(r851_n70) );
  NAND2X0 r851_U60 ( .IN1(r851_n69), .IN2(r851_n70), .QN(P2_N3904) );
  NAND2X0 r851_U245 ( .IN1(r851_n240), .IN2(r851_n241), .QN(r851_n234) );
  NAND2X0 r851_U244 ( .IN1(r851_n239), .IN2(r851_n234), .QN(r851_n237) );
  OR2X1 r851_U243 ( .IN2(r851_n234), .IN1(r851_n239), .Q(r851_n238) );
  NAND2X0 r851_U242 ( .IN1(r851_n237), .IN2(r851_n238), .QN(P2_N3888) );
  INVX0 r851_U241 ( .ZN(r851_n223), .INP(P2_N3737) );
  NAND2X0 r851_U240 ( .IN1(n7209), .IN2(r851_n223), .QN(r851_n235) );
  OR2X1 r851_U239 ( .IN2(n7209), .IN1(r851_n223), .Q(r851_n236) );
  NAND2X0 r851_U238 ( .IN1(r851_n235), .IN2(r851_n236), .QN(r851_n229) );
  NAND2X0 r851_U237 ( .IN1(n7210), .IN2(r851_n234), .QN(r851_n230) );
  OR2X1 r851_U236 ( .IN2(n7210), .IN1(r851_n234), .Q(r851_n232) );
  NAND2X0 r851_U235 ( .IN1(r851_n232), .IN2(r851_n233), .QN(r851_n231) );
  NAND2X0 r851_U234 ( .IN1(r851_n230), .IN2(r851_n231), .QN(r851_n224) );
  NAND2X0 r851_U233 ( .IN1(r851_n229), .IN2(r851_n224), .QN(r851_n227) );
  OR2X1 r851_U232 ( .IN2(r851_n224), .IN1(r851_n229), .Q(r851_n228) );
  NAND2X0 r851_U231 ( .IN1(r851_n227), .IN2(r851_n228), .QN(P2_N3889) );
  INVX0 r851_U230 ( .ZN(r851_n213), .INP(P2_N3738) );
  NAND2X0 r851_U229 ( .IN1(n7206), .IN2(r851_n213), .QN(r851_n225) );
  OR2X1 r851_U228 ( .IN2(n7206), .IN1(r851_n213), .Q(r851_n226) );
  NAND2X0 r851_U227 ( .IN1(r851_n225), .IN2(r851_n226), .QN(r851_n219) );
  NAND2X0 r851_U226 ( .IN1(n7209), .IN2(r851_n224), .QN(r851_n220) );
  OR2X1 r851_U225 ( .IN2(n7209), .IN1(r851_n224), .Q(r851_n222) );
  NAND2X0 r851_U224 ( .IN1(r851_n222), .IN2(r851_n223), .QN(r851_n221) );
  NAND2X0 r851_U223 ( .IN1(r851_n220), .IN2(r851_n221), .QN(r851_n214) );
  NAND2X0 r851_U222 ( .IN1(r851_n219), .IN2(r851_n214), .QN(r851_n217) );
  OR2X1 r851_U221 ( .IN2(r851_n214), .IN1(r851_n219), .Q(r851_n218) );
  NAND2X0 r851_U220 ( .IN1(r851_n217), .IN2(r851_n218), .QN(P2_N3890) );
  INVX0 r851_U219 ( .ZN(r851_n203), .INP(P2_N3739) );
  NAND2X0 r851_U218 ( .IN1(P2_N5086), .IN2(r851_n203), .QN(r851_n215) );
  OR2X1 r851_U217 ( .IN2(P2_N5086), .IN1(r851_n203), .Q(r851_n216) );
  NAND2X0 r851_U216 ( .IN1(r851_n215), .IN2(r851_n216), .QN(r851_n209) );
  NAND2X0 r851_U215 ( .IN1(n7206), .IN2(r851_n214), .QN(r851_n210) );
  OR2X1 r851_U214 ( .IN2(n7206), .IN1(r851_n214), .Q(r851_n212) );
  NAND2X0 r851_U213 ( .IN1(r851_n212), .IN2(r851_n213), .QN(r851_n211) );
  NAND2X0 r851_U212 ( .IN1(r851_n210), .IN2(r851_n211), .QN(r851_n204) );
  NAND2X0 r851_U211 ( .IN1(r851_n209), .IN2(r851_n204), .QN(r851_n207) );
  OR2X1 r851_U210 ( .IN2(r851_n204), .IN1(r851_n209), .Q(r851_n208) );
  NAND2X0 r851_U209 ( .IN1(r851_n207), .IN2(r851_n208), .QN(P2_N3891) );
  INVX0 r851_U208 ( .ZN(r851_n193), .INP(P2_N3740) );
  NAND2X0 r851_U207 ( .IN1(n7198), .IN2(r851_n193), .QN(r851_n205) );
  OR2X1 r851_U206 ( .IN2(n7198), .IN1(r851_n193), .Q(r851_n206) );
  NAND2X0 r851_U205 ( .IN1(r851_n205), .IN2(r851_n206), .QN(r851_n199) );
  NAND2X0 r851_U204 ( .IN1(P2_N5086), .IN2(r851_n204), .QN(r851_n200) );
  OR2X1 r851_U203 ( .IN2(P2_N5086), .IN1(r851_n204), .Q(r851_n202) );
  NAND2X0 r851_U202 ( .IN1(r851_n202), .IN2(r851_n203), .QN(r851_n201) );
  NAND2X0 r851_U201 ( .IN1(r851_n200), .IN2(r851_n201), .QN(r851_n194) );
  NAND2X0 r851_U200 ( .IN1(r851_n199), .IN2(r851_n194), .QN(r851_n197) );
  OR2X1 r851_U199 ( .IN2(r851_n194), .IN1(r851_n199), .Q(r851_n198) );
  NAND2X0 r851_U198 ( .IN1(r851_n197), .IN2(r851_n198), .QN(P2_N3892) );
  INVX0 r851_U197 ( .ZN(r851_n183), .INP(P2_N3741) );
  NAND2X0 r851_U196 ( .IN1(n7194), .IN2(r851_n183), .QN(r851_n195) );
  OR2X1 r851_U195 ( .IN2(n7194), .IN1(r851_n183), .Q(r851_n196) );
  NAND2X0 r851_U194 ( .IN1(r851_n195), .IN2(r851_n196), .QN(r851_n189) );
  NAND2X0 r851_U193 ( .IN1(n7198), .IN2(r851_n194), .QN(r851_n190) );
  OR2X1 r851_U192 ( .IN2(n7198), .IN1(r851_n194), .Q(r851_n192) );
  NAND2X0 r851_U191 ( .IN1(r851_n192), .IN2(r851_n193), .QN(r851_n191) );
  NAND2X0 r851_U190 ( .IN1(r851_n190), .IN2(r851_n191), .QN(r851_n184) );
  NAND2X0 r851_U189 ( .IN1(r851_n189), .IN2(r851_n184), .QN(r851_n187) );
  OR2X1 r851_U188 ( .IN2(r851_n184), .IN1(r851_n189), .Q(r851_n188) );
  NAND2X0 r851_U187 ( .IN1(r851_n187), .IN2(r851_n188), .QN(P2_N3893) );
  INVX0 r851_U186 ( .ZN(r851_n173), .INP(P2_N3742) );
  NAND2X0 r851_U185 ( .IN1(n7187), .IN2(r851_n173), .QN(r851_n185) );
  OR2X1 r851_U184 ( .IN2(n7187), .IN1(r851_n173), .Q(r851_n186) );
  NAND2X0 r851_U183 ( .IN1(r851_n185), .IN2(r851_n186), .QN(r851_n179) );
  NAND2X0 r851_U182 ( .IN1(n7194), .IN2(r851_n184), .QN(r851_n180) );
  OR2X1 r851_U181 ( .IN2(n7194), .IN1(r851_n184), .Q(r851_n182) );
  NAND2X0 r851_U180 ( .IN1(r851_n182), .IN2(r851_n183), .QN(r851_n181) );
  NAND2X0 r851_U179 ( .IN1(r851_n180), .IN2(r851_n181), .QN(r851_n174) );
  NAND2X0 r851_U178 ( .IN1(r851_n179), .IN2(r851_n174), .QN(r851_n177) );
  OR2X1 r851_U177 ( .IN2(r851_n174), .IN1(r851_n179), .Q(r851_n178) );
  NAND2X0 r851_U176 ( .IN1(r851_n177), .IN2(r851_n178), .QN(P2_N3894) );
  INVX0 r851_U175 ( .ZN(r851_n155), .INP(P2_N3743) );
  NAND2X0 r851_U174 ( .IN1(P2_N5090), .IN2(r851_n155), .QN(r851_n175) );
  OR2X1 r851_U173 ( .IN2(P2_N5090), .IN1(r851_n155), .Q(r851_n176) );
  NAND2X0 r851_U172 ( .IN1(r851_n175), .IN2(r851_n176), .QN(r851_n169) );
  NAND2X0 r851_U171 ( .IN1(n7187), .IN2(r851_n174), .QN(r851_n170) );
  OR2X1 r851_U170 ( .IN2(n7187), .IN1(r851_n174), .Q(r851_n172) );
  NAND2X0 r851_U169 ( .IN1(r851_n172), .IN2(r851_n173), .QN(r851_n171) );
  NAND2X0 r851_U168 ( .IN1(r851_n170), .IN2(r851_n171), .QN(r851_n156) );
  NAND2X0 r851_U167 ( .IN1(r851_n169), .IN2(r851_n156), .QN(r851_n167) );
  OR2X1 r851_U166 ( .IN2(r851_n156), .IN1(r851_n169), .Q(r851_n168) );
  NAND2X0 r851_U165 ( .IN1(r851_n167), .IN2(r851_n168), .QN(P2_N3895) );
  NAND2X0 r851_U164 ( .IN1(P2_N5072), .IN2(r851_n166), .QN(r851_n163) );
  NAND2X0 r851_U163 ( .IN1(P2_N3725), .IN2(n7184), .QN(r851_n164) );
  NAND2X0 r851_U162 ( .IN1(r851_n163), .IN2(r851_n164), .QN(r851_n161) );
  NAND2X0 r851_U161 ( .IN1(r851_n161), .IN2(r851_n162), .QN(r851_n159) );
  OR2X1 r851_U160 ( .IN2(r851_n162), .IN1(r851_n161), .Q(r851_n160) );
  NAND2X0 r851_U159 ( .IN1(r851_n159), .IN2(r851_n160), .QN(P2_N3877) );
  INVX0 r851_U158 ( .ZN(r851_n145), .INP(P2_N3744) );
  NAND2X0 r851_U157 ( .IN1(P2_N5091), .IN2(r851_n145), .QN(r851_n157) );
  OR2X1 r851_U156 ( .IN2(P2_N5091), .IN1(r851_n145), .Q(r851_n158) );
  NAND2X0 r851_U155 ( .IN1(r851_n157), .IN2(r851_n158), .QN(r851_n151) );
  NAND2X0 r851_U154 ( .IN1(P2_N5090), .IN2(r851_n156), .QN(r851_n152) );
  OR2X1 r851_U153 ( .IN2(P2_N5090), .IN1(r851_n156), .Q(r851_n154) );
  INVX0 r851_U321 ( .ZN(r851_n291), .INP(P2_N3724) );
  NOR2X0 r851_U320 ( .QN(r851_n287), .IN1(r851_n291), .IN2(n7035) );
  INVX0 r851_U319 ( .ZN(r851_n162), .INP(r851_n287) );
  NAND2X0 r851_U318 ( .IN1(n7035), .IN2(r851_n291), .QN(r851_n290) );
  NAND2X0 r851_U317 ( .IN1(r851_n162), .IN2(r851_n290), .QN(P2_N3876) );
  INVX0 r851_U316 ( .ZN(r851_n253), .INP(P2_N3734) );
  NAND2X0 r851_U315 ( .IN1(P2_N5081), .IN2(r851_n253), .QN(r851_n288) );
  OR2X1 r851_U314 ( .IN2(P2_N5081), .IN1(r851_n253), .Q(r851_n289) );
  NAND2X0 r851_U313 ( .IN1(r851_n288), .IN2(r851_n289), .QN(r851_n259) );
  NAND2X0 r851_U312 ( .IN1(P2_N5072), .IN2(r851_n162), .QN(r851_n284) );
  NAND2X0 r851_U310 ( .IN1(r851_n287), .IN2(n7184), .QN(r851_n286) );
  INVX0 r851_U309 ( .ZN(r851_n166), .INP(P2_N3725) );
  NAND2X0 r851_U308 ( .IN1(r851_n286), .IN2(r851_n166), .QN(r851_n285) );
  NAND2X0 r851_U307 ( .IN1(r851_n284), .IN2(r851_n285), .QN(r851_n53) );
  NAND2X0 r851_U306 ( .IN1(P2_N5073), .IN2(r851_n53), .QN(r851_n281) );
  OR2X1 r851_U305 ( .IN2(P2_N5073), .IN1(r851_n53), .Q(r851_n283) );
  INVX0 r851_U304 ( .ZN(r851_n56), .INP(P2_N3726) );
  NAND2X0 r851_U303 ( .IN1(r851_n283), .IN2(r851_n56), .QN(r851_n282) );
  NAND2X0 r851_U302 ( .IN1(r851_n281), .IN2(r851_n282), .QN(r851_n46) );
  NAND2X0 r851_U301 ( .IN1(n7177), .IN2(r851_n46), .QN(r851_n278) );
  OR2X1 r851_U300 ( .IN2(n7177), .IN1(r851_n46), .Q(r851_n280) );
  INVX0 r851_U299 ( .ZN(r851_n49), .INP(P2_N3727) );
  NAND2X0 r851_U298 ( .IN1(r851_n280), .IN2(r851_n49), .QN(r851_n279) );
  NAND2X0 r851_U297 ( .IN1(r851_n278), .IN2(r851_n279), .QN(r851_n39) );
  NAND2X0 r851_U296 ( .IN1(n7173), .IN2(r851_n39), .QN(r851_n275) );
  OR2X1 r851_U295 ( .IN2(n7173), .IN1(r851_n39), .Q(r851_n277) );
  INVX0 r851_U294 ( .ZN(r851_n42), .INP(P2_N3728) );
  NAND2X0 r851_U293 ( .IN1(r851_n277), .IN2(r851_n42), .QN(r851_n276) );
  NAND2X0 r851_U292 ( .IN1(r851_n275), .IN2(r851_n276), .QN(r851_n32) );
  NAND2X0 r851_U291 ( .IN1(P2_N5076), .IN2(r851_n32), .QN(r851_n272) );
  OR2X1 r851_U290 ( .IN2(P2_N5076), .IN1(r851_n32), .Q(r851_n274) );
  INVX0 r851_U289 ( .ZN(r851_n35), .INP(P2_N3729) );
  NAND2X0 r851_U288 ( .IN1(r851_n274), .IN2(r851_n35), .QN(r851_n273) );
  NAND2X0 r851_U287 ( .IN1(r851_n272), .IN2(r851_n273), .QN(r851_n25) );
  NAND2X0 r851_U286 ( .IN1(n7162), .IN2(r851_n25), .QN(r851_n269) );
  OR2X1 r851_U285 ( .IN2(n7162), .IN1(r851_n25), .Q(r851_n271) );
  INVX0 r851_U284 ( .ZN(r851_n28), .INP(P2_N3730) );
  NAND2X0 r851_U283 ( .IN1(r851_n271), .IN2(r851_n28), .QN(r851_n270) );
  NAND2X0 r851_U282 ( .IN1(r851_n269), .IN2(r851_n270), .QN(r851_n18) );
  NAND2X0 r851_U281 ( .IN1(P2_N5078), .IN2(r851_n18), .QN(r851_n266) );
  OR2X1 r851_U280 ( .IN2(P2_N5078), .IN1(r851_n18), .Q(r851_n268) );
  INVX0 r851_U279 ( .ZN(r851_n21), .INP(P2_N3731) );
  NAND2X0 r851_U278 ( .IN1(r851_n268), .IN2(r851_n21), .QN(r851_n267) );
  NAND2X0 r851_U277 ( .IN1(r851_n266), .IN2(r851_n267), .QN(r851_n11) );
  NAND2X0 r851_U276 ( .IN1(n7154), .IN2(r851_n11), .QN(r851_n263) );
  OR2X1 r851_U275 ( .IN2(n7154), .IN1(r851_n11), .Q(r851_n265) );
  INVX0 r851_U274 ( .ZN(r851_n14), .INP(P2_N3732) );
  NAND2X0 r851_U273 ( .IN1(r851_n265), .IN2(r851_n14), .QN(r851_n264) );
  NAND2X0 r851_U272 ( .IN1(r851_n263), .IN2(r851_n264), .QN(r851_n4) );
  NAND2X0 r851_U271 ( .IN1(n7151), .IN2(r851_n4), .QN(r851_n260) );
  OR2X1 r851_U270 ( .IN2(n7151), .IN1(r851_n4), .Q(r851_n262) );
  INVX0 r851_U269 ( .ZN(r851_n7), .INP(P2_N3733) );
  NAND2X0 r851_U268 ( .IN1(r851_n262), .IN2(r851_n7), .QN(r851_n261) );
  NAND2X0 r851_U267 ( .IN1(r851_n260), .IN2(r851_n261), .QN(r851_n254) );
  NAND2X0 r851_U266 ( .IN1(r851_n259), .IN2(r851_n254), .QN(r851_n257) );
  OR2X1 r851_U265 ( .IN2(r851_n254), .IN1(r851_n259), .Q(r851_n258) );
  NAND2X0 r851_U264 ( .IN1(r851_n257), .IN2(r851_n258), .QN(P2_N3886) );
  INVX0 r851_U263 ( .ZN(r851_n243), .INP(P2_N3735) );
  NAND2X0 r851_U262 ( .IN1(P2_N5082), .IN2(r851_n243), .QN(r851_n255) );
  OR2X1 r851_U261 ( .IN2(P2_N5082), .IN1(r851_n243), .Q(r851_n256) );
  NAND2X0 r851_U260 ( .IN1(r851_n255), .IN2(r851_n256), .QN(r851_n249) );
  NAND2X0 r851_U259 ( .IN1(P2_N5081), .IN2(r851_n254), .QN(r851_n250) );
  OR2X1 r851_U258 ( .IN2(P2_N5081), .IN1(r851_n254), .Q(r851_n252) );
  NAND2X0 r851_U257 ( .IN1(r851_n252), .IN2(r851_n253), .QN(r851_n251) );
  NAND2X0 r851_U256 ( .IN1(r851_n250), .IN2(r851_n251), .QN(r851_n244) );
  NAND2X0 r851_U255 ( .IN1(r851_n249), .IN2(r851_n244), .QN(r851_n247) );
  OR2X1 r851_U254 ( .IN2(r851_n244), .IN1(r851_n249), .Q(r851_n248) );
  NAND2X0 r851_U253 ( .IN1(r851_n247), .IN2(r851_n248), .QN(P2_N3887) );
  INVX0 r851_U252 ( .ZN(r851_n233), .INP(P2_N3736) );
  NAND2X0 r851_U251 ( .IN1(n7210), .IN2(r851_n233), .QN(r851_n245) );
  OR2X1 r851_U250 ( .IN2(n7210), .IN1(r851_n233), .Q(r851_n246) );
  NAND2X0 r851_U249 ( .IN1(r851_n245), .IN2(r851_n246), .QN(r851_n239) );
  NAND2X0 r851_U248 ( .IN1(P2_N5082), .IN2(r851_n244), .QN(r851_n240) );
  OR2X1 r851_U247 ( .IN2(P2_N5082), .IN1(r851_n244), .Q(r851_n242) );
  NAND2X0 r851_U246 ( .IN1(r851_n242), .IN2(r851_n243), .QN(r851_n241) );
  OR2X1 r854_U6 ( .IN2(P2_N4106), .IN1(n7149), .Q(r854_n5) );
  NAND2X0 r854_U5 ( .IN1(P2_N4106), .IN2(n7149), .QN(r854_n6) );
  NAND2X0 r854_U4 ( .IN1(r854_n5), .IN2(r854_n6), .QN(r854_n4) );
  NOR2X0 r854_U3 ( .QN(r854_n1), .IN1(r854_n3), .IN2(r854_n4) );
  AND2X1 r854_U2 ( .IN1(r854_n3), .IN2(r854_n4), .Q(r854_n2) );
  NOR2X0 r854_U1 ( .QN(P2_N4287), .IN1(r854_n1), .IN2(r854_n2) );
  NAND2X0 r854_U100 ( .IN1(n7237), .IN2(r854_n97), .QN(r854_n94) );
  OR2X1 r854_U99 ( .IN2(n7237), .IN1(r854_n97), .Q(r854_n96) );
  NAND2X0 r854_U98 ( .IN1(P2_N4122), .IN2(r854_n96), .QN(r854_n95) );
  NAND2X0 r854_U97 ( .IN1(r854_n94), .IN2(r854_n95), .QN(r854_n87) );
  OR2X1 r854_U95 ( .IN2(P2_N4123), .IN1(n7229), .Q(r854_n91) );
  NAND2X0 r854_U94 ( .IN1(P2_N4123), .IN2(n7229), .QN(r854_n92) );
  NAND2X0 r854_U93 ( .IN1(r854_n91), .IN2(r854_n92), .QN(r854_n90) );
  NOR2X0 r854_U92 ( .QN(r854_n88), .IN1(r854_n87), .IN2(r854_n90) );
  AND2X1 r854_U91 ( .IN1(r854_n87), .IN2(r854_n90), .Q(r854_n89) );
  NOR2X0 r854_U90 ( .QN(P2_N4304), .IN1(r854_n88), .IN2(r854_n89) );
  NAND2X0 r854_U89 ( .IN1(n7231), .IN2(r854_n87), .QN(r854_n84) );
  OR2X1 r854_U88 ( .IN2(n7231), .IN1(r854_n87), .Q(r854_n86) );
  NAND2X0 r854_U87 ( .IN1(P2_N4123), .IN2(r854_n86), .QN(r854_n85) );
  NAND2X0 r854_U86 ( .IN1(r854_n84), .IN2(r854_n85), .QN(r854_n77) );
  OR2X1 r854_U84 ( .IN2(P2_N4124), .IN1(n7224), .Q(r854_n81) );
  NAND2X0 r854_U83 ( .IN1(P2_N4124), .IN2(n7224), .QN(r854_n82) );
  NAND2X0 r854_U82 ( .IN1(r854_n81), .IN2(r854_n82), .QN(r854_n80) );
  NOR2X0 r854_U81 ( .QN(r854_n78), .IN1(r854_n77), .IN2(r854_n80) );
  AND2X1 r854_U80 ( .IN1(r854_n77), .IN2(r854_n80), .Q(r854_n79) );
  NOR2X0 r854_U79 ( .QN(P2_N4305), .IN1(r854_n78), .IN2(r854_n79) );
  NAND2X0 r854_U78 ( .IN1(n7227), .IN2(r854_n77), .QN(r854_n74) );
  OR2X1 r854_U77 ( .IN2(n7227), .IN1(r854_n77), .Q(r854_n76) );
  NAND2X0 r854_U76 ( .IN1(P2_N4124), .IN2(r854_n76), .QN(r854_n75) );
  NAND2X0 r854_U75 ( .IN1(r854_n74), .IN2(r854_n75), .QN(r854_n64) );
  OR2X1 r854_U73 ( .IN2(P2_N4125), .IN1(n7222), .Q(r854_n71) );
  NAND2X0 r854_U72 ( .IN1(P2_N4125), .IN2(n7222), .QN(r854_n72) );
  NAND2X0 r854_U71 ( .IN1(r854_n71), .IN2(r854_n72), .QN(r854_n70) );
  NOR2X0 r854_U70 ( .QN(r854_n68), .IN1(r854_n64), .IN2(r854_n70) );
  AND2X1 r854_U69 ( .IN1(r854_n64), .IN2(r854_n70), .Q(r854_n69) );
  NOR2X0 r854_U68 ( .QN(P2_N4306), .IN1(r854_n68), .IN2(r854_n69) );
  OR2X1 r854_U66 ( .IN2(P2_N4126), .IN1(n7266), .Q(r854_n65) );
  NAND2X0 r854_U65 ( .IN1(P2_N4126), .IN2(n7266), .QN(r854_n66) );
  NAND2X0 r854_U64 ( .IN1(r854_n65), .IN2(r854_n66), .QN(r854_n60) );
  NAND2X0 r854_U63 ( .IN1(P2_N5099), .IN2(r854_n64), .QN(r854_n61) );
  OR2X1 r854_U62 ( .IN2(P2_N5099), .IN1(r854_n64), .Q(r854_n63) );
  NAND2X0 r854_U61 ( .IN1(P2_N4125), .IN2(r854_n63), .QN(r854_n62) );
  NAND2X0 r854_U60 ( .IN1(r854_n61), .IN2(r854_n62), .QN(r854_n59) );
  NOR2X0 r854_U59 ( .QN(r854_n57), .IN1(r854_n60), .IN2(r854_n59) );
  AND2X1 r854_U58 ( .IN1(r854_n59), .IN2(r854_n60), .Q(r854_n58) );
  NOR2X0 r854_U57 ( .QN(P2_N4307), .IN1(r854_n57), .IN2(r854_n58) );
  OR2X1 r854_U55 ( .IN2(P2_N4099), .IN1(n7182), .Q(r854_n54) );
  NAND2X0 r854_U54 ( .IN1(P2_N4099), .IN2(n7182), .QN(r854_n55) );
  NAND2X0 r854_U53 ( .IN1(r854_n54), .IN2(r854_n55), .QN(r854_n53) );
  NOR2X0 r854_U52 ( .QN(r854_n50), .IN1(r854_n52), .IN2(r854_n53) );
  AND2X1 r854_U51 ( .IN1(r854_n52), .IN2(r854_n53), .Q(r854_n51) );
  NOR2X0 r854_U50 ( .QN(P2_N4280), .IN1(r854_n50), .IN2(r854_n51) );
  OR2X1 r854_U48 ( .IN2(P2_N4100), .IN1(n7178), .Q(r854_n47) );
  NAND2X0 r854_U47 ( .IN1(P2_N4100), .IN2(n7178), .QN(r854_n48) );
  NAND2X0 r854_U46 ( .IN1(r854_n47), .IN2(r854_n48), .QN(r854_n46) );
  NOR2X0 r854_U45 ( .QN(r854_n43), .IN1(r854_n45), .IN2(r854_n46) );
  AND2X1 r854_U44 ( .IN1(r854_n45), .IN2(r854_n46), .Q(r854_n44) );
  NOR2X0 r854_U43 ( .QN(P2_N4281), .IN1(r854_n43), .IN2(r854_n44) );
  OR2X1 r854_U41 ( .IN2(P2_N4101), .IN1(n7174), .Q(r854_n40) );
  NAND2X0 r854_U40 ( .IN1(P2_N4101), .IN2(n7174), .QN(r854_n41) );
  NAND2X0 r854_U39 ( .IN1(r854_n40), .IN2(r854_n41), .QN(r854_n39) );
  NOR2X0 r854_U38 ( .QN(r854_n36), .IN1(r854_n38), .IN2(r854_n39) );
  AND2X1 r854_U37 ( .IN1(r854_n38), .IN2(r854_n39), .Q(r854_n37) );
  NOR2X0 r854_U36 ( .QN(P2_N4282), .IN1(r854_n36), .IN2(r854_n37) );
  OR2X1 r854_U34 ( .IN2(P2_N4102), .IN1(n7166), .Q(r854_n33) );
  NAND2X0 r854_U33 ( .IN1(P2_N4102), .IN2(n7166), .QN(r854_n34) );
  NAND2X0 r854_U32 ( .IN1(r854_n33), .IN2(r854_n34), .QN(r854_n32) );
  NOR2X0 r854_U31 ( .QN(r854_n29), .IN1(r854_n31), .IN2(r854_n32) );
  AND2X1 r854_U30 ( .IN1(r854_n31), .IN2(r854_n32), .Q(r854_n30) );
  NOR2X0 r854_U29 ( .QN(P2_N4283), .IN1(r854_n29), .IN2(r854_n30) );
  OR2X1 r854_U27 ( .IN2(P2_N4103), .IN1(n7164), .Q(r854_n26) );
  NAND2X0 r854_U26 ( .IN1(P2_N4103), .IN2(n7164), .QN(r854_n27) );
  NAND2X0 r854_U25 ( .IN1(r854_n26), .IN2(r854_n27), .QN(r854_n25) );
  NOR2X0 r854_U24 ( .QN(r854_n22), .IN1(r854_n24), .IN2(r854_n25) );
  AND2X1 r854_U23 ( .IN1(r854_n24), .IN2(r854_n25), .Q(r854_n23) );
  NOR2X0 r854_U22 ( .QN(P2_N4284), .IN1(r854_n22), .IN2(r854_n23) );
  OR2X1 r854_U20 ( .IN2(P2_N4104), .IN1(n7157), .Q(r854_n19) );
  NAND2X0 r854_U19 ( .IN1(P2_N4104), .IN2(n7157), .QN(r854_n20) );
  NAND2X0 r854_U18 ( .IN1(r854_n19), .IN2(r854_n20), .QN(r854_n18) );
  NOR2X0 r854_U17 ( .QN(r854_n15), .IN1(r854_n17), .IN2(r854_n18) );
  AND2X1 r854_U16 ( .IN1(r854_n17), .IN2(r854_n18), .Q(r854_n16) );
  NOR2X0 r854_U15 ( .QN(P2_N4285), .IN1(r854_n15), .IN2(r854_n16) );
  OR2X1 r854_U13 ( .IN2(P2_N4105), .IN1(n7153), .Q(r854_n12) );
  NAND2X0 r854_U12 ( .IN1(P2_N4105), .IN2(n7153), .QN(r854_n13) );
  NAND2X0 r854_U11 ( .IN1(r854_n12), .IN2(r854_n13), .QN(r854_n11) );
  NOR2X0 r854_U10 ( .QN(r854_n8), .IN1(r854_n10), .IN2(r854_n11) );
  AND2X1 r854_U9 ( .IN1(r854_n10), .IN2(r854_n11), .Q(r854_n9) );
  NOR2X0 r854_U8 ( .QN(P2_N4286), .IN1(r854_n8), .IN2(r854_n9) );
  OR2X1 r854_U193 ( .IN2(n7194), .IN1(r854_n184), .Q(r854_n183) );
  NAND2X0 r854_U192 ( .IN1(P2_N4114), .IN2(r854_n183), .QN(r854_n182) );
  NAND2X0 r854_U191 ( .IN1(r854_n181), .IN2(r854_n182), .QN(r854_n174) );
  OR2X1 r854_U189 ( .IN2(P2_N4115), .IN1(n7188), .Q(r854_n178) );
  NAND2X0 r854_U188 ( .IN1(P2_N4115), .IN2(n7188), .QN(r854_n179) );
  NAND2X0 r854_U187 ( .IN1(r854_n178), .IN2(r854_n179), .QN(r854_n177) );
  NOR2X0 r854_U186 ( .QN(r854_n175), .IN1(r854_n174), .IN2(r854_n177) );
  AND2X1 r854_U185 ( .IN1(r854_n174), .IN2(r854_n177), .Q(r854_n176) );
  NOR2X0 r854_U184 ( .QN(P2_N4296), .IN1(r854_n175), .IN2(r854_n176) );
  NAND2X0 r854_U183 ( .IN1(n7187), .IN2(r854_n174), .QN(r854_n171) );
  OR2X1 r854_U182 ( .IN2(n7187), .IN1(r854_n174), .Q(r854_n173) );
  NAND2X0 r854_U181 ( .IN1(P2_N4115), .IN2(r854_n173), .QN(r854_n172) );
  NAND2X0 r854_U180 ( .IN1(r854_n171), .IN2(r854_n172), .QN(r854_n157) );
  OR2X1 r854_U178 ( .IN2(P2_N4116), .IN1(n7264), .Q(r854_n168) );
  NAND2X0 r854_U177 ( .IN1(P2_N4116), .IN2(n7264), .QN(r854_n169) );
  NAND2X0 r854_U176 ( .IN1(r854_n168), .IN2(r854_n169), .QN(r854_n167) );
  NOR2X0 r854_U175 ( .QN(r854_n165), .IN1(r854_n157), .IN2(r854_n167) );
  AND2X1 r854_U174 ( .IN1(r854_n157), .IN2(r854_n167), .Q(r854_n166) );
  NOR2X0 r854_U173 ( .QN(P2_N4297), .IN1(r854_n165), .IN2(r854_n166) );
  OR2X1 r854_U172 ( .IN2(P2_N4098), .IN1(n7186), .Q(r854_n162) );
  NAND2X0 r854_U171 ( .IN1(P2_N4098), .IN2(n7186), .QN(r854_n163) );
  NAND2X0 r854_U170 ( .IN1(r854_n162), .IN2(r854_n163), .QN(r854_n160) );
  NAND2X0 r854_U169 ( .IN1(r854_n160), .IN2(r854_n161), .QN(r854_n158) );
  OR2X1 r854_U168 ( .IN2(r854_n161), .IN1(r854_n160), .Q(r854_n159) );
  NAND2X0 r854_U167 ( .IN1(r854_n158), .IN2(r854_n159), .QN(P2_N4279) );
  NAND2X0 r854_U166 ( .IN1(n7263), .IN2(r854_n157), .QN(r854_n154) );
  OR2X1 r854_U165 ( .IN2(n7263), .IN1(r854_n157), .Q(r854_n156) );
  NAND2X0 r854_U164 ( .IN1(P2_N4116), .IN2(r854_n156), .QN(r854_n155) );
  NAND2X0 r854_U163 ( .IN1(r854_n154), .IN2(r854_n155), .QN(r854_n147) );
  OR2X1 r854_U161 ( .IN2(P2_N4117), .IN1(n7260), .Q(r854_n151) );
  NAND2X0 r854_U160 ( .IN1(P2_N4117), .IN2(n7260), .QN(r854_n152) );
  NAND2X0 r854_U159 ( .IN1(r854_n151), .IN2(r854_n152), .QN(r854_n150) );
  NOR2X0 r854_U158 ( .QN(r854_n148), .IN1(r854_n147), .IN2(r854_n150) );
  AND2X1 r854_U157 ( .IN1(r854_n147), .IN2(r854_n150), .Q(r854_n149) );
  NOR2X0 r854_U156 ( .QN(P2_N4298), .IN1(r854_n148), .IN2(r854_n149) );
  NAND2X0 r854_U155 ( .IN1(n7259), .IN2(r854_n147), .QN(r854_n144) );
  OR2X1 r854_U154 ( .IN2(n7259), .IN1(r854_n147), .Q(r854_n146) );
  NAND2X0 r854_U153 ( .IN1(P2_N4117), .IN2(r854_n146), .QN(r854_n145) );
  NAND2X0 r854_U152 ( .IN1(r854_n144), .IN2(r854_n145), .QN(r854_n137) );
  OR2X1 r854_U150 ( .IN2(P2_N4118), .IN1(n7253), .Q(r854_n141) );
  NAND2X0 r854_U149 ( .IN1(P2_N4118), .IN2(n7253), .QN(r854_n142) );
  NAND2X0 r854_U148 ( .IN1(r854_n141), .IN2(r854_n142), .QN(r854_n140) );
  NOR2X0 r854_U147 ( .QN(r854_n138), .IN1(r854_n137), .IN2(r854_n140) );
  AND2X1 r854_U146 ( .IN1(r854_n137), .IN2(r854_n140), .Q(r854_n139) );
  NOR2X0 r854_U145 ( .QN(P2_N4299), .IN1(r854_n138), .IN2(r854_n139) );
  NAND2X0 r854_U144 ( .IN1(n7252), .IN2(r854_n137), .QN(r854_n134) );
  OR2X1 r854_U143 ( .IN2(n7252), .IN1(r854_n137), .Q(r854_n136) );
  NAND2X0 r854_U142 ( .IN1(P2_N4118), .IN2(r854_n136), .QN(r854_n135) );
  NAND2X0 r854_U141 ( .IN1(r854_n134), .IN2(r854_n135), .QN(r854_n127) );
  OR2X1 r854_U139 ( .IN2(P2_N4119), .IN1(n7248), .Q(r854_n131) );
  NAND2X0 r854_U138 ( .IN1(P2_N4119), .IN2(n7248), .QN(r854_n132) );
  NAND2X0 r854_U137 ( .IN1(r854_n131), .IN2(r854_n132), .QN(r854_n130) );
  NOR2X0 r854_U136 ( .QN(r854_n128), .IN1(r854_n127), .IN2(r854_n130) );
  AND2X1 r854_U135 ( .IN1(r854_n127), .IN2(r854_n130), .Q(r854_n129) );
  NOR2X0 r854_U134 ( .QN(P2_N4300), .IN1(r854_n128), .IN2(r854_n129) );
  NAND2X0 r854_U133 ( .IN1(P2_N5093), .IN2(r854_n127), .QN(r854_n124) );
  OR2X1 r854_U132 ( .IN2(n7247), .IN1(r854_n127), .Q(r854_n126) );
  NAND2X0 r854_U131 ( .IN1(P2_N4119), .IN2(r854_n126), .QN(r854_n125) );
  NAND2X0 r854_U130 ( .IN1(r854_n124), .IN2(r854_n125), .QN(r854_n117) );
  OR2X1 r854_U128 ( .IN2(P2_N4120), .IN1(n7243), .Q(r854_n121) );
  NAND2X0 r854_U127 ( .IN1(P2_N4120), .IN2(n7243), .QN(r854_n122) );
  NAND2X0 r854_U126 ( .IN1(r854_n121), .IN2(r854_n122), .QN(r854_n120) );
  NOR2X0 r854_U125 ( .QN(r854_n118), .IN1(r854_n117), .IN2(r854_n120) );
  AND2X1 r854_U124 ( .IN1(r854_n117), .IN2(r854_n120), .Q(r854_n119) );
  NOR2X0 r854_U123 ( .QN(P2_N4301), .IN1(r854_n118), .IN2(r854_n119) );
  NAND2X0 r854_U122 ( .IN1(n7242), .IN2(r854_n117), .QN(r854_n114) );
  OR2X1 r854_U121 ( .IN2(n7242), .IN1(r854_n117), .Q(r854_n116) );
  NAND2X0 r854_U120 ( .IN1(P2_N4120), .IN2(r854_n116), .QN(r854_n115) );
  NAND2X0 r854_U119 ( .IN1(r854_n114), .IN2(r854_n115), .QN(r854_n107) );
  OR2X1 r854_U117 ( .IN2(P2_N4121), .IN1(n7239), .Q(r854_n111) );
  NAND2X0 r854_U116 ( .IN1(P2_N4121), .IN2(n7239), .QN(r854_n112) );
  NAND2X0 r854_U115 ( .IN1(r854_n111), .IN2(r854_n112), .QN(r854_n110) );
  NOR2X0 r854_U114 ( .QN(r854_n108), .IN1(r854_n107), .IN2(r854_n110) );
  AND2X1 r854_U113 ( .IN1(r854_n107), .IN2(r854_n110), .Q(r854_n109) );
  NOR2X0 r854_U112 ( .QN(P2_N4302), .IN1(r854_n108), .IN2(r854_n109) );
  NAND2X0 r854_U111 ( .IN1(n7238), .IN2(r854_n107), .QN(r854_n104) );
  OR2X1 r854_U110 ( .IN2(n7238), .IN1(r854_n107), .Q(r854_n106) );
  NAND2X0 r854_U109 ( .IN1(P2_N4121), .IN2(r854_n106), .QN(r854_n105) );
  NAND2X0 r854_U108 ( .IN1(r854_n104), .IN2(r854_n105), .QN(r854_n97) );
  OR2X1 r854_U106 ( .IN2(P2_N4122), .IN1(n7234), .Q(r854_n101) );
  NAND2X0 r854_U105 ( .IN1(P2_N4122), .IN2(n7234), .QN(r854_n102) );
  NAND2X0 r854_U104 ( .IN1(r854_n101), .IN2(r854_n102), .QN(r854_n100) );
  NOR2X0 r854_U103 ( .QN(r854_n98), .IN1(r854_n97), .IN2(r854_n100) );
  AND2X1 r854_U102 ( .IN1(r854_n97), .IN2(r854_n100), .Q(r854_n99) );
  NOR2X0 r854_U101 ( .QN(P2_N4303), .IN1(r854_n98), .IN2(r854_n99) );
  NAND2X0 r854_U286 ( .IN1(P2_N5079), .IN2(r854_n10), .QN(r854_n264) );
  OR2X1 r854_U285 ( .IN2(P2_N5079), .IN1(r854_n10), .Q(r854_n266) );
  NAND2X0 r854_U284 ( .IN1(P2_N4105), .IN2(r854_n266), .QN(r854_n265) );
  NAND2X0 r854_U283 ( .IN1(r854_n264), .IN2(r854_n265), .QN(r854_n3) );
  NAND2X0 r854_U282 ( .IN1(n7151), .IN2(r854_n3), .QN(r854_n261) );
  OR2X1 r854_U281 ( .IN2(n7151), .IN1(r854_n3), .Q(r854_n263) );
  NAND2X0 r854_U280 ( .IN1(P2_N4106), .IN2(r854_n263), .QN(r854_n262) );
  NAND2X0 r854_U279 ( .IN1(r854_n261), .IN2(r854_n262), .QN(r854_n254) );
  OR2X1 r854_U277 ( .IN2(P2_N4107), .IN1(n7219), .Q(r854_n258) );
  NAND2X0 r854_U276 ( .IN1(P2_N4107), .IN2(n7219), .QN(r854_n259) );
  NAND2X0 r854_U275 ( .IN1(r854_n258), .IN2(r854_n259), .QN(r854_n257) );
  NOR2X0 r854_U274 ( .QN(r854_n255), .IN1(r854_n254), .IN2(r854_n257) );
  AND2X1 r854_U273 ( .IN1(r854_n254), .IN2(r854_n257), .Q(r854_n256) );
  NOR2X0 r854_U272 ( .QN(P2_N4288), .IN1(r854_n255), .IN2(r854_n256) );
  NAND2X0 r854_U271 ( .IN1(P2_N5081), .IN2(r854_n254), .QN(r854_n251) );
  OR2X1 r854_U270 ( .IN2(P2_N5081), .IN1(r854_n254), .Q(r854_n253) );
  NAND2X0 r854_U269 ( .IN1(P2_N4107), .IN2(r854_n253), .QN(r854_n252) );
  NAND2X0 r854_U268 ( .IN1(r854_n251), .IN2(r854_n252), .QN(r854_n244) );
  OR2X1 r854_U266 ( .IN2(P2_N4108), .IN1(n7214), .Q(r854_n248) );
  NAND2X0 r854_U265 ( .IN1(P2_N4108), .IN2(n7214), .QN(r854_n249) );
  NAND2X0 r854_U264 ( .IN1(r854_n248), .IN2(r854_n249), .QN(r854_n247) );
  NOR2X0 r854_U263 ( .QN(r854_n245), .IN1(r854_n244), .IN2(r854_n247) );
  AND2X1 r854_U262 ( .IN1(r854_n244), .IN2(r854_n247), .Q(r854_n246) );
  NOR2X0 r854_U261 ( .QN(P2_N4289), .IN1(r854_n245), .IN2(r854_n246) );
  NAND2X0 r854_U260 ( .IN1(P2_N5082), .IN2(r854_n244), .QN(r854_n241) );
  OR2X1 r854_U259 ( .IN2(P2_N5082), .IN1(r854_n244), .Q(r854_n243) );
  NAND2X0 r854_U258 ( .IN1(P2_N4108), .IN2(r854_n243), .QN(r854_n242) );
  NAND2X0 r854_U257 ( .IN1(r854_n241), .IN2(r854_n242), .QN(r854_n234) );
  OR2X1 r854_U255 ( .IN2(P2_N4109), .IN1(n7211), .Q(r854_n238) );
  NAND2X0 r854_U254 ( .IN1(P2_N4109), .IN2(n7211), .QN(r854_n239) );
  NAND2X0 r854_U253 ( .IN1(r854_n238), .IN2(r854_n239), .QN(r854_n237) );
  NOR2X0 r854_U252 ( .QN(r854_n235), .IN1(r854_n234), .IN2(r854_n237) );
  AND2X1 r854_U251 ( .IN1(r854_n234), .IN2(r854_n237), .Q(r854_n236) );
  NOR2X0 r854_U250 ( .QN(P2_N4290), .IN1(r854_n235), .IN2(r854_n236) );
  NAND2X0 r854_U249 ( .IN1(n7210), .IN2(r854_n234), .QN(r854_n231) );
  OR2X1 r854_U248 ( .IN2(n7210), .IN1(r854_n234), .Q(r854_n233) );
  NAND2X0 r854_U247 ( .IN1(P2_N4109), .IN2(r854_n233), .QN(r854_n232) );
  NAND2X0 r854_U246 ( .IN1(r854_n231), .IN2(r854_n232), .QN(r854_n224) );
  OR2X1 r854_U244 ( .IN2(P2_N4110), .IN1(n7208), .Q(r854_n228) );
  NAND2X0 r854_U243 ( .IN1(P2_N4110), .IN2(n7208), .QN(r854_n229) );
  NAND2X0 r854_U242 ( .IN1(r854_n228), .IN2(r854_n229), .QN(r854_n227) );
  NOR2X0 r854_U241 ( .QN(r854_n225), .IN1(r854_n224), .IN2(r854_n227) );
  AND2X1 r854_U240 ( .IN1(r854_n224), .IN2(r854_n227), .Q(r854_n226) );
  NOR2X0 r854_U239 ( .QN(P2_N4291), .IN1(r854_n225), .IN2(r854_n226) );
  NAND2X0 r854_U238 ( .IN1(P2_N5084), .IN2(r854_n224), .QN(r854_n221) );
  OR2X1 r854_U237 ( .IN2(P2_N5084), .IN1(r854_n224), .Q(r854_n223) );
  NAND2X0 r854_U236 ( .IN1(P2_N4110), .IN2(r854_n223), .QN(r854_n222) );
  NAND2X0 r854_U235 ( .IN1(r854_n221), .IN2(r854_n222), .QN(r854_n214) );
  OR2X1 r854_U233 ( .IN2(P2_N4111), .IN1(n7205), .Q(r854_n218) );
  NAND2X0 r854_U232 ( .IN1(P2_N4111), .IN2(n7205), .QN(r854_n219) );
  NAND2X0 r854_U231 ( .IN1(r854_n218), .IN2(r854_n219), .QN(r854_n217) );
  NOR2X0 r854_U230 ( .QN(r854_n215), .IN1(r854_n214), .IN2(r854_n217) );
  AND2X1 r854_U229 ( .IN1(r854_n214), .IN2(r854_n217), .Q(r854_n216) );
  NOR2X0 r854_U228 ( .QN(P2_N4292), .IN1(r854_n215), .IN2(r854_n216) );
  NAND2X0 r854_U227 ( .IN1(P2_N5085), .IN2(r854_n214), .QN(r854_n211) );
  OR2X1 r854_U226 ( .IN2(P2_N5085), .IN1(r854_n214), .Q(r854_n213) );
  NAND2X0 r854_U225 ( .IN1(P2_N4111), .IN2(r854_n213), .QN(r854_n212) );
  NAND2X0 r854_U224 ( .IN1(r854_n211), .IN2(r854_n212), .QN(r854_n204) );
  OR2X1 r854_U222 ( .IN2(P2_N4112), .IN1(n7201), .Q(r854_n208) );
  NAND2X0 r854_U221 ( .IN1(P2_N4112), .IN2(n7201), .QN(r854_n209) );
  NAND2X0 r854_U220 ( .IN1(r854_n208), .IN2(r854_n209), .QN(r854_n207) );
  NOR2X0 r854_U219 ( .QN(r854_n205), .IN1(r854_n204), .IN2(r854_n207) );
  AND2X1 r854_U218 ( .IN1(r854_n204), .IN2(r854_n207), .Q(r854_n206) );
  NOR2X0 r854_U217 ( .QN(P2_N4293), .IN1(r854_n205), .IN2(r854_n206) );
  NAND2X0 r854_U216 ( .IN1(P2_N5086), .IN2(r854_n204), .QN(r854_n201) );
  OR2X1 r854_U215 ( .IN2(P2_N5086), .IN1(r854_n204), .Q(r854_n203) );
  NAND2X0 r854_U214 ( .IN1(P2_N4112), .IN2(r854_n203), .QN(r854_n202) );
  NAND2X0 r854_U213 ( .IN1(r854_n201), .IN2(r854_n202), .QN(r854_n194) );
  OR2X1 r854_U211 ( .IN2(P2_N4113), .IN1(n7197), .Q(r854_n198) );
  NAND2X0 r854_U210 ( .IN1(P2_N4113), .IN2(n7197), .QN(r854_n199) );
  NAND2X0 r854_U209 ( .IN1(r854_n198), .IN2(r854_n199), .QN(r854_n197) );
  NOR2X0 r854_U208 ( .QN(r854_n195), .IN1(r854_n194), .IN2(r854_n197) );
  AND2X1 r854_U207 ( .IN1(r854_n194), .IN2(r854_n197), .Q(r854_n196) );
  NOR2X0 r854_U206 ( .QN(P2_N4294), .IN1(r854_n195), .IN2(r854_n196) );
  NAND2X0 r854_U205 ( .IN1(P2_N5087), .IN2(r854_n194), .QN(r854_n191) );
  OR2X1 r854_U204 ( .IN2(P2_N5087), .IN1(r854_n194), .Q(r854_n193) );
  NAND2X0 r854_U203 ( .IN1(P2_N4113), .IN2(r854_n193), .QN(r854_n192) );
  NAND2X0 r854_U202 ( .IN1(r854_n191), .IN2(r854_n192), .QN(r854_n184) );
  OR2X1 r854_U200 ( .IN2(P2_N4114), .IN1(n7195), .Q(r854_n188) );
  NAND2X0 r854_U199 ( .IN1(P2_N4114), .IN2(n7195), .QN(r854_n189) );
  NAND2X0 r854_U198 ( .IN1(r854_n188), .IN2(r854_n189), .QN(r854_n187) );
  NOR2X0 r854_U197 ( .QN(r854_n185), .IN1(r854_n184), .IN2(r854_n187) );
  AND2X1 r854_U196 ( .IN1(r854_n184), .IN2(r854_n187), .Q(r854_n186) );
  NOR2X0 r854_U195 ( .QN(P2_N4295), .IN1(r854_n185), .IN2(r854_n186) );
  NAND2X0 r854_U194 ( .IN1(n7194), .IN2(r854_n184), .QN(r854_n181) );
  OR2X1 r854_U319 ( .IN2(P2_N4097), .IN1(n2919), .Q(r854_n288) );
  NAND2X0 r854_U318 ( .IN1(P2_N4097), .IN2(n2919), .QN(r854_n289) );
  NAND2X0 r854_U317 ( .IN1(r854_n288), .IN2(r854_n289), .QN(P2_N4278) );
  NAND2X0 r854_U315 ( .IN1(P2_N4097), .IN2(n7035), .QN(r854_n161) );
  OR2X1 r854_U314 ( .IN2(r854_n161), .IN1(n7186), .Q(r854_n285) );
  NAND2X0 r854_U313 ( .IN1(n7186), .IN2(r854_n161), .QN(r854_n287) );
  NAND2X0 r854_U312 ( .IN1(P2_N4098), .IN2(r854_n287), .QN(r854_n286) );
  NAND2X0 r854_U311 ( .IN1(r854_n285), .IN2(r854_n286), .QN(r854_n52) );
  NAND2X0 r854_U310 ( .IN1(n7181), .IN2(r854_n52), .QN(r854_n282) );
  OR2X1 r854_U309 ( .IN2(n7181), .IN1(r854_n52), .Q(r854_n284) );
  NAND2X0 r854_U308 ( .IN1(P2_N4099), .IN2(r854_n284), .QN(r854_n283) );
  NAND2X0 r854_U307 ( .IN1(r854_n282), .IN2(r854_n283), .QN(r854_n45) );
  NAND2X0 r854_U306 ( .IN1(n7177), .IN2(r854_n45), .QN(r854_n279) );
  OR2X1 r854_U305 ( .IN2(n7177), .IN1(r854_n45), .Q(r854_n281) );
  NAND2X0 r854_U304 ( .IN1(P2_N4100), .IN2(r854_n281), .QN(r854_n280) );
  NAND2X0 r854_U303 ( .IN1(r854_n279), .IN2(r854_n280), .QN(r854_n38) );
  NAND2X0 r854_U302 ( .IN1(n7173), .IN2(r854_n38), .QN(r854_n276) );
  OR2X1 r854_U301 ( .IN2(n7173), .IN1(r854_n38), .Q(r854_n278) );
  NAND2X0 r854_U300 ( .IN1(P2_N4101), .IN2(r854_n278), .QN(r854_n277) );
  NAND2X0 r854_U299 ( .IN1(r854_n276), .IN2(r854_n277), .QN(r854_n31) );
  NAND2X0 r854_U298 ( .IN1(n7165), .IN2(r854_n31), .QN(r854_n273) );
  OR2X1 r854_U297 ( .IN2(n7165), .IN1(r854_n31), .Q(r854_n275) );
  NAND2X0 r854_U296 ( .IN1(P2_N4102), .IN2(r854_n275), .QN(r854_n274) );
  NAND2X0 r854_U295 ( .IN1(r854_n273), .IN2(r854_n274), .QN(r854_n24) );
  NAND2X0 r854_U294 ( .IN1(P2_N5077), .IN2(r854_n24), .QN(r854_n270) );
  OR2X1 r854_U293 ( .IN2(P2_N5077), .IN1(r854_n24), .Q(r854_n272) );
  NAND2X0 r854_U292 ( .IN1(P2_N4103), .IN2(r854_n272), .QN(r854_n271) );
  NAND2X0 r854_U291 ( .IN1(r854_n270), .IN2(r854_n271), .QN(r854_n17) );
  NAND2X0 r854_U290 ( .IN1(P2_N5078), .IN2(r854_n17), .QN(r854_n267) );
  OR2X1 r854_U289 ( .IN2(P2_N5078), .IN1(r854_n17), .Q(r854_n269) );
  NAND2X0 r854_U288 ( .IN1(P2_N4104), .IN2(r854_n269), .QN(r854_n268) );
  NAND2X0 r854_U287 ( .IN1(r854_n267), .IN2(r854_n268), .QN(r854_n10) );
  OR2X1 r855_U69 ( .IN2(r855_n58), .IN1(n7243), .Q(r855_n62) );
  OR2X1 r855_U68 ( .IN2(n7238), .IN1(r855_n62), .Q(r855_n60) );
  NAND2X0 r855_U67 ( .IN1(n7238), .IN2(r855_n62), .QN(r855_n61) );
  NAND2X0 r855_U66 ( .IN1(r855_n60), .IN2(r855_n61), .QN(P2_N4454) );
  NOR2X0 r855_U65 ( .QN(r855_n57), .IN1(r855_n58), .IN2(n7243) );
  NAND2X0 r855_U64 ( .IN1(r855_n57), .IN2(n7238), .QN(r855_n50) );
  OR2X1 r855_U63 ( .IN2(P2_N5096), .IN1(r855_n50), .Q(r855_n55) );
  NAND2X0 r855_U62 ( .IN1(P2_N5096), .IN2(r855_n50), .QN(r855_n56) );
  NAND2X0 r855_U61 ( .IN1(r855_n55), .IN2(r855_n56), .QN(P2_N4455) );
  OR2X1 r855_U59 ( .IN2(r855_n50), .IN1(n7234), .Q(r855_n54) );
  OR2X1 r855_U58 ( .IN2(P2_N5097), .IN1(r855_n54), .Q(r855_n52) );
  NAND2X0 r855_U57 ( .IN1(P2_N5097), .IN2(r855_n54), .QN(r855_n53) );
  NAND2X0 r855_U56 ( .IN1(r855_n52), .IN2(r855_n53), .QN(P2_N4456) );
  NOR2X0 r855_U55 ( .QN(r855_n49), .IN1(r855_n50), .IN2(n7234) );
  NAND2X0 r855_U54 ( .IN1(r855_n49), .IN2(P2_N5097), .QN(r855_n42) );
  OR2X1 r855_U53 ( .IN2(n7227), .IN1(r855_n42), .Q(r855_n47) );
  NAND2X0 r855_U52 ( .IN1(n7227), .IN2(r855_n42), .QN(r855_n48) );
  NAND2X0 r855_U51 ( .IN1(r855_n47), .IN2(r855_n48), .QN(P2_N4457) );
  OR2X1 r855_U49 ( .IN2(r855_n42), .IN1(n7224), .Q(r855_n46) );
  OR2X1 r855_U48 ( .IN2(P2_N5099), .IN1(r855_n46), .Q(r855_n44) );
  NAND2X0 r855_U47 ( .IN1(P2_N5099), .IN2(r855_n46), .QN(r855_n45) );
  NAND2X0 r855_U46 ( .IN1(r855_n44), .IN2(r855_n45), .QN(P2_N4458) );
  NOR2X0 r855_U45 ( .QN(r855_n41), .IN1(r855_n42), .IN2(n7224) );
  NAND2X0 r855_U44 ( .IN1(r855_n41), .IN2(P2_N5099), .QN(r855_n32) );
  OR2X1 r855_U43 ( .IN2(P2_N5100), .IN1(r855_n32), .Q(r855_n39) );
  NAND2X0 r855_U42 ( .IN1(P2_N5100), .IN2(r855_n32), .QN(r855_n40) );
  NAND2X0 r855_U41 ( .IN1(r855_n39), .IN2(r855_n40), .QN(P2_N4459) );
  OR2X1 r855_U39 ( .IN2(r855_n32), .IN1(n7266), .Q(r855_n38) );
  OR2X1 r855_U38 ( .IN2(P2_N497), .IN1(r855_n38), .Q(r855_n36) );
  NAND2X0 r855_U37 ( .IN1(P2_N497), .IN2(r855_n38), .QN(r855_n37) );
  NAND2X0 r855_U36 ( .IN1(r855_n36), .IN2(r855_n37), .QN(P2_N4460) );
  OR2X1 r855_U35 ( .IN2(n7177), .IN1(r855_n26), .Q(r855_n34) );
  NAND2X0 r855_U34 ( .IN1(n7177), .IN2(r855_n26), .QN(r855_n35) );
  NAND2X0 r855_U33 ( .IN1(r855_n34), .IN2(r855_n35), .QN(P2_N4433) );
  NOR2X0 r855_U31 ( .QN(r855_n31), .IN1(r855_n32), .IN2(n7266) );
  AND2X1 r855_U30 ( .IN1(r855_n31), .IN2(P2_N497), .Q(r855_n29) );
  NOR2X0 r855_U29 ( .QN(P2_N4462), .IN1(n2562), .IN2(r855_n29) );
  INVX0 r855_U28 ( .ZN(r855_n27), .INP(P2_N4462) );
  NAND2X0 r855_U27 ( .IN1(r855_n29), .IN2(n2562), .QN(r855_n28) );
  NAND2X0 r855_U26 ( .IN1(r855_n27), .IN2(r855_n28), .QN(P2_N4461) );
  OR2X1 r855_U25 ( .IN2(r855_n26), .IN1(n7178), .Q(r855_n24) );
  OR2X1 r855_U24 ( .IN2(P2_N5075), .IN1(r855_n24), .Q(r855_n22) );
  NAND2X0 r855_U23 ( .IN1(P2_N5075), .IN2(r855_n24), .QN(r855_n23) );
  NAND2X0 r855_U22 ( .IN1(r855_n22), .IN2(r855_n23), .QN(P2_N4434) );
  OR2X1 r855_U21 ( .IN2(P2_N5076), .IN1(r855_n19), .Q(r855_n20) );
  NAND2X0 r855_U20 ( .IN1(P2_N5076), .IN2(r855_n19), .QN(r855_n21) );
  NAND2X0 r855_U19 ( .IN1(r855_n20), .IN2(r855_n21), .QN(P2_N4435) );
  OR2X1 r855_U18 ( .IN2(r855_n19), .IN1(r855_n51), .Q(r855_n17) );
  OR2X1 r855_U17 ( .IN2(n7162), .IN1(r855_n17), .Q(r855_n15) );
  NAND2X0 r855_U16 ( .IN1(n7162), .IN2(r855_n17), .QN(r855_n16) );
  NAND2X0 r855_U15 ( .IN1(r855_n15), .IN2(r855_n16), .QN(P2_N4436) );
  OR2X1 r855_U14 ( .IN2(n7158), .IN1(r855_n12), .Q(r855_n13) );
  NAND2X0 r855_U13 ( .IN1(n7158), .IN2(r855_n12), .QN(r855_n14) );
  NAND2X0 r855_U12 ( .IN1(r855_n13), .IN2(r855_n14), .QN(P2_N4437) );
  OR2X1 r855_U11 ( .IN2(r855_n12), .IN1(r855_n30), .Q(r855_n10) );
  OR2X1 r855_U10 ( .IN2(n7154), .IN1(r855_n10), .Q(r855_n8) );
  NAND2X0 r855_U9 ( .IN1(n7154), .IN2(r855_n10), .QN(r855_n9) );
  NAND2X0 r855_U8 ( .IN1(r855_n8), .IN2(r855_n9), .QN(P2_N4438) );
  OR2X1 r855_U7 ( .IN2(P2_N5080), .IN1(r855_n5), .Q(r855_n6) );
  NAND2X0 r855_U6 ( .IN1(P2_N5080), .IN2(r855_n5), .QN(r855_n7) );
  NAND2X0 r855_U5 ( .IN1(r855_n6), .IN2(r855_n7), .QN(P2_N4439) );
  OR2X1 r855_U4 ( .IN2(r855_n5), .IN1(r855_n11), .Q(r855_n3) );
  OR2X1 r855_U3 ( .IN2(n7220), .IN1(r855_n3), .Q(r855_n1) );
  NAND2X0 r855_U2 ( .IN1(n7220), .IN2(r855_n3), .QN(r855_n2) );
  NAND2X0 r855_U1 ( .IN1(r855_n1), .IN2(r855_n2), .QN(P2_N4440) );
  NAND2X0 r855_U155 ( .IN1(P2_N4430), .IN2(n7186), .QN(r855_n123) );
  INVX0 r855_U154 ( .ZN(r855_n121), .INP(P2_N4430) );
  NAND2X0 r855_U153 ( .IN1(P2_N5072), .IN2(r855_n121), .QN(r855_n124) );
  NAND2X0 r855_U152 ( .IN1(r855_n123), .IN2(r855_n124), .QN(P2_N4431) );
  NOR2X0 r855_U151 ( .QN(r855_n120), .IN1(r855_n121), .IN2(n7186) );
  NAND2X0 r855_U150 ( .IN1(r855_n120), .IN2(n7181), .QN(r855_n26) );
  NOR2X0 r855_U148 ( .QN(r855_n119), .IN1(r855_n26), .IN2(n7178) );
  NAND2X0 r855_U147 ( .IN1(r855_n119), .IN2(P2_N5075), .QN(r855_n19) );
  NOR2X0 r855_U145 ( .QN(r855_n118), .IN1(r855_n19), .IN2(r855_n51) );
  NAND2X0 r855_U144 ( .IN1(r855_n118), .IN2(n7162), .QN(r855_n12) );
  NOR2X0 r855_U142 ( .QN(r855_n117), .IN1(r855_n12), .IN2(r855_n30) );
  NAND2X0 r855_U141 ( .IN1(r855_n117), .IN2(n7154), .QN(r855_n5) );
  NOR2X0 r855_U139 ( .QN(r855_n116), .IN1(r855_n5), .IN2(r855_n11) );
  NAND2X0 r855_U138 ( .IN1(r855_n116), .IN2(n7220), .QN(r855_n109) );
  OR2X1 r855_U137 ( .IN2(n7216), .IN1(r855_n109), .Q(r855_n114) );
  NAND2X0 r855_U136 ( .IN1(n7216), .IN2(r855_n109), .QN(r855_n115) );
  NAND2X0 r855_U135 ( .IN1(r855_n114), .IN2(r855_n115), .QN(P2_N4441) );
  OR2X1 r855_U133 ( .IN2(r855_n109), .IN1(r855_n134), .Q(r855_n113) );
  OR2X1 r855_U132 ( .IN2(P2_N5083), .IN1(r855_n113), .Q(r855_n111) );
  NAND2X0 r855_U131 ( .IN1(P2_N5083), .IN2(r855_n113), .QN(r855_n112) );
  NAND2X0 r855_U130 ( .IN1(r855_n111), .IN2(r855_n112), .QN(P2_N4442) );
  NOR2X0 r855_U129 ( .QN(r855_n108), .IN1(r855_n109), .IN2(r855_n134) );
  NAND2X0 r855_U128 ( .IN1(r855_n108), .IN2(P2_N5083), .QN(r855_n101) );
  OR2X1 r855_U127 ( .IN2(n7209), .IN1(r855_n101), .Q(r855_n106) );
  NAND2X0 r855_U126 ( .IN1(n7209), .IN2(r855_n101), .QN(r855_n107) );
  NAND2X0 r855_U125 ( .IN1(r855_n106), .IN2(r855_n107), .QN(P2_N4443) );
  OR2X1 r855_U123 ( .IN2(r855_n101), .IN1(r855_n131), .Q(r855_n105) );
  OR2X1 r855_U122 ( .IN2(n7206), .IN1(r855_n105), .Q(r855_n103) );
  NAND2X0 r855_U121 ( .IN1(n7206), .IN2(r855_n105), .QN(r855_n104) );
  NAND2X0 r855_U120 ( .IN1(r855_n103), .IN2(r855_n104), .QN(P2_N4444) );
  NOR2X0 r855_U119 ( .QN(r855_n100), .IN1(r855_n101), .IN2(r855_n131) );
  NAND2X0 r855_U118 ( .IN1(r855_n100), .IN2(n7206), .QN(r855_n93) );
  OR2X1 r855_U117 ( .IN2(n7202), .IN1(r855_n93), .Q(r855_n98) );
  NAND2X0 r855_U116 ( .IN1(n7202), .IN2(r855_n93), .QN(r855_n99) );
  NAND2X0 r855_U115 ( .IN1(r855_n98), .IN2(r855_n99), .QN(P2_N4445) );
  OR2X1 r855_U113 ( .IN2(r855_n93), .IN1(r855_n128), .Q(r855_n97) );
  OR2X1 r855_U112 ( .IN2(n7198), .IN1(r855_n97), .Q(r855_n95) );
  NAND2X0 r855_U111 ( .IN1(n7198), .IN2(r855_n97), .QN(r855_n96) );
  NAND2X0 r855_U110 ( .IN1(r855_n95), .IN2(r855_n96), .QN(P2_N4446) );
  NOR2X0 r855_U109 ( .QN(r855_n92), .IN1(r855_n93), .IN2(r855_n128) );
  NAND2X0 r855_U108 ( .IN1(r855_n92), .IN2(n7198), .QN(r855_n85) );
  OR2X1 r855_U107 ( .IN2(P2_N5088), .IN1(r855_n85), .Q(r855_n90) );
  NAND2X0 r855_U106 ( .IN1(P2_N5088), .IN2(r855_n85), .QN(r855_n91) );
  NAND2X0 r855_U105 ( .IN1(r855_n90), .IN2(r855_n91), .QN(P2_N4447) );
  OR2X1 r855_U103 ( .IN2(r855_n85), .IN1(r855_n125), .Q(r855_n89) );
  OR2X1 r855_U102 ( .IN2(P2_N5089), .IN1(r855_n89), .Q(r855_n87) );
  NAND2X0 r855_U101 ( .IN1(P2_N5089), .IN2(r855_n89), .QN(r855_n88) );
  NAND2X0 r855_U100 ( .IN1(r855_n87), .IN2(r855_n88), .QN(P2_N4448) );
  NOR2X0 r855_U99 ( .QN(r855_n84), .IN1(r855_n85), .IN2(r855_n125) );
  NAND2X0 r855_U98 ( .IN1(r855_n84), .IN2(P2_N5089), .QN(r855_n74) );
  OR2X1 r855_U97 ( .IN2(n7263), .IN1(r855_n74), .Q(r855_n82) );
  NAND2X0 r855_U96 ( .IN1(n7263), .IN2(r855_n74), .QN(r855_n83) );
  NAND2X0 r855_U95 ( .IN1(r855_n82), .IN2(r855_n83), .QN(P2_N4449) );
  OR2X1 r855_U93 ( .IN2(r855_n74), .IN1(n7264), .Q(r855_n81) );
  OR2X1 r855_U92 ( .IN2(n7259), .IN1(r855_n81), .Q(r855_n79) );
  NAND2X0 r855_U91 ( .IN1(n7259), .IN2(r855_n81), .QN(r855_n80) );
  NAND2X0 r855_U90 ( .IN1(r855_n79), .IN2(r855_n80), .QN(P2_N4450) );
  NAND2X0 r855_U89 ( .IN1(P2_N5072), .IN2(P2_N4430), .QN(r855_n78) );
  OR2X1 r855_U88 ( .IN2(n7181), .IN1(r855_n78), .Q(r855_n76) );
  NAND2X0 r855_U87 ( .IN1(n7181), .IN2(r855_n78), .QN(r855_n77) );
  NAND2X0 r855_U86 ( .IN1(r855_n76), .IN2(r855_n77), .QN(P2_N4432) );
  NOR2X0 r855_U85 ( .QN(r855_n73), .IN1(r855_n74), .IN2(n7264) );
  NAND2X0 r855_U84 ( .IN1(r855_n73), .IN2(n7259), .QN(r855_n66) );
  OR2X1 r855_U83 ( .IN2(P2_N5092), .IN1(r855_n66), .Q(r855_n71) );
  NAND2X0 r855_U82 ( .IN1(P2_N5092), .IN2(r855_n66), .QN(r855_n72) );
  NAND2X0 r855_U81 ( .IN1(r855_n71), .IN2(r855_n72), .QN(P2_N4451) );
  OR2X1 r855_U79 ( .IN2(r855_n66), .IN1(r855_n146), .Q(r855_n70) );
  OR2X1 r855_U78 ( .IN2(P2_N5093), .IN1(r855_n70), .Q(r855_n68) );
  NAND2X0 r855_U77 ( .IN1(P2_N5093), .IN2(r855_n70), .QN(r855_n69) );
  NAND2X0 r855_U76 ( .IN1(r855_n68), .IN2(r855_n69), .QN(P2_N4452) );
  NOR2X0 r855_U75 ( .QN(r855_n65), .IN1(r855_n66), .IN2(r855_n146) );
  NAND2X0 r855_U74 ( .IN1(r855_n65), .IN2(P2_N5093), .QN(r855_n58) );
  OR2X1 r855_U73 ( .IN2(P2_N5094), .IN1(r855_n58), .Q(r855_n63) );
  NAND2X0 r855_U72 ( .IN1(P2_N5094), .IN2(r855_n58), .QN(r855_n64) );
  NAND2X0 r855_U71 ( .IN1(r855_n63), .IN2(r855_n64), .QN(P2_N4453) );
  INVX0 r855_U32 ( .ZN(r855_n11), .INP(P2_N5080) );
  INVX0 r855_U40 ( .ZN(r855_n30), .INP(n7158) );
  INVX0 r855_U50 ( .ZN(r855_n51), .INP(P2_N5076) );
  INVX0 r855_U60 ( .ZN(r855_n125), .INP(P2_N5088) );
  INVX0 r855_U70 ( .ZN(r855_n128), .INP(n7202) );
  INVX0 r855_U80 ( .ZN(r855_n131), .INP(n7209) );
  INVX0 r855_U94 ( .ZN(r855_n134), .INP(n7216) );
  INVX0 r855_U104 ( .ZN(r855_n146), .INP(P2_N5092) );
  NAND2X0 r860_U59 ( .IN1(r860_n108), .IN2(r860_n109), .QN(r860_n107) );
  NOR2X0 r860_U58 ( .QN(r860_n101), .IN1(r860_n106), .IN2(r860_n107) );
  INVX0 r860_U57 ( .ZN(r860_n103), .INP(r860_n105) );
  NAND2X0 r860_U56 ( .IN1(r860_n103), .IN2(r860_n104), .QN(r860_n102) );
  NOR2X0 r860_U55 ( .QN(r860_n100), .IN1(r860_n101), .IN2(r860_n102) );
  NOR2X0 r860_U54 ( .QN(r860_n97), .IN1(r860_n99), .IN2(r860_n100) );
  NAND2X0 r860_U53 ( .IN1(r860_n97), .IN2(r860_n98), .QN(r860_n96) );
  NAND2X0 r860_U52 ( .IN1(r860_n95), .IN2(r860_n96), .QN(r860_n93) );
  NAND2X0 r860_U51 ( .IN1(r860_n93), .IN2(r860_n94), .QN(r860_n92) );
  NOR2X0 r860_U50 ( .QN(r860_n86), .IN1(r860_n91), .IN2(r860_n92) );
  INVX0 r860_U49 ( .ZN(r860_n88), .INP(r860_n90) );
  NAND2X0 r860_U48 ( .IN1(r860_n88), .IN2(r860_n89), .QN(r860_n87) );
  NOR2X0 r860_U47 ( .QN(r860_n85), .IN1(r860_n86), .IN2(r860_n87) );
  NOR2X0 r860_U46 ( .QN(r860_n82), .IN1(r860_n84), .IN2(r860_n85) );
  NAND2X0 r860_U45 ( .IN1(r860_n82), .IN2(r860_n83), .QN(r860_n81) );
  NAND2X0 r860_U44 ( .IN1(r860_n80), .IN2(r860_n81), .QN(r860_n78) );
  NAND2X0 r860_U43 ( .IN1(r860_n78), .IN2(r860_n79), .QN(r860_n77) );
  NOR2X0 r860_U42 ( .QN(r860_n71), .IN1(r860_n76), .IN2(r860_n77) );
  INVX0 r860_U41 ( .ZN(r860_n73), .INP(r860_n75) );
  NAND2X0 r860_U40 ( .IN1(r860_n73), .IN2(r860_n74), .QN(r860_n72) );
  NOR2X0 r860_U39 ( .QN(r860_n70), .IN1(r860_n71), .IN2(r860_n72) );
  NOR2X0 r860_U38 ( .QN(r860_n67), .IN1(r860_n69), .IN2(r860_n70) );
  NAND2X0 r860_U37 ( .IN1(r860_n67), .IN2(r860_n68), .QN(r860_n66) );
  NAND2X0 r860_U36 ( .IN1(r860_n65), .IN2(r860_n66), .QN(r860_n63) );
  NAND2X0 r860_U35 ( .IN1(r860_n63), .IN2(r860_n64), .QN(r860_n62) );
  NOR2X0 r860_U34 ( .QN(r860_n56), .IN1(r860_n61), .IN2(r860_n62) );
  INVX0 r860_U33 ( .ZN(r860_n58), .INP(r860_n60) );
  NAND2X0 r860_U32 ( .IN1(r860_n58), .IN2(r860_n59), .QN(r860_n57) );
  NOR2X0 r860_U31 ( .QN(r860_n55), .IN1(r860_n56), .IN2(r860_n57) );
  NOR2X0 r860_U30 ( .QN(r860_n52), .IN1(r860_n54), .IN2(r860_n55) );
  NAND2X0 r860_U29 ( .IN1(r860_n52), .IN2(r860_n53), .QN(r860_n51) );
  NAND2X0 r860_U28 ( .IN1(r860_n50), .IN2(r860_n51), .QN(r860_n48) );
  NAND2X0 r860_U27 ( .IN1(r860_n48), .IN2(r860_n49), .QN(r860_n47) );
  NOR2X0 r860_U26 ( .QN(r860_n41), .IN1(r860_n46), .IN2(r860_n47) );
  INVX0 r860_U25 ( .ZN(r860_n43), .INP(r860_n45) );
  NAND2X0 r860_U24 ( .IN1(r860_n43), .IN2(r860_n44), .QN(r860_n42) );
  NOR2X0 r860_U23 ( .QN(r860_n40), .IN1(r860_n41), .IN2(r860_n42) );
  NOR2X0 r860_U22 ( .QN(r860_n37), .IN1(r860_n39), .IN2(r860_n40) );
  NAND2X0 r860_U21 ( .IN1(r860_n37), .IN2(r860_n38), .QN(r860_n36) );
  NAND2X0 r860_U20 ( .IN1(r860_n35), .IN2(r860_n36), .QN(r860_n33) );
  NAND2X0 r860_U19 ( .IN1(r860_n33), .IN2(r860_n34), .QN(r860_n32) );
  NOR2X0 r860_U18 ( .QN(r860_n26), .IN1(r860_n31), .IN2(r860_n32) );
  INVX0 r860_U17 ( .ZN(r860_n28), .INP(r860_n30) );
  NAND2X0 r860_U16 ( .IN1(r860_n28), .IN2(r860_n29), .QN(r860_n27) );
  NOR2X0 r860_U15 ( .QN(r860_n25), .IN1(r860_n26), .IN2(r860_n27) );
  NOR2X0 r860_U14 ( .QN(r860_n22), .IN1(r860_n24), .IN2(r860_n25) );
  NAND2X0 r860_U13 ( .IN1(r860_n22), .IN2(r860_n23), .QN(r860_n21) );
  NAND2X0 r860_U12 ( .IN1(r860_n20), .IN2(r860_n21), .QN(r860_n18) );
  NAND2X0 r860_U11 ( .IN1(r860_n18), .IN2(r860_n19), .QN(r860_n17) );
  NOR2X0 r860_U10 ( .QN(r860_n11), .IN1(r860_n16), .IN2(r860_n17) );
  INVX0 r860_U9 ( .ZN(r860_n13), .INP(r860_n15) );
  NAND2X0 r860_U8 ( .IN1(r860_n13), .IN2(r860_n14), .QN(r860_n12) );
  NOR2X0 r860_U7 ( .QN(r860_n10), .IN1(r860_n11), .IN2(r860_n12) );
  NOR2X0 r860_U6 ( .QN(r860_n7), .IN1(r860_n9), .IN2(r860_n10) );
  NAND2X0 r860_U5 ( .IN1(r860_n7), .IN2(r860_n8), .QN(r860_n5) );
  NAND2X0 r860_U4 ( .IN1(r860_n5), .IN2(r860_n6), .QN(r860_n3) );
  NAND2X0 r860_U3 ( .IN1(r860_n3), .IN2(r860_n4), .QN(r860_n2) );
  NAND2X0 r860_U2 ( .IN1(r860_n1), .IN2(r860_n2), .QN(P2_N5065) );
  NOR2X0 r860_U1 ( .QN(P2_N5062), .IN1(P2_N5059), .IN2(P2_N5065) );
  NOR2X0 r860_U152 ( .QN(r860_n68), .IN1(r860_n127), .IN2(r860_n201) );
  NAND2X0 r860_U151 ( .IN1(r860_n200), .IN2(r860_n68), .QN(r860_n198) );
  NAND2X0 r860_U150 ( .IN1(r860_n198), .IN2(r860_n199), .QN(r860_n197) );
  NOR2X0 r860_U149 ( .QN(r860_n195), .IN1(r860_n196), .IN2(r860_n197) );
  NOR2X0 r860_U148 ( .QN(r860_n192), .IN1(r860_n128), .IN2(r860_n195) );
  OR2X1 r860_U146 ( .IN2(P2_N5022), .IN1(n7197), .Q(r860_n59) );
  NAND2X0 r860_U145 ( .IN1(P2_N5022), .IN2(n7197), .QN(r860_n191) );
  NAND2X0 r860_U144 ( .IN1(r860_n59), .IN2(r860_n191), .QN(r860_n61) );
  INVX0 r860_U143 ( .ZN(r860_n193), .INP(r860_n61) );
  NAND2X0 r860_U142 ( .IN1(r860_n192), .IN2(r860_n193), .QN(r860_n190) );
  NAND2X0 r860_U141 ( .IN1(r860_n190), .IN2(r860_n191), .QN(r860_n189) );
  NOR2X0 r860_U140 ( .QN(r860_n188), .IN1(r860_n54), .IN2(r860_n189) );
  NOR2X0 r860_U139 ( .QN(r860_n185), .IN1(r860_n60), .IN2(r860_n188) );
  NOR2X0 r860_U137 ( .QN(r860_n129), .IN1(n7188), .IN2(P2_N5024) );
  NAND2X0 r860_U136 ( .IN1(P2_N5024), .IN2(n7188), .QN(r860_n184) );
  INVX0 r860_U135 ( .ZN(r860_n186), .INP(r860_n184) );
  NOR2X0 r860_U134 ( .QN(r860_n53), .IN1(r860_n129), .IN2(r860_n186) );
  NAND2X0 r860_U133 ( .IN1(r860_n185), .IN2(r860_n53), .QN(r860_n183) );
  NAND2X0 r860_U132 ( .IN1(r860_n183), .IN2(r860_n184), .QN(r860_n182) );
  NOR2X0 r860_U131 ( .QN(r860_n180), .IN1(r860_n181), .IN2(r860_n182) );
  NOR2X0 r860_U130 ( .QN(r860_n177), .IN1(r860_n130), .IN2(r860_n180) );
  OR2X1 r860_U128 ( .IN2(P2_N5026), .IN1(n7260), .Q(r860_n44) );
  NAND2X0 r860_U127 ( .IN1(P2_N5026), .IN2(n7260), .QN(r860_n176) );
  NAND2X0 r860_U126 ( .IN1(r860_n44), .IN2(r860_n176), .QN(r860_n46) );
  INVX0 r860_U125 ( .ZN(r860_n178), .INP(r860_n46) );
  NAND2X0 r860_U124 ( .IN1(r860_n177), .IN2(r860_n178), .QN(r860_n175) );
  NAND2X0 r860_U123 ( .IN1(r860_n175), .IN2(r860_n176), .QN(r860_n174) );
  NOR2X0 r860_U122 ( .QN(r860_n173), .IN1(r860_n39), .IN2(r860_n174) );
  NOR2X0 r860_U121 ( .QN(r860_n170), .IN1(r860_n45), .IN2(r860_n173) );
  NOR2X0 r860_U119 ( .QN(r860_n131), .IN1(r860_n303), .IN2(P2_N5028) );
  NAND2X0 r860_U118 ( .IN1(P2_N5028), .IN2(r860_n303), .QN(r860_n169) );
  INVX0 r860_U117 ( .ZN(r860_n171), .INP(r860_n169) );
  NOR2X0 r860_U116 ( .QN(r860_n38), .IN1(r860_n131), .IN2(r860_n171) );
  NAND2X0 r860_U115 ( .IN1(r860_n170), .IN2(r860_n38), .QN(r860_n168) );
  NAND2X0 r860_U114 ( .IN1(r860_n168), .IN2(r860_n169), .QN(r860_n167) );
  NOR2X0 r860_U113 ( .QN(r860_n165), .IN1(r860_n166), .IN2(r860_n167) );
  NOR2X0 r860_U112 ( .QN(r860_n162), .IN1(r860_n132), .IN2(r860_n165) );
  OR2X1 r860_U110 ( .IN2(P2_N5030), .IN1(r860_n300), .Q(r860_n29) );
  NAND2X0 r860_U109 ( .IN1(P2_N5030), .IN2(r860_n300), .QN(r860_n161) );
  NAND2X0 r860_U108 ( .IN1(r860_n29), .IN2(r860_n161), .QN(r860_n31) );
  INVX0 r860_U107 ( .ZN(r860_n163), .INP(r860_n31) );
  NAND2X0 r860_U106 ( .IN1(r860_n162), .IN2(r860_n163), .QN(r860_n160) );
  NAND2X0 r860_U105 ( .IN1(r860_n160), .IN2(r860_n161), .QN(r860_n159) );
  NOR2X0 r860_U104 ( .QN(r860_n158), .IN1(r860_n24), .IN2(r860_n159) );
  NOR2X0 r860_U103 ( .QN(r860_n155), .IN1(r860_n30), .IN2(r860_n158) );
  NOR2X0 r860_U101 ( .QN(r860_n133), .IN1(r860_n297), .IN2(P2_N5032) );
  NAND2X0 r860_U100 ( .IN1(P2_N5032), .IN2(r860_n297), .QN(r860_n154) );
  INVX0 r860_U99 ( .ZN(r860_n156), .INP(r860_n154) );
  NOR2X0 r860_U98 ( .QN(r860_n23), .IN1(r860_n133), .IN2(r860_n156) );
  NAND2X0 r860_U97 ( .IN1(r860_n155), .IN2(r860_n23), .QN(r860_n153) );
  NAND2X0 r860_U96 ( .IN1(r860_n153), .IN2(r860_n154), .QN(r860_n152) );
  NOR2X0 r860_U95 ( .QN(r860_n150), .IN1(r860_n151), .IN2(r860_n152) );
  NOR2X0 r860_U94 ( .QN(r860_n147), .IN1(r860_n134), .IN2(r860_n150) );
  OR2X1 r860_U92 ( .IN2(P2_N5034), .IN1(n7222), .Q(r860_n14) );
  NAND2X0 r860_U91 ( .IN1(P2_N5034), .IN2(n7222), .QN(r860_n146) );
  NAND2X0 r860_U90 ( .IN1(r860_n14), .IN2(r860_n146), .QN(r860_n16) );
  INVX0 r860_U89 ( .ZN(r860_n148), .INP(r860_n16) );
  NAND2X0 r860_U88 ( .IN1(r860_n147), .IN2(r860_n148), .QN(r860_n145) );
  NAND2X0 r860_U87 ( .IN1(r860_n145), .IN2(r860_n146), .QN(r860_n144) );
  NOR2X0 r860_U86 ( .QN(r860_n143), .IN1(r860_n9), .IN2(r860_n144) );
  NOR2X0 r860_U85 ( .QN(r860_n140), .IN1(r860_n15), .IN2(r860_n143) );
  NAND2X0 r860_U83 ( .IN1(P2_N497), .IN2(r860_n309), .QN(r860_n6) );
  NAND2X0 r860_U81 ( .IN1(P2_N5036), .IN2(n7265), .QN(r860_n139) );
  AND2X1 r860_U80 ( .IN1(r860_n6), .IN2(r860_n139), .Q(r860_n8) );
  NAND2X0 r860_U79 ( .IN1(r860_n140), .IN2(r860_n8), .QN(r860_n138) );
  NAND2X0 r860_U78 ( .IN1(r860_n138), .IN2(r860_n139), .QN(r860_n136) );
  NAND2X0 r860_U77 ( .IN1(P2_N5037), .IN2(n2562), .QN(r860_n1) );
  NAND2X0 r860_U76 ( .IN1(r860_n136), .IN2(r860_n1), .QN(r860_n135) );
  NAND2X0 r860_U75 ( .IN1(r860_n4), .IN2(r860_n135), .QN(P2_N5059) );
  NOR2X0 r860_U74 ( .QN(r860_n20), .IN1(r860_n133), .IN2(r860_n134) );
  NOR2X0 r860_U73 ( .QN(r860_n35), .IN1(r860_n131), .IN2(r860_n132) );
  NOR2X0 r860_U72 ( .QN(r860_n50), .IN1(r860_n129), .IN2(r860_n130) );
  NOR2X0 r860_U71 ( .QN(r860_n65), .IN1(r860_n127), .IN2(r860_n128) );
  NOR2X0 r860_U70 ( .QN(r860_n80), .IN1(r860_n125), .IN2(r860_n126) );
  NOR2X0 r860_U69 ( .QN(r860_n95), .IN1(r860_n123), .IN2(r860_n124) );
  NOR2X0 r860_U68 ( .QN(r860_n110), .IN1(r860_n121), .IN2(r860_n122) );
  NAND2X0 r860_U67 ( .IN1(n7035), .IN2(r860_n120), .QN(r860_n117) );
  NOR2X0 r860_U66 ( .QN(r860_n118), .IN1(n7184), .IN2(r860_n117) );
  INVX0 r860_U65 ( .ZN(r860_n119), .INP(P2_N5007) );
  NOR2X0 r860_U64 ( .QN(r860_n114), .IN1(r860_n118), .IN2(r860_n119) );
  AND2X1 r860_U63 ( .IN1(n7184), .IN2(r860_n117), .Q(r860_n115) );
  NOR2X0 r860_U62 ( .QN(r860_n112), .IN1(r860_n114), .IN2(r860_n115) );
  NAND2X0 r860_U61 ( .IN1(r860_n112), .IN2(r860_n113), .QN(r860_n111) );
  NAND2X0 r860_U60 ( .IN1(r860_n110), .IN2(r860_n111), .QN(r860_n108) );
  NOR2X0 r860_U244 ( .QN(r860_n60), .IN1(n7195), .IN2(P2_N5023) );
  AND2X1 r860_U243 ( .IN1(P2_N5023), .IN2(n7195), .Q(r860_n54) );
  NOR2X0 r860_U241 ( .QN(r860_n128), .IN1(n7201), .IN2(P2_N5021) );
  NAND2X0 r860_U240 ( .IN1(P2_N5021), .IN2(n7201), .QN(r860_n64) );
  INVX0 r860_U239 ( .ZN(r860_n196), .INP(r860_n64) );
  NOR2X0 r860_U237 ( .QN(r860_n75), .IN1(n7208), .IN2(P2_N5019) );
  AND2X1 r860_U236 ( .IN1(P2_N5019), .IN2(n7208), .Q(r860_n69) );
  NOR2X0 r860_U234 ( .QN(r860_n126), .IN1(n7214), .IN2(P2_N5017) );
  NAND2X0 r860_U233 ( .IN1(P2_N5017), .IN2(n7214), .QN(r860_n79) );
  INVX0 r860_U232 ( .ZN(r860_n211), .INP(r860_n79) );
  NOR2X0 r860_U230 ( .QN(r860_n90), .IN1(n7149), .IN2(P2_N5015) );
  AND2X1 r860_U229 ( .IN1(P2_N5015), .IN2(n7149), .Q(r860_n84) );
  NOR2X0 r860_U227 ( .QN(r860_n124), .IN1(n7157), .IN2(P2_N5013) );
  NAND2X0 r860_U226 ( .IN1(P2_N5013), .IN2(n7157), .QN(r860_n94) );
  INVX0 r860_U225 ( .ZN(r860_n226), .INP(r860_n94) );
  NOR2X0 r860_U223 ( .QN(r860_n105), .IN1(n7166), .IN2(P2_N5011) );
  AND2X1 r860_U222 ( .IN1(P2_N5011), .IN2(n7166), .Q(r860_n99) );
  NOR2X0 r860_U220 ( .QN(r860_n122), .IN1(n7178), .IN2(P2_N5009) );
  NAND2X0 r860_U219 ( .IN1(P2_N5009), .IN2(n7178), .QN(r860_n109) );
  INVX0 r860_U218 ( .ZN(r860_n241), .INP(r860_n109) );
  INVX0 r860_U216 ( .ZN(r860_n120), .INP(P2_N5006) );
  NOR2X0 r860_U215 ( .QN(r860_n250), .IN1(r860_n120), .IN2(n7035) );
  AND2X1 r860_U214 ( .IN1(n7184), .IN2(r860_n250), .Q(r860_n251) );
  NOR2X0 r860_U213 ( .QN(r860_n248), .IN1(P2_N5007), .IN2(r860_n251) );
  NOR2X0 r860_U212 ( .QN(r860_n249), .IN1(r860_n250), .IN2(n7184) );
  NOR2X0 r860_U211 ( .QN(r860_n245), .IN1(r860_n248), .IN2(r860_n249) );
  NOR2X0 r860_U209 ( .QN(r860_n121), .IN1(n7182), .IN2(P2_N5008) );
  NAND2X0 r860_U208 ( .IN1(P2_N5008), .IN2(n7182), .QN(r860_n244) );
  INVX0 r860_U207 ( .ZN(r860_n246), .INP(r860_n244) );
  NOR2X0 r860_U206 ( .QN(r860_n113), .IN1(r860_n121), .IN2(r860_n246) );
  NAND2X0 r860_U205 ( .IN1(r860_n245), .IN2(r860_n113), .QN(r860_n243) );
  NAND2X0 r860_U204 ( .IN1(r860_n243), .IN2(r860_n244), .QN(r860_n242) );
  NOR2X0 r860_U203 ( .QN(r860_n240), .IN1(r860_n241), .IN2(r860_n242) );
  NOR2X0 r860_U202 ( .QN(r860_n237), .IN1(r860_n122), .IN2(r860_n240) );
  OR2X1 r860_U200 ( .IN2(P2_N5010), .IN1(n7174), .Q(r860_n104) );
  NAND2X0 r860_U199 ( .IN1(P2_N5010), .IN2(n7174), .QN(r860_n236) );
  NAND2X0 r860_U198 ( .IN1(r860_n104), .IN2(r860_n236), .QN(r860_n106) );
  INVX0 r860_U197 ( .ZN(r860_n238), .INP(r860_n106) );
  NAND2X0 r860_U196 ( .IN1(r860_n237), .IN2(r860_n238), .QN(r860_n235) );
  NAND2X0 r860_U195 ( .IN1(r860_n235), .IN2(r860_n236), .QN(r860_n234) );
  NOR2X0 r860_U194 ( .QN(r860_n233), .IN1(r860_n99), .IN2(r860_n234) );
  NOR2X0 r860_U193 ( .QN(r860_n230), .IN1(r860_n105), .IN2(r860_n233) );
  NOR2X0 r860_U191 ( .QN(r860_n123), .IN1(n7164), .IN2(P2_N5012) );
  NAND2X0 r860_U190 ( .IN1(P2_N5012), .IN2(n7164), .QN(r860_n229) );
  INVX0 r860_U189 ( .ZN(r860_n231), .INP(r860_n229) );
  NOR2X0 r860_U188 ( .QN(r860_n98), .IN1(r860_n123), .IN2(r860_n231) );
  NAND2X0 r860_U187 ( .IN1(r860_n230), .IN2(r860_n98), .QN(r860_n228) );
  NAND2X0 r860_U186 ( .IN1(r860_n228), .IN2(r860_n229), .QN(r860_n227) );
  NOR2X0 r860_U185 ( .QN(r860_n225), .IN1(r860_n226), .IN2(r860_n227) );
  NOR2X0 r860_U184 ( .QN(r860_n222), .IN1(r860_n124), .IN2(r860_n225) );
  OR2X1 r860_U182 ( .IN2(P2_N5014), .IN1(n7153), .Q(r860_n89) );
  NAND2X0 r860_U181 ( .IN1(P2_N5014), .IN2(n7153), .QN(r860_n221) );
  NAND2X0 r860_U180 ( .IN1(r860_n89), .IN2(r860_n221), .QN(r860_n91) );
  INVX0 r860_U179 ( .ZN(r860_n223), .INP(r860_n91) );
  NAND2X0 r860_U178 ( .IN1(r860_n222), .IN2(r860_n223), .QN(r860_n220) );
  NAND2X0 r860_U177 ( .IN1(r860_n220), .IN2(r860_n221), .QN(r860_n219) );
  NOR2X0 r860_U176 ( .QN(r860_n218), .IN1(r860_n84), .IN2(r860_n219) );
  NOR2X0 r860_U175 ( .QN(r860_n215), .IN1(r860_n90), .IN2(r860_n218) );
  NOR2X0 r860_U173 ( .QN(r860_n125), .IN1(n7219), .IN2(P2_N5016) );
  NAND2X0 r860_U172 ( .IN1(P2_N5016), .IN2(n7219), .QN(r860_n214) );
  INVX0 r860_U171 ( .ZN(r860_n216), .INP(r860_n214) );
  NOR2X0 r860_U170 ( .QN(r860_n83), .IN1(r860_n125), .IN2(r860_n216) );
  NAND2X0 r860_U169 ( .IN1(r860_n215), .IN2(r860_n83), .QN(r860_n213) );
  NAND2X0 r860_U168 ( .IN1(r860_n213), .IN2(r860_n214), .QN(r860_n212) );
  NOR2X0 r860_U167 ( .QN(r860_n210), .IN1(r860_n211), .IN2(r860_n212) );
  NOR2X0 r860_U166 ( .QN(r860_n207), .IN1(r860_n126), .IN2(r860_n210) );
  OR2X1 r860_U164 ( .IN2(P2_N5018), .IN1(n7211), .Q(r860_n74) );
  NAND2X0 r860_U163 ( .IN1(P2_N5018), .IN2(n7211), .QN(r860_n206) );
  NAND2X0 r860_U162 ( .IN1(r860_n74), .IN2(r860_n206), .QN(r860_n76) );
  INVX0 r860_U161 ( .ZN(r860_n208), .INP(r860_n76) );
  NAND2X0 r860_U160 ( .IN1(r860_n207), .IN2(r860_n208), .QN(r860_n205) );
  NAND2X0 r860_U159 ( .IN1(r860_n205), .IN2(r860_n206), .QN(r860_n204) );
  NOR2X0 r860_U158 ( .QN(r860_n203), .IN1(r860_n69), .IN2(r860_n204) );
  NOR2X0 r860_U157 ( .QN(r860_n200), .IN1(r860_n75), .IN2(r860_n203) );
  NOR2X0 r860_U155 ( .QN(r860_n127), .IN1(n7205), .IN2(P2_N5020) );
  NAND2X0 r860_U154 ( .IN1(P2_N5020), .IN2(n7205), .QN(r860_n199) );
  INVX0 r860_U153 ( .ZN(r860_n201), .INP(r860_n199) );
  OR2X1 r860_U267 ( .IN2(P2_N5037), .IN1(n2562), .Q(r860_n4) );
  NOR2X0 r860_U265 ( .QN(r860_n15), .IN1(n7266), .IN2(P2_N5035) );
  AND2X1 r860_U264 ( .IN1(P2_N5035), .IN2(n7266), .Q(r860_n9) );
  NOR2X0 r860_U262 ( .QN(r860_n134), .IN1(n7224), .IN2(P2_N5033) );
  NAND2X0 r860_U261 ( .IN1(P2_N5033), .IN2(n7224), .QN(r860_n19) );
  INVX0 r860_U260 ( .ZN(r860_n151), .INP(r860_n19) );
  NOR2X0 r860_U258 ( .QN(r860_n30), .IN1(n7234), .IN2(P2_N5031) );
  AND2X1 r860_U257 ( .IN1(P2_N5031), .IN2(n7234), .Q(r860_n24) );
  NOR2X0 r860_U255 ( .QN(r860_n132), .IN1(n7243), .IN2(P2_N5029) );
  NAND2X0 r860_U254 ( .IN1(P2_N5029), .IN2(n7243), .QN(r860_n34) );
  INVX0 r860_U253 ( .ZN(r860_n166), .INP(r860_n34) );
  NOR2X0 r860_U251 ( .QN(r860_n45), .IN1(n7253), .IN2(P2_N5027) );
  AND2X1 r860_U250 ( .IN1(P2_N5027), .IN2(n7253), .Q(r860_n39) );
  NOR2X0 r860_U248 ( .QN(r860_n130), .IN1(n7264), .IN2(P2_N5025) );
  NAND2X0 r860_U247 ( .IN1(P2_N5025), .IN2(n7264), .QN(r860_n49) );
  INVX0 r860_U246 ( .ZN(r860_n181), .INP(r860_n49) );
  INVX0 r860_U82 ( .ZN(r860_n297), .INP(P2_N5097) );
  INVX0 r860_U84 ( .ZN(r860_n300), .INP(P2_N5095) );
  INVX0 r860_U93 ( .ZN(r860_n303), .INP(P2_N5093) );
  INVX0 r860_U102 ( .ZN(r860_n309), .INP(P2_N5036) );
  NAND2X0 add_1095_U203 ( .IN1(add_1095_n63), .IN2(add_1095_n60), 
        .QN(add_1095_n187) );
  OR2X1 add_1095_U204 ( .IN2(add_1095_n60), .IN1(add_1095_n63), 
        .Q(add_1095_n185) );
  NAND2X0 add_1095_U205 ( .IN1(n9489), .IN2(n9329), .QN(add_1095_n60) );
  INVX0 add_1095_U206 ( .ZN(add_1095_n63), .INP(n9318) );
  NAND2X0 add_1095_U207 ( .IN1(add_1095_n188), .IN2(add_1095_n189), .QN(so_0_)
         );
  NAND2X0 add_1095_U208 ( .IN1(n9489), .IN2(add_1095_n190), .QN(add_1095_n189)
         );
  OR2X1 add_1095_U209 ( .IN2(n9489), .IN1(add_1095_n190), .Q(add_1095_n188) );
  INVX0 add_1095_U210 ( .ZN(add_1095_n190), .INP(n9329) );
  OR2X1 add_1095_U195 ( .IN2(n9625), .IN1(add_1095_n45), .Q(add_1095_n181) );
  NAND2X0 add_1095_U196 ( .IN1(n9625), .IN2(add_1095_n45), .QN(add_1095_n179)
         );
  NAND2X0 add_1095_U197 ( .IN1(add_1095_n182), .IN2(add_1095_n183), 
        .QN(add_1095_n45) );
  NAND2X0 add_1095_U198 ( .IN1(n9481), .IN2(add_1095_n184), .QN(add_1095_n183)
         );
  OR2X1 add_1095_U199 ( .IN2(n9629), .IN1(add_1095_n52), .Q(add_1095_n184) );
  NAND2X0 add_1095_U200 ( .IN1(n9629), .IN2(add_1095_n52), .QN(add_1095_n182)
         );
  NAND2X0 add_1095_U201 ( .IN1(add_1095_n185), .IN2(add_1095_n186), 
        .QN(add_1095_n52) );
  NAND2X0 add_1095_U202 ( .IN1(n9485), .IN2(add_1095_n187), .QN(add_1095_n186)
         );
  OR2X1 add_1095_U187 ( .IN2(n9617), .IN1(add_1095_n31), .Q(add_1095_n175) );
  NAND2X0 add_1095_U188 ( .IN1(n9617), .IN2(add_1095_n31), .QN(add_1095_n173)
         );
  NAND2X0 add_1095_U189 ( .IN1(add_1095_n176), .IN2(add_1095_n177), 
        .QN(add_1095_n31) );
  NAND2X0 add_1095_U190 ( .IN1(n9473), .IN2(add_1095_n178), .QN(add_1095_n177)
         );
  OR2X1 add_1095_U191 ( .IN2(n9621), .IN1(add_1095_n38), .Q(add_1095_n178) );
  NAND2X0 add_1095_U192 ( .IN1(n9621), .IN2(add_1095_n38), .QN(add_1095_n176)
         );
  NAND2X0 add_1095_U193 ( .IN1(add_1095_n179), .IN2(add_1095_n180), 
        .QN(add_1095_n38) );
  NAND2X0 add_1095_U194 ( .IN1(n9477), .IN2(add_1095_n181), .QN(add_1095_n180)
         );
  OR2X1 add_1095_U179 ( .IN2(n9609), .IN1(add_1095_n17), .Q(add_1095_n169) );
  NAND2X0 add_1095_U180 ( .IN1(n9609), .IN2(add_1095_n17), .QN(add_1095_n167)
         );
  NAND2X0 add_1095_U181 ( .IN1(add_1095_n170), .IN2(add_1095_n171), 
        .QN(add_1095_n17) );
  NAND2X0 add_1095_U182 ( .IN1(n9465), .IN2(add_1095_n172), .QN(add_1095_n171)
         );
  OR2X1 add_1095_U183 ( .IN2(n9613), .IN1(add_1095_n24), .Q(add_1095_n172) );
  NAND2X0 add_1095_U184 ( .IN1(n9613), .IN2(add_1095_n24), .QN(add_1095_n170)
         );
  NAND2X0 add_1095_U185 ( .IN1(add_1095_n173), .IN2(add_1095_n174), 
        .QN(add_1095_n24) );
  NAND2X0 add_1095_U186 ( .IN1(n9469), .IN2(add_1095_n175), .QN(add_1095_n174)
         );
  OR2X1 add_1095_U171 ( .IN2(n9601), .IN1(add_1095_n3), .Q(add_1095_n163) );
  NAND2X0 add_1095_U172 ( .IN1(n9601), .IN2(add_1095_n3), .QN(add_1095_n161)
         );
  NAND2X0 add_1095_U173 ( .IN1(add_1095_n164), .IN2(add_1095_n165), 
        .QN(add_1095_n3) );
  NAND2X0 add_1095_U174 ( .IN1(n9457), .IN2(add_1095_n166), .QN(add_1095_n165)
         );
  OR2X1 add_1095_U175 ( .IN2(n9605), .IN1(add_1095_n10), .Q(add_1095_n166) );
  NAND2X0 add_1095_U176 ( .IN1(n9605), .IN2(add_1095_n10), .QN(add_1095_n164)
         );
  NAND2X0 add_1095_U177 ( .IN1(add_1095_n167), .IN2(add_1095_n168), 
        .QN(add_1095_n10) );
  NAND2X0 add_1095_U178 ( .IN1(n9461), .IN2(add_1095_n169), .QN(add_1095_n168)
         );
  AND2X1 add_1095_U163 ( .IN1(add_1095_n154), .IN2(add_1095_n157), 
        .Q(add_1095_n156) );
  NOR2X0 add_1095_U164 ( .QN(add_1095_n155), .IN1(add_1095_n154), 
        .IN2(add_1095_n157) );
  NAND2X0 add_1095_U165 ( .IN1(add_1095_n158), .IN2(add_1095_n159), 
        .QN(add_1095_n157) );
  NAND2X0 add_1095_U166 ( .IN1(n9449), .IN2(add_1095_n160), .QN(add_1095_n159)
         );
  OR2X1 add_1095_U167 ( .IN2(n9449), .IN1(add_1095_n160), .Q(add_1095_n158) );
  INVX0 add_1095_U168 ( .ZN(add_1095_n160), .INP(n9597) );
  NAND2X0 add_1095_U169 ( .IN1(add_1095_n161), .IN2(add_1095_n162), 
        .QN(add_1095_n154) );
  NAND2X0 add_1095_U170 ( .IN1(n9453), .IN2(add_1095_n163), .QN(add_1095_n162)
         );
  NAND2X0 add_1095_U155 ( .IN1(n9445), .IN2(add_1095_n150), .QN(add_1095_n149)
         );
  OR2X1 add_1095_U156 ( .IN2(n9445), .IN1(add_1095_n150), .Q(add_1095_n148) );
  INVX0 add_1095_U157 ( .ZN(add_1095_n150), .INP(n9593) );
  NAND2X0 add_1095_U158 ( .IN1(add_1095_n151), .IN2(add_1095_n152), 
        .QN(add_1095_n144) );
  NAND2X0 add_1095_U159 ( .IN1(n9449), .IN2(add_1095_n153), .QN(add_1095_n152)
         );
  OR2X1 add_1095_U160 ( .IN2(n9597), .IN1(add_1095_n154), .Q(add_1095_n153) );
  NAND2X0 add_1095_U161 ( .IN1(n9597), .IN2(add_1095_n154), .QN(add_1095_n151)
         );
  NOR2X0 add_1095_U162 ( .QN(so_10_), .IN1(add_1095_n155), .IN2(add_1095_n156)
         );
  NAND2X0 add_1095_U147 ( .IN1(add_1095_n141), .IN2(add_1095_n142), 
        .QN(add_1095_n134) );
  NAND2X0 add_1095_U148 ( .IN1(n9445), .IN2(add_1095_n143), .QN(add_1095_n142)
         );
  OR2X1 add_1095_U149 ( .IN2(n9593), .IN1(add_1095_n144), .Q(add_1095_n143) );
  NAND2X0 add_1095_U150 ( .IN1(n9593), .IN2(add_1095_n144), .QN(add_1095_n141)
         );
  NOR2X0 add_1095_U151 ( .QN(so_11_), .IN1(add_1095_n145), .IN2(add_1095_n146)
         );
  AND2X1 add_1095_U152 ( .IN1(add_1095_n144), .IN2(add_1095_n147), 
        .Q(add_1095_n146) );
  NOR2X0 add_1095_U153 ( .QN(add_1095_n145), .IN1(add_1095_n144), 
        .IN2(add_1095_n147) );
  NAND2X0 add_1095_U154 ( .IN1(add_1095_n148), .IN2(add_1095_n149), 
        .QN(add_1095_n147) );
  NAND2X0 add_1095_U139 ( .IN1(n9589), .IN2(add_1095_n134), .QN(add_1095_n131)
         );
  NOR2X0 add_1095_U140 ( .QN(so_12_), .IN1(add_1095_n135), .IN2(add_1095_n136)
         );
  AND2X1 add_1095_U141 ( .IN1(add_1095_n134), .IN2(add_1095_n137), 
        .Q(add_1095_n136) );
  NOR2X0 add_1095_U142 ( .QN(add_1095_n135), .IN1(add_1095_n134), 
        .IN2(add_1095_n137) );
  NAND2X0 add_1095_U143 ( .IN1(add_1095_n138), .IN2(add_1095_n139), 
        .QN(add_1095_n137) );
  NAND2X0 add_1095_U144 ( .IN1(n9441), .IN2(add_1095_n140), .QN(add_1095_n139)
         );
  OR2X1 add_1095_U145 ( .IN2(n9441), .IN1(add_1095_n140), .Q(add_1095_n138) );
  INVX0 add_1095_U146 ( .ZN(add_1095_n140), .INP(n9589) );
  NOR2X0 add_1095_U131 ( .QN(add_1095_n125), .IN1(add_1095_n124), 
        .IN2(add_1095_n127) );
  NAND2X0 add_1095_U132 ( .IN1(add_1095_n128), .IN2(add_1095_n129), 
        .QN(add_1095_n127) );
  NAND2X0 add_1095_U133 ( .IN1(n9437), .IN2(add_1095_n130), .QN(add_1095_n129)
         );
  OR2X1 add_1095_U134 ( .IN2(n9437), .IN1(add_1095_n130), .Q(add_1095_n128) );
  INVX0 add_1095_U135 ( .ZN(add_1095_n130), .INP(n9585) );
  NAND2X0 add_1095_U136 ( .IN1(add_1095_n131), .IN2(add_1095_n132), 
        .QN(add_1095_n124) );
  NAND2X0 add_1095_U137 ( .IN1(n9441), .IN2(add_1095_n133), .QN(add_1095_n132)
         );
  OR2X1 add_1095_U138 ( .IN2(n9589), .IN1(add_1095_n134), .Q(add_1095_n133) );
  OR2X1 add_1095_U123 ( .IN2(n9433), .IN1(add_1095_n120), .Q(add_1095_n118) );
  INVX0 add_1095_U124 ( .ZN(add_1095_n120), .INP(n9581) );
  NAND2X0 add_1095_U125 ( .IN1(add_1095_n121), .IN2(add_1095_n122), 
        .QN(add_1095_n114) );
  NAND2X0 add_1095_U126 ( .IN1(n9437), .IN2(add_1095_n123), .QN(add_1095_n122)
         );
  OR2X1 add_1095_U127 ( .IN2(n9585), .IN1(add_1095_n124), .Q(add_1095_n123) );
  NAND2X0 add_1095_U128 ( .IN1(n9585), .IN2(add_1095_n124), .QN(add_1095_n121)
         );
  NOR2X0 add_1095_U129 ( .QN(so_13_), .IN1(add_1095_n125), .IN2(add_1095_n126)
         );
  AND2X1 add_1095_U130 ( .IN1(add_1095_n124), .IN2(add_1095_n127), 
        .Q(add_1095_n126) );
  NAND2X0 add_1095_U115 ( .IN1(n9433), .IN2(add_1095_n113), .QN(add_1095_n112)
         );
  OR2X1 add_1095_U116 ( .IN2(n9581), .IN1(add_1095_n114), .Q(add_1095_n113) );
  NAND2X0 add_1095_U117 ( .IN1(n9581), .IN2(add_1095_n114), .QN(add_1095_n111)
         );
  NOR2X0 add_1095_U118 ( .QN(so_14_), .IN1(add_1095_n115), .IN2(add_1095_n116)
         );
  AND2X1 add_1095_U119 ( .IN1(add_1095_n114), .IN2(add_1095_n117), 
        .Q(add_1095_n116) );
  NOR2X0 add_1095_U120 ( .QN(add_1095_n115), .IN1(add_1095_n114), 
        .IN2(add_1095_n117) );
  NAND2X0 add_1095_U121 ( .IN1(add_1095_n118), .IN2(add_1095_n119), 
        .QN(add_1095_n117) );
  NAND2X0 add_1095_U122 ( .IN1(n9433), .IN2(add_1095_n120), .QN(add_1095_n119)
         );
  NOR2X0 add_1095_U107 ( .QN(so_15_), .IN1(add_1095_n105), .IN2(add_1095_n106)
         );
  AND2X1 add_1095_U108 ( .IN1(add_1095_n104), .IN2(add_1095_n107), 
        .Q(add_1095_n106) );
  NOR2X0 add_1095_U109 ( .QN(add_1095_n105), .IN1(add_1095_n104), 
        .IN2(add_1095_n107) );
  NAND2X0 add_1095_U110 ( .IN1(add_1095_n108), .IN2(add_1095_n109), 
        .QN(add_1095_n107) );
  NAND2X0 add_1095_U111 ( .IN1(n9429), .IN2(add_1095_n110), .QN(add_1095_n109)
         );
  OR2X1 add_1095_U112 ( .IN2(n9429), .IN1(add_1095_n110), .Q(add_1095_n108) );
  INVX0 add_1095_U113 ( .ZN(add_1095_n110), .INP(n9577) );
  NAND2X0 add_1095_U114 ( .IN1(add_1095_n111), .IN2(add_1095_n112), 
        .QN(add_1095_n104) );
  NAND2X0 add_1095_U99 ( .IN1(add_1095_n98), .IN2(add_1095_n99), 
        .QN(add_1095_n97) );
  NAND2X0 add_1095_U100 ( .IN1(n9425), .IN2(add_1095_n100), .QN(add_1095_n99)
         );
  OR2X1 add_1095_U101 ( .IN2(n9425), .IN1(add_1095_n100), .Q(add_1095_n98) );
  INVX0 add_1095_U102 ( .ZN(add_1095_n100), .INP(n9573) );
  NAND2X0 add_1095_U103 ( .IN1(add_1095_n101), .IN2(add_1095_n102), 
        .QN(add_1095_n94) );
  NAND2X0 add_1095_U104 ( .IN1(n9429), .IN2(add_1095_n103), .QN(add_1095_n102)
         );
  OR2X1 add_1095_U105 ( .IN2(n9577), .IN1(add_1095_n104), .Q(add_1095_n103) );
  NAND2X0 add_1095_U106 ( .IN1(n9577), .IN2(add_1095_n104), .QN(add_1095_n101)
         );
  INVX0 add_1095_U91 ( .ZN(add_1095_n90), .INP(n9569) );
  NAND2X0 add_1095_U92 ( .IN1(add_1095_n91), .IN2(add_1095_n92), 
        .QN(add_1095_n84) );
  NAND2X0 add_1095_U93 ( .IN1(n9425), .IN2(add_1095_n93), .QN(add_1095_n92) );
  OR2X1 add_1095_U94 ( .IN2(n9573), .IN1(add_1095_n94), .Q(add_1095_n93) );
  NAND2X0 add_1095_U95 ( .IN1(n9573), .IN2(add_1095_n94), .QN(add_1095_n91) );
  NOR2X0 add_1095_U96 ( .QN(so_16_), .IN1(add_1095_n95), .IN2(add_1095_n96) );
  AND2X1 add_1095_U97 ( .IN1(add_1095_n94), .IN2(add_1095_n97), 
        .Q(add_1095_n96) );
  NOR2X0 add_1095_U98 ( .QN(add_1095_n95), .IN1(add_1095_n94), 
        .IN2(add_1095_n97) );
  OR2X1 add_1095_U83 ( .IN2(n9569), .IN1(add_1095_n84), .Q(add_1095_n83) );
  NAND2X0 add_1095_U84 ( .IN1(n9569), .IN2(add_1095_n84), .QN(add_1095_n81) );
  NOR2X0 add_1095_U85 ( .QN(so_17_), .IN1(add_1095_n85), .IN2(add_1095_n86) );
  AND2X1 add_1095_U86 ( .IN1(add_1095_n84), .IN2(add_1095_n87), 
        .Q(add_1095_n86) );
  NOR2X0 add_1095_U87 ( .QN(add_1095_n85), .IN1(add_1095_n84), 
        .IN2(add_1095_n87) );
  NAND2X0 add_1095_U88 ( .IN1(add_1095_n88), .IN2(add_1095_n89), 
        .QN(add_1095_n87) );
  NAND2X0 add_1095_U89 ( .IN1(n9421), .IN2(add_1095_n90), .QN(add_1095_n89) );
  OR2X1 add_1095_U90 ( .IN2(n9421), .IN1(add_1095_n90), .Q(add_1095_n88) );
  AND2X1 add_1095_U75 ( .IN1(add_1095_n71), .IN2(add_1095_n77), 
        .Q(add_1095_n76) );
  NOR2X0 add_1095_U76 ( .QN(add_1095_n75), .IN1(add_1095_n71), 
        .IN2(add_1095_n77) );
  NAND2X0 add_1095_U77 ( .IN1(add_1095_n78), .IN2(add_1095_n79), 
        .QN(add_1095_n77) );
  NAND2X0 add_1095_U78 ( .IN1(n9417), .IN2(add_1095_n80), .QN(add_1095_n79) );
  OR2X1 add_1095_U79 ( .IN2(n9417), .IN1(add_1095_n80), .Q(add_1095_n78) );
  INVX0 add_1095_U80 ( .ZN(add_1095_n80), .INP(n9565) );
  NAND2X0 add_1095_U81 ( .IN1(add_1095_n81), .IN2(add_1095_n82), 
        .QN(add_1095_n71) );
  NAND2X0 add_1095_U82 ( .IN1(n9421), .IN2(add_1095_n83), .QN(add_1095_n82) );
  NAND2X0 add_1095_U67 ( .IN1(n9417), .IN2(add_1095_n70), .QN(add_1095_n69) );
  OR2X1 add_1095_U68 ( .IN2(n9565), .IN1(add_1095_n71), .Q(add_1095_n70) );
  NAND2X0 add_1095_U69 ( .IN1(n9565), .IN2(add_1095_n71), .QN(add_1095_n68) );
  NAND2X0 add_1095_U70 ( .IN1(add_1095_n72), .IN2(add_1095_n73), 
        .QN(add_1095_n67) );
  NAND2X0 add_1095_U71 ( .IN1(n18209), .IN2(add_1095_n74), .QN(add_1095_n73)
         );
  OR2X1 add_1095_U72 ( .IN2(n18209), .IN1(add_1095_n74), .Q(add_1095_n72) );
  INVX0 add_1095_U73 ( .ZN(add_1095_n74), .INP(n18245) );
  NOR2X0 add_1095_U74 ( .QN(so_18_), .IN1(add_1095_n75), .IN2(add_1095_n76) );
  NAND2X0 add_1095_U59 ( .IN1(add_1095_n59), .IN2(add_1095_n60), 
        .QN(add_1095_n57) );
  NAND2X0 add_1095_U60 ( .IN1(add_1095_n61), .IN2(add_1095_n62), 
        .QN(add_1095_n59) );
  NAND2X0 add_1095_U61 ( .IN1(n9485), .IN2(add_1095_n63), .QN(add_1095_n62) );
  OR2X1 add_1095_U62 ( .IN2(n9485), .IN1(add_1095_n63), .Q(add_1095_n61) );
  NOR2X0 add_1095_U63 ( .QN(so_19_), .IN1(add_1095_n64), .IN2(add_1095_n65) );
  AND2X1 add_1095_U64 ( .IN1(add_1095_n66), .IN2(add_1095_n67), 
        .Q(add_1095_n65) );
  NOR2X0 add_1095_U65 ( .QN(add_1095_n64), .IN1(add_1095_n67), 
        .IN2(add_1095_n66) );
  NAND2X0 add_1095_U66 ( .IN1(add_1095_n68), .IN2(add_1095_n69), 
        .QN(add_1095_n66) );
  AND2X1 add_1095_U51 ( .IN1(add_1095_n52), .IN2(add_1095_n53), 
        .Q(add_1095_n51) );
  NOR2X0 add_1095_U52 ( .QN(add_1095_n50), .IN1(add_1095_n52), 
        .IN2(add_1095_n53) );
  NAND2X0 add_1095_U53 ( .IN1(add_1095_n54), .IN2(add_1095_n55), 
        .QN(add_1095_n53) );
  NAND2X0 add_1095_U54 ( .IN1(n9481), .IN2(add_1095_n56), .QN(add_1095_n55) );
  OR2X1 add_1095_U55 ( .IN2(n9481), .IN1(add_1095_n56), .Q(add_1095_n54) );
  INVX0 add_1095_U56 ( .ZN(add_1095_n56), .INP(n9629) );
  NAND2X0 add_1095_U57 ( .IN1(add_1095_n57), .IN2(add_1095_n58), .QN(so_1_) );
  OR2X1 add_1095_U58 ( .IN2(add_1095_n60), .IN1(add_1095_n59), 
        .Q(add_1095_n58) );
  NOR2X0 add_1095_U43 ( .QN(so_3_), .IN1(add_1095_n43), .IN2(add_1095_n44) );
  AND2X1 add_1095_U44 ( .IN1(add_1095_n45), .IN2(add_1095_n46), 
        .Q(add_1095_n44) );
  NOR2X0 add_1095_U45 ( .QN(add_1095_n43), .IN1(add_1095_n45), 
        .IN2(add_1095_n46) );
  NAND2X0 add_1095_U46 ( .IN1(add_1095_n47), .IN2(add_1095_n48), 
        .QN(add_1095_n46) );
  NAND2X0 add_1095_U47 ( .IN1(n9477), .IN2(add_1095_n49), .QN(add_1095_n48) );
  OR2X1 add_1095_U48 ( .IN2(n9477), .IN1(add_1095_n49), .Q(add_1095_n47) );
  INVX0 add_1095_U49 ( .ZN(add_1095_n49), .INP(n9625) );
  NOR2X0 add_1095_U50 ( .QN(so_2_), .IN1(add_1095_n50), .IN2(add_1095_n51) );
  INVX0 add_1095_U35 ( .ZN(add_1095_n35), .INP(n9617) );
  NOR2X0 add_1095_U36 ( .QN(so_4_), .IN1(add_1095_n36), .IN2(add_1095_n37) );
  AND2X1 add_1095_U37 ( .IN1(add_1095_n38), .IN2(add_1095_n39), 
        .Q(add_1095_n37) );
  NOR2X0 add_1095_U38 ( .QN(add_1095_n36), .IN1(add_1095_n38), 
        .IN2(add_1095_n39) );
  NAND2X0 add_1095_U39 ( .IN1(add_1095_n40), .IN2(add_1095_n41), 
        .QN(add_1095_n39) );
  NAND2X0 add_1095_U40 ( .IN1(n9473), .IN2(add_1095_n42), .QN(add_1095_n41) );
  OR2X1 add_1095_U41 ( .IN2(n9473), .IN1(add_1095_n42), .Q(add_1095_n40) );
  INVX0 add_1095_U42 ( .ZN(add_1095_n42), .INP(n9621) );
  OR2X1 add_1095_U27 ( .IN2(n9465), .IN1(add_1095_n28), .Q(add_1095_n26) );
  INVX0 add_1095_U28 ( .ZN(add_1095_n28), .INP(n9613) );
  NOR2X0 add_1095_U29 ( .QN(so_5_), .IN1(add_1095_n29), .IN2(add_1095_n30) );
  AND2X1 add_1095_U30 ( .IN1(add_1095_n31), .IN2(add_1095_n32), 
        .Q(add_1095_n30) );
  NOR2X0 add_1095_U31 ( .QN(add_1095_n29), .IN1(add_1095_n31), 
        .IN2(add_1095_n32) );
  NAND2X0 add_1095_U32 ( .IN1(add_1095_n33), .IN2(add_1095_n34), 
        .QN(add_1095_n32) );
  NAND2X0 add_1095_U33 ( .IN1(n9469), .IN2(add_1095_n35), .QN(add_1095_n34) );
  OR2X1 add_1095_U34 ( .IN2(n9469), .IN1(add_1095_n35), .Q(add_1095_n33) );
  NAND2X0 add_1095_U19 ( .IN1(n9461), .IN2(add_1095_n21), .QN(add_1095_n20) );
  OR2X1 add_1095_U20 ( .IN2(n9461), .IN1(add_1095_n21), .Q(add_1095_n19) );
  INVX0 add_1095_U21 ( .ZN(add_1095_n21), .INP(n9609) );
  NOR2X0 add_1095_U22 ( .QN(so_6_), .IN1(add_1095_n22), .IN2(add_1095_n23) );
  AND2X1 add_1095_U23 ( .IN1(add_1095_n24), .IN2(add_1095_n25), 
        .Q(add_1095_n23) );
  NOR2X0 add_1095_U24 ( .QN(add_1095_n22), .IN1(add_1095_n24), 
        .IN2(add_1095_n25) );
  NAND2X0 add_1095_U25 ( .IN1(add_1095_n26), .IN2(add_1095_n27), 
        .QN(add_1095_n25) );
  NAND2X0 add_1095_U26 ( .IN1(n9465), .IN2(add_1095_n28), .QN(add_1095_n27) );
  NAND2X0 add_1095_U11 ( .IN1(add_1095_n12), .IN2(add_1095_n13), 
        .QN(add_1095_n11) );
  NAND2X0 add_1095_U12 ( .IN1(n9457), .IN2(add_1095_n14), .QN(add_1095_n13) );
  OR2X1 add_1095_U13 ( .IN2(n9457), .IN1(add_1095_n14), .Q(add_1095_n12) );
  INVX0 add_1095_U14 ( .ZN(add_1095_n14), .INP(n9605) );
  NOR2X0 add_1095_U15 ( .QN(so_7_), .IN1(add_1095_n15), .IN2(add_1095_n16) );
  AND2X1 add_1095_U16 ( .IN1(add_1095_n17), .IN2(add_1095_n18), 
        .Q(add_1095_n16) );
  NOR2X0 add_1095_U17 ( .QN(add_1095_n15), .IN1(add_1095_n17), 
        .IN2(add_1095_n18) );
  NAND2X0 add_1095_U18 ( .IN1(add_1095_n19), .IN2(add_1095_n20), 
        .QN(add_1095_n18) );
  NOR2X0 add_1095_U3 ( .QN(add_1095_n1), .IN1(add_1095_n3), .IN2(add_1095_n4)
         );
  NAND2X0 add_1095_U4 ( .IN1(add_1095_n5), .IN2(add_1095_n6), .QN(add_1095_n4)
         );
  NAND2X0 add_1095_U5 ( .IN1(n9453), .IN2(add_1095_n7), .QN(add_1095_n6) );
  OR2X1 add_1095_U6 ( .IN2(n9453), .IN1(add_1095_n7), .Q(add_1095_n5) );
  INVX0 add_1095_U7 ( .ZN(add_1095_n7), .INP(n9601) );
  NOR2X0 add_1095_U8 ( .QN(so_8_), .IN1(add_1095_n8), .IN2(add_1095_n9) );
  AND2X1 add_1095_U9 ( .IN1(add_1095_n10), .IN2(add_1095_n11), .Q(add_1095_n9)
         );
  NOR2X0 add_1095_U10 ( .QN(add_1095_n8), .IN1(add_1095_n10), 
        .IN2(add_1095_n11) );
  NOR2X0 add_1095_U1 ( .QN(so_9_), .IN1(add_1095_n1), .IN2(add_1095_n2) );
  AND2X1 add_1095_U2 ( .IN1(add_1095_n3), .IN2(add_1095_n4), .Q(add_1095_n2)
         );
  NOR2X0 P2_sub_621_U39 ( .QN(P2_N131), .IN1(P2_sub_621_n34), 
        .IN2(P2_sub_621_n35) );
  OR2X1 P2_sub_621_U38 ( .IN2(n6595), .IN1(n6596), .Q(P2_sub_621_n33) );
  AND2X1 P2_sub_621_U37 ( .IN1(P2_sub_621_n33), .IN2(n6597), 
        .Q(P2_sub_621_n31) );
  NOR2X0 P2_sub_621_U36 ( .QN(P2_sub_621_n32), .IN1(n6597), 
        .IN2(P2_sub_621_n33) );
  NOR2X0 P2_sub_621_U35 ( .QN(P2_N104), .IN1(P2_sub_621_n31), 
        .IN2(P2_sub_621_n32) );
  OR2X1 P2_sub_621_U34 ( .IN2(n10133), .IN1(P2_sub_621_n30), 
        .Q(P2_sub_621_n27) );
  AND2X1 P2_sub_621_U33 ( .IN1(P2_sub_621_n27), .IN2(n10137), 
        .Q(P2_sub_621_n28) );
  NOR2X0 P2_sub_621_U32 ( .QN(P2_sub_621_n29), .IN1(n10137), 
        .IN2(P2_sub_621_n27) );
  NOR2X0 P2_sub_621_U31 ( .QN(P2_N132), .IN1(P2_sub_621_n28), 
        .IN2(P2_sub_621_n29) );
  OR2X1 P2_sub_621_U30 ( .IN2(n10137), .IN1(P2_sub_621_n27), 
        .Q(P2_sub_621_n26) );
  AND2X1 P2_sub_621_U29 ( .IN1(P2_sub_621_n26), .IN2(n6688), 
        .Q(P2_sub_621_n24) );
  NOR2X0 P2_sub_621_U28 ( .QN(P2_sub_621_n25), .IN1(n6688), 
        .IN2(P2_sub_621_n26) );
  NOR2X0 P2_sub_621_U27 ( .QN(P2_N133), .IN1(P2_sub_621_n24), 
        .IN2(P2_sub_621_n25) );
  AND2X1 P2_sub_621_U26 ( .IN1(P2_sub_621_n21), .IN2(n6598), 
        .Q(P2_sub_621_n22) );
  NOR2X0 P2_sub_621_U25 ( .QN(P2_sub_621_n23), .IN1(n6598), 
        .IN2(P2_sub_621_n21) );
  NOR2X0 P2_sub_621_U24 ( .QN(P2_N105), .IN1(P2_sub_621_n22), 
        .IN2(P2_sub_621_n23) );
  OR2X1 P2_sub_621_U23 ( .IN2(n6598), .IN1(P2_sub_621_n21), .Q(P2_sub_621_n20)
         );
  AND2X1 P2_sub_621_U22 ( .IN1(P2_sub_621_n20), .IN2(n6599), 
        .Q(P2_sub_621_n18) );
  NOR2X0 P2_sub_621_U21 ( .QN(P2_sub_621_n19), .IN1(n6599), 
        .IN2(P2_sub_621_n20) );
  NOR2X0 P2_sub_621_U20 ( .QN(P2_N106), .IN1(P2_sub_621_n18), 
        .IN2(P2_sub_621_n19) );
  INVX0 P2_sub_621_U19 ( .ZN(P2_sub_621_n14), .INP(P2_sub_621_n17) );
  AND2X1 P2_sub_621_U18 ( .IN1(P2_sub_621_n14), .IN2(n6600), 
        .Q(P2_sub_621_n15) );
  NOR2X0 P2_sub_621_U17 ( .QN(P2_sub_621_n16), .IN1(n6600), 
        .IN2(P2_sub_621_n14) );
  NOR2X0 P2_sub_621_U16 ( .QN(P2_N107), .IN1(P2_sub_621_n15), 
        .IN2(P2_sub_621_n16) );
  OR2X1 P2_sub_621_U15 ( .IN2(n6600), .IN1(P2_sub_621_n14), .Q(P2_sub_621_n13)
         );
  AND2X1 P2_sub_621_U14 ( .IN1(P2_sub_621_n13), .IN2(n6601), 
        .Q(P2_sub_621_n11) );
  NOR2X0 P2_sub_621_U13 ( .QN(P2_sub_621_n12), .IN1(n6601), 
        .IN2(P2_sub_621_n13) );
  NOR2X0 P2_sub_621_U12 ( .QN(P2_N108), .IN1(P2_sub_621_n11), 
        .IN2(P2_sub_621_n12) );
  AND2X1 P2_sub_621_U11 ( .IN1(P2_sub_621_n8), .IN2(n6602), .Q(P2_sub_621_n9)
         );
  NOR2X0 P2_sub_621_U10 ( .QN(P2_sub_621_n10), .IN1(n6602), 
        .IN2(P2_sub_621_n8) );
  NOR2X0 P2_sub_621_U9 ( .QN(P2_N109), .IN1(P2_sub_621_n9), 
        .IN2(P2_sub_621_n10) );
  OR2X1 P2_sub_621_U8 ( .IN2(n6602), .IN1(P2_sub_621_n8), .Q(P2_sub_621_n7) );
  AND2X1 P2_sub_621_U7 ( .IN1(P2_sub_621_n7), .IN2(n6603), .Q(P2_sub_621_n5)
         );
  NOR2X0 P2_sub_621_U6 ( .QN(P2_sub_621_n6), .IN1(n6603), .IN2(P2_sub_621_n7)
         );
  NOR2X0 P2_sub_621_U5 ( .QN(P2_N110), .IN1(P2_sub_621_n5), 
        .IN2(P2_sub_621_n6) );
  AND2X1 P2_sub_621_U4 ( .IN1(P2_sub_621_n4), .IN2(n6604), .Q(P2_sub_621_n2)
         );
  NOR2X0 P2_sub_621_U3 ( .QN(P2_sub_621_n3), .IN1(n6604), .IN2(P2_sub_621_n4)
         );
  NOR2X0 P2_sub_621_U2 ( .QN(P2_N111), .IN1(P2_sub_621_n2), 
        .IN2(P2_sub_621_n3) );
  NOR2X0 P2_sub_621_U132 ( .QN(P2_sub_621_n107), .IN1(n6604), .IN2(n6605) );
  NAND2X0 P2_sub_621_U131 ( .IN1(P2_sub_621_n107), .IN2(P2_sub_621_n108), 
        .QN(P2_sub_621_n101) );
  AND2X1 P2_sub_621_U130 ( .IN1(P2_sub_621_n101), .IN2(n6606), 
        .Q(P2_sub_621_n105) );
  NOR2X0 P2_sub_621_U129 ( .QN(P2_sub_621_n106), .IN1(n6606), 
        .IN2(P2_sub_621_n101) );
  NOR2X0 P2_sub_621_U128 ( .QN(P2_N113), .IN1(P2_sub_621_n105), 
        .IN2(P2_sub_621_n106) );
  OR2X1 P2_sub_621_U127 ( .IN2(n6606), .IN1(P2_sub_621_n101), 
        .Q(P2_sub_621_n104) );
  AND2X1 P2_sub_621_U126 ( .IN1(P2_sub_621_n104), .IN2(n6607), 
        .Q(P2_sub_621_n102) );
  NOR2X0 P2_sub_621_U125 ( .QN(P2_sub_621_n103), .IN1(n6607), 
        .IN2(P2_sub_621_n104) );
  NOR2X0 P2_sub_621_U124 ( .QN(P2_N114), .IN1(P2_sub_621_n102), 
        .IN2(P2_sub_621_n103) );
  OR2X1 P2_sub_621_U123 ( .IN2(n6606), .IN1(n6607), .Q(P2_sub_621_n100) );
  NOR2X0 P2_sub_621_U122 ( .QN(P2_sub_621_n93), .IN1(P2_sub_621_n100), 
        .IN2(P2_sub_621_n101) );
  INVX0 P2_sub_621_U121 ( .ZN(P2_sub_621_n97), .INP(P2_sub_621_n93) );
  AND2X1 P2_sub_621_U120 ( .IN1(P2_sub_621_n97), .IN2(n6617), 
        .Q(P2_sub_621_n98) );
  NOR2X0 P2_sub_621_U119 ( .QN(P2_sub_621_n99), .IN1(n6617), 
        .IN2(P2_sub_621_n97) );
  NOR2X0 P2_sub_621_U118 ( .QN(P2_N115), .IN1(P2_sub_621_n98), 
        .IN2(P2_sub_621_n99) );
  OR2X1 P2_sub_621_U117 ( .IN2(n6617), .IN1(P2_sub_621_n97), 
        .Q(P2_sub_621_n96) );
  AND2X1 P2_sub_621_U116 ( .IN1(P2_sub_621_n96), .IN2(n6616), 
        .Q(P2_sub_621_n94) );
  NOR2X0 P2_sub_621_U115 ( .QN(P2_sub_621_n95), .IN1(n6616), 
        .IN2(P2_sub_621_n96) );
  NOR2X0 P2_sub_621_U114 ( .QN(P2_N116), .IN1(P2_sub_621_n94), 
        .IN2(P2_sub_621_n95) );
  NOR2X0 P2_sub_621_U113 ( .QN(P2_sub_621_n92), .IN1(n6616), .IN2(n6617) );
  NAND2X0 P2_sub_621_U112 ( .IN1(P2_sub_621_n92), .IN2(P2_sub_621_n93), 
        .QN(P2_sub_621_n86) );
  AND2X1 P2_sub_621_U111 ( .IN1(P2_sub_621_n86), .IN2(n6615), 
        .Q(P2_sub_621_n90) );
  NOR2X0 P2_sub_621_U110 ( .QN(P2_sub_621_n91), .IN1(n6615), 
        .IN2(P2_sub_621_n86) );
  NOR2X0 P2_sub_621_U109 ( .QN(P2_N117), .IN1(P2_sub_621_n90), 
        .IN2(P2_sub_621_n91) );
  OR2X1 P2_sub_621_U108 ( .IN2(n6615), .IN1(P2_sub_621_n86), 
        .Q(P2_sub_621_n89) );
  AND2X1 P2_sub_621_U107 ( .IN1(P2_sub_621_n89), .IN2(n6614), 
        .Q(P2_sub_621_n87) );
  NOR2X0 P2_sub_621_U106 ( .QN(P2_sub_621_n88), .IN1(n6614), 
        .IN2(P2_sub_621_n89) );
  NOR2X0 P2_sub_621_U105 ( .QN(P2_N118), .IN1(P2_sub_621_n87), 
        .IN2(P2_sub_621_n88) );
  OR2X1 P2_sub_621_U104 ( .IN2(n6615), .IN1(n6614), .Q(P2_sub_621_n85) );
  NOR2X0 P2_sub_621_U103 ( .QN(P2_sub_621_n78), .IN1(P2_sub_621_n85), 
        .IN2(P2_sub_621_n86) );
  INVX0 P2_sub_621_U102 ( .ZN(P2_sub_621_n82), .INP(P2_sub_621_n78) );
  AND2X1 P2_sub_621_U101 ( .IN1(P2_sub_621_n82), .IN2(n6613), 
        .Q(P2_sub_621_n83) );
  NOR2X0 P2_sub_621_U100 ( .QN(P2_sub_621_n84), .IN1(n6613), 
        .IN2(P2_sub_621_n82) );
  NOR2X0 P2_sub_621_U99 ( .QN(P2_N119), .IN1(P2_sub_621_n83), 
        .IN2(P2_sub_621_n84) );
  OR2X1 P2_sub_621_U98 ( .IN2(n6613), .IN1(P2_sub_621_n82), .Q(P2_sub_621_n81)
         );
  AND2X1 P2_sub_621_U97 ( .IN1(P2_sub_621_n81), .IN2(n6612), 
        .Q(P2_sub_621_n79) );
  NOR2X0 P2_sub_621_U96 ( .QN(P2_sub_621_n80), .IN1(n6612), 
        .IN2(P2_sub_621_n81) );
  NOR2X0 P2_sub_621_U95 ( .QN(P2_N120), .IN1(P2_sub_621_n79), 
        .IN2(P2_sub_621_n80) );
  NOR2X0 P2_sub_621_U94 ( .QN(P2_sub_621_n77), .IN1(n6612), .IN2(n6613) );
  NAND2X0 P2_sub_621_U93 ( .IN1(P2_sub_621_n77), .IN2(P2_sub_621_n78), 
        .QN(P2_sub_621_n68) );
  AND2X1 P2_sub_621_U92 ( .IN1(P2_sub_621_n68), .IN2(n6611), 
        .Q(P2_sub_621_n75) );
  NOR2X0 P2_sub_621_U91 ( .QN(P2_sub_621_n76), .IN1(n6611), 
        .IN2(P2_sub_621_n68) );
  NOR2X0 P2_sub_621_U90 ( .QN(P2_N121), .IN1(P2_sub_621_n75), 
        .IN2(P2_sub_621_n76) );
  OR2X1 P2_sub_621_U89 ( .IN2(n6596), .IN1(n18347), .Q(P2_sub_621_n72) );
  NAND2X0 P2_sub_621_U88 ( .IN1(n6596), .IN2(n18347), .QN(P2_sub_621_n73) );
  NAND2X0 P2_sub_621_U87 ( .IN1(P2_sub_621_n72), .IN2(P2_sub_621_n73), 
        .QN(P2_N103) );
  OR2X1 P2_sub_621_U86 ( .IN2(n6611), .IN1(P2_sub_621_n68), .Q(P2_sub_621_n71)
         );
  AND2X1 P2_sub_621_U85 ( .IN1(P2_sub_621_n71), .IN2(n6610), 
        .Q(P2_sub_621_n69) );
  NOR2X0 P2_sub_621_U84 ( .QN(P2_sub_621_n70), .IN1(n6610), 
        .IN2(P2_sub_621_n71) );
  NOR2X0 P2_sub_621_U83 ( .QN(P2_N122), .IN1(P2_sub_621_n69), 
        .IN2(P2_sub_621_n70) );
  OR2X1 P2_sub_621_U82 ( .IN2(n6611), .IN1(n6610), .Q(P2_sub_621_n67) );
  NOR2X0 P2_sub_621_U81 ( .QN(P2_sub_621_n60), .IN1(P2_sub_621_n67), 
        .IN2(P2_sub_621_n68) );
  INVX0 P2_sub_621_U80 ( .ZN(P2_sub_621_n64), .INP(P2_sub_621_n60) );
  AND2X1 P2_sub_621_U79 ( .IN1(P2_sub_621_n64), .IN2(n6609), 
        .Q(P2_sub_621_n65) );
  NOR2X0 P2_sub_621_U78 ( .QN(P2_sub_621_n66), .IN1(n6609), 
        .IN2(P2_sub_621_n64) );
  NOR2X0 P2_sub_621_U77 ( .QN(P2_N123), .IN1(P2_sub_621_n65), 
        .IN2(P2_sub_621_n66) );
  OR2X1 P2_sub_621_U76 ( .IN2(n6609), .IN1(P2_sub_621_n64), .Q(P2_sub_621_n63)
         );
  AND2X1 P2_sub_621_U75 ( .IN1(P2_sub_621_n63), .IN2(n6608), 
        .Q(P2_sub_621_n61) );
  NOR2X0 P2_sub_621_U74 ( .QN(P2_sub_621_n62), .IN1(n6608), 
        .IN2(P2_sub_621_n63) );
  NOR2X0 P2_sub_621_U73 ( .QN(P2_N124), .IN1(P2_sub_621_n61), 
        .IN2(P2_sub_621_n62) );
  NOR2X0 P2_sub_621_U72 ( .QN(P2_sub_621_n59), .IN1(n6608), .IN2(n6609) );
  NAND2X0 P2_sub_621_U71 ( .IN1(P2_sub_621_n59), .IN2(P2_sub_621_n60), 
        .QN(P2_sub_621_n53) );
  AND2X1 P2_sub_621_U70 ( .IN1(P2_sub_621_n53), .IN2(n6719), 
        .Q(P2_sub_621_n57) );
  NOR2X0 P2_sub_621_U69 ( .QN(P2_sub_621_n58), .IN1(n6719), 
        .IN2(P2_sub_621_n53) );
  NOR2X0 P2_sub_621_U68 ( .QN(P2_N125), .IN1(P2_sub_621_n57), 
        .IN2(P2_sub_621_n58) );
  OR2X1 P2_sub_621_U67 ( .IN2(n6719), .IN1(P2_sub_621_n53), .Q(P2_sub_621_n56)
         );
  AND2X1 P2_sub_621_U66 ( .IN1(P2_sub_621_n56), .IN2(n10191), 
        .Q(P2_sub_621_n54) );
  NOR2X0 P2_sub_621_U65 ( .QN(P2_sub_621_n55), .IN1(n10191), 
        .IN2(P2_sub_621_n56) );
  NOR2X0 P2_sub_621_U64 ( .QN(P2_N126), .IN1(P2_sub_621_n54), 
        .IN2(P2_sub_621_n55) );
  OR2X1 P2_sub_621_U63 ( .IN2(n6719), .IN1(n10191), .Q(P2_sub_621_n52) );
  NOR2X0 P2_sub_621_U62 ( .QN(P2_sub_621_n45), .IN1(P2_sub_621_n52), 
        .IN2(P2_sub_621_n53) );
  INVX0 P2_sub_621_U61 ( .ZN(P2_sub_621_n49), .INP(P2_sub_621_n45) );
  AND2X1 P2_sub_621_U60 ( .IN1(P2_sub_621_n49), .IN2(n10377), 
        .Q(P2_sub_621_n50) );
  NOR2X0 P2_sub_621_U59 ( .QN(P2_sub_621_n51), .IN1(n10377), 
        .IN2(P2_sub_621_n49) );
  NOR2X0 P2_sub_621_U58 ( .QN(P2_N127), .IN1(P2_sub_621_n50), 
        .IN2(P2_sub_621_n51) );
  OR2X1 P2_sub_621_U57 ( .IN2(n10377), .IN1(P2_sub_621_n49), 
        .Q(P2_sub_621_n48) );
  AND2X1 P2_sub_621_U56 ( .IN1(P2_sub_621_n48), .IN2(n10183), 
        .Q(P2_sub_621_n46) );
  NOR2X0 P2_sub_621_U55 ( .QN(P2_sub_621_n47), .IN1(n10183), 
        .IN2(P2_sub_621_n48) );
  NOR2X0 P2_sub_621_U54 ( .QN(P2_N128), .IN1(P2_sub_621_n46), 
        .IN2(P2_sub_621_n47) );
  NOR2X0 P2_sub_621_U53 ( .QN(P2_sub_621_n44), .IN1(n10183), .IN2(n10377) );
  NAND2X0 P2_sub_621_U52 ( .IN1(P2_sub_621_n44), .IN2(P2_sub_621_n45), 
        .QN(P2_sub_621_n38) );
  AND2X1 P2_sub_621_U51 ( .IN1(P2_sub_621_n38), .IN2(n10369), 
        .Q(P2_sub_621_n42) );
  NOR2X0 P2_sub_621_U50 ( .QN(P2_sub_621_n43), .IN1(n10369), 
        .IN2(P2_sub_621_n38) );
  NOR2X0 P2_sub_621_U49 ( .QN(P2_N129), .IN1(P2_sub_621_n42), 
        .IN2(P2_sub_621_n43) );
  OR2X1 P2_sub_621_U48 ( .IN2(n10369), .IN1(P2_sub_621_n38), 
        .Q(P2_sub_621_n41) );
  AND2X1 P2_sub_621_U47 ( .IN1(P2_sub_621_n41), .IN2(n10141), 
        .Q(P2_sub_621_n39) );
  NOR2X0 P2_sub_621_U46 ( .QN(P2_sub_621_n40), .IN1(n10141), 
        .IN2(P2_sub_621_n41) );
  NOR2X0 P2_sub_621_U45 ( .QN(P2_N130), .IN1(P2_sub_621_n39), 
        .IN2(P2_sub_621_n40) );
  NOR2X0 P2_sub_621_U44 ( .QN(P2_sub_621_n36), .IN1(n10141), .IN2(n10369) );
  INVX0 P2_sub_621_U43 ( .ZN(P2_sub_621_n37), .INP(P2_sub_621_n38) );
  NAND2X0 P2_sub_621_U42 ( .IN1(P2_sub_621_n36), .IN2(P2_sub_621_n37), 
        .QN(P2_sub_621_n30) );
  AND2X1 P2_sub_621_U41 ( .IN1(P2_sub_621_n30), .IN2(n10133), 
        .Q(P2_sub_621_n34) );
  NOR2X0 P2_sub_621_U40 ( .QN(P2_sub_621_n35), .IN1(n10133), 
        .IN2(P2_sub_621_n30) );
  OR2X1 P2_sub_621_U146 ( .IN2(n6602), .IN1(n6603), .Q(P2_sub_621_n112) );
  NOR2X0 P2_sub_621_U145 ( .QN(P2_sub_621_n113), .IN1(n6601), .IN2(n6600) );
  OR2X1 P2_sub_621_U144 ( .IN2(n6598), .IN1(n6599), .Q(P2_sub_621_n114) );
  NOR2X0 P2_sub_621_U143 ( .QN(P2_sub_621_n115), .IN1(n6597), .IN2(n6596) );
  NAND2X0 P2_sub_621_U141 ( .IN1(P2_sub_621_n115), .IN2(n18347), 
        .QN(P2_sub_621_n21) );
  NOR2X0 P2_sub_621_U140 ( .QN(P2_sub_621_n17), .IN1(P2_sub_621_n114), 
        .IN2(P2_sub_621_n21) );
  NAND2X0 P2_sub_621_U139 ( .IN1(P2_sub_621_n113), .IN2(P2_sub_621_n17), 
        .QN(P2_sub_621_n8) );
  NOR2X0 P2_sub_621_U138 ( .QN(P2_sub_621_n108), .IN1(P2_sub_621_n112), 
        .IN2(P2_sub_621_n8) );
  INVX0 P2_sub_621_U137 ( .ZN(P2_sub_621_n4), .INP(P2_sub_621_n108) );
  OR2X1 P2_sub_621_U136 ( .IN2(n6604), .IN1(P2_sub_621_n4), 
        .Q(P2_sub_621_n111) );
  AND2X1 P2_sub_621_U135 ( .IN1(P2_sub_621_n111), .IN2(n6605), 
        .Q(P2_sub_621_n109) );
  NOR2X0 P2_sub_621_U134 ( .QN(P2_sub_621_n110), .IN1(n6605), 
        .IN2(P2_sub_621_n111) );
  NOR2X0 P2_sub_621_U133 ( .QN(P2_N112), .IN1(P2_sub_621_n109), 
        .IN2(P2_sub_621_n110) );
  OR2X1 r837_U64 ( .IN2(n10112), .IN1(n6771), .Q(r837_n74) );
  NAND2X0 r837_U63 ( .IN1(n10112), .IN2(n6771), .QN(r837_n75) );
  NAND2X0 r837_U62 ( .IN1(r837_n74), .IN2(r837_n75), .QN(r837_n68) );
  NAND2X0 r837_U61 ( .IN1(P2_N345), .IN2(r837_n73), .QN(r837_n69) );
  OR2X1 r837_U60 ( .IN2(P2_N345), .IN1(r837_n73), .Q(r837_n71) );
  NAND2X0 r837_U59 ( .IN1(r837_n71), .IN2(n18907), .QN(r837_n70) );
  NAND2X0 r837_U58 ( .IN1(r837_n69), .IN2(r837_n70), .QN(r837_n67) );
  NAND2X0 r837_U57 ( .IN1(r837_n68), .IN2(r837_n67), .QN(r837_n65) );
  OR2X1 r837_U56 ( .IN2(r837_n68), .IN1(r837_n67), .Q(r837_n66) );
  NAND2X0 r837_U55 ( .IN1(r837_n65), .IN2(r837_n66), .QN(n116) );
  NAND2X0 r837_U54 ( .IN1(P2_N362), .IN2(n18939), .QN(r837_n61) );
  NAND2X0 r837_U53 ( .IN1(n6664), .IN2(n6733), .QN(r837_n62) );
  NAND2X0 r837_U52 ( .IN1(r837_n61), .IN2(r837_n62), .QN(r837_n59) );
  NAND2X0 r837_U51 ( .IN1(r837_n59), .IN2(r837_n60), .QN(r837_n57) );
  OR2X1 r837_U50 ( .IN2(r837_n60), .IN1(r837_n59), .Q(r837_n58) );
  NAND2X0 r837_U49 ( .IN1(r837_n57), .IN2(r837_n58), .QN(n134) );
  NAND2X0 r837_U48 ( .IN1(P2_N361), .IN2(n18937), .QN(r837_n54) );
  OR2X1 r837_U47 ( .IN2(P2_N361), .IN1(n18937), .Q(r837_n55) );
  NAND2X0 r837_U46 ( .IN1(r837_n54), .IN2(r837_n55), .QN(r837_n52) );
  NAND2X0 r837_U45 ( .IN1(r837_n52), .IN2(r837_n53), .QN(r837_n50) );
  OR2X1 r837_U44 ( .IN2(r837_n53), .IN1(r837_n52), .Q(r837_n51) );
  NAND2X0 r837_U43 ( .IN1(r837_n50), .IN2(r837_n51), .QN(n133) );
  NAND2X0 r837_U42 ( .IN1(P2_N360), .IN2(n18935), .QN(r837_n47) );
  OR2X1 r837_U41 ( .IN2(P2_N360), .IN1(n18935), .Q(r837_n48) );
  NAND2X0 r837_U40 ( .IN1(r837_n47), .IN2(r837_n48), .QN(r837_n45) );
  NAND2X0 r837_U39 ( .IN1(r837_n45), .IN2(r837_n46), .QN(r837_n43) );
  OR2X1 r837_U38 ( .IN2(r837_n46), .IN1(r837_n45), .Q(r837_n44) );
  NAND2X0 r837_U37 ( .IN1(r837_n43), .IN2(r837_n44), .QN(n132) );
  NAND2X0 r837_U36 ( .IN1(P2_N359), .IN2(n18933), .QN(r837_n40) );
  OR2X1 r837_U35 ( .IN2(P2_N359), .IN1(n18933), .Q(r837_n41) );
  NAND2X0 r837_U34 ( .IN1(r837_n40), .IN2(r837_n41), .QN(r837_n38) );
  NAND2X0 r837_U33 ( .IN1(r837_n38), .IN2(r837_n39), .QN(r837_n36) );
  OR2X1 r837_U32 ( .IN2(r837_n39), .IN1(r837_n38), .Q(r837_n37) );
  NAND2X0 r837_U31 ( .IN1(r837_n36), .IN2(r837_n37), .QN(n131) );
  NAND2X0 r837_U30 ( .IN1(P2_N358), .IN2(n18931), .QN(r837_n33) );
  OR2X1 r837_U29 ( .IN2(P2_N358), .IN1(n18931), .Q(r837_n34) );
  NAND2X0 r837_U28 ( .IN1(r837_n33), .IN2(r837_n34), .QN(r837_n31) );
  NAND2X0 r837_U27 ( .IN1(r837_n31), .IN2(r837_n32), .QN(r837_n29) );
  OR2X1 r837_U26 ( .IN2(r837_n32), .IN1(r837_n31), .Q(r837_n30) );
  NAND2X0 r837_U25 ( .IN1(r837_n29), .IN2(r837_n30), .QN(n130) );
  NAND2X0 r837_U24 ( .IN1(P2_N357), .IN2(n18929), .QN(r837_n26) );
  OR2X1 r837_U23 ( .IN2(P2_N357), .IN1(n18929), .Q(r837_n27) );
  NAND2X0 r837_U22 ( .IN1(r837_n26), .IN2(r837_n27), .QN(r837_n24) );
  NAND2X0 r837_U21 ( .IN1(r837_n24), .IN2(r837_n25), .QN(r837_n22) );
  OR2X1 r837_U20 ( .IN2(r837_n25), .IN1(r837_n24), .Q(r837_n23) );
  NAND2X0 r837_U19 ( .IN1(r837_n22), .IN2(r837_n23), .QN(n129) );
  NAND2X0 r837_U18 ( .IN1(P2_N356), .IN2(n18927), .QN(r837_n19) );
  OR2X1 r837_U17 ( .IN2(P2_N356), .IN1(n18927), .Q(r837_n20) );
  NAND2X0 r837_U16 ( .IN1(r837_n19), .IN2(r837_n20), .QN(r837_n17) );
  NAND2X0 r837_U15 ( .IN1(r837_n17), .IN2(r837_n18), .QN(r837_n15) );
  OR2X1 r837_U14 ( .IN2(r837_n18), .IN1(r837_n17), .Q(r837_n16) );
  NAND2X0 r837_U13 ( .IN1(r837_n15), .IN2(r837_n16), .QN(n128) );
  NAND2X0 r837_U12 ( .IN1(P2_N355), .IN2(r837_n14), .QN(r837_n12) );
  OR2X1 r837_U11 ( .IN2(P2_N355), .IN1(r837_n14), .Q(r837_n13) );
  NAND2X0 r837_U10 ( .IN1(r837_n12), .IN2(r837_n13), .QN(r837_n10) );
  NAND2X0 r837_U9 ( .IN1(r837_n10), .IN2(r837_n11), .QN(r837_n8) );
  OR2X1 r837_U8 ( .IN2(r837_n11), .IN1(r837_n10), .Q(r837_n9) );
  NAND2X0 r837_U7 ( .IN1(r837_n8), .IN2(r837_n9), .QN(n127) );
  NAND2X0 r837_U6 ( .IN1(P2_N354), .IN2(n18925), .QN(r837_n5) );
  OR2X1 r837_U5 ( .IN2(P2_N354), .IN1(n18925), .Q(r837_n6) );
  NAND2X0 r837_U4 ( .IN1(r837_n5), .IN2(r837_n6), .QN(r837_n3) );
  NAND2X0 r837_U3 ( .IN1(r837_n3), .IN2(r837_n4), .QN(r837_n1) );
  OR2X1 r837_U2 ( .IN2(r837_n4), .IN1(r837_n3), .Q(r837_n2) );
  NAND2X0 r837_U1 ( .IN1(r837_n1), .IN2(r837_n2), .QN(n126) );
  NAND2X0 r837_U157 ( .IN1(r837_n160), .IN2(r837_n161), .QN(r837_n154) );
  NAND2X0 r837_U156 ( .IN1(r837_n159), .IN2(r837_n154), .QN(r837_n157) );
  OR2X1 r837_U155 ( .IN2(r837_n154), .IN1(r837_n159), .Q(r837_n158) );
  NAND2X0 r837_U154 ( .IN1(r837_n157), .IN2(r837_n158), .QN(n125) );
  NAND2X0 r837_U152 ( .IN1(P2_N352), .IN2(n18921), .QN(r837_n155) );
  OR2X1 r837_U151 ( .IN2(P2_N352), .IN1(n18921), .Q(r837_n156) );
  NAND2X0 r837_U150 ( .IN1(r837_n155), .IN2(r837_n156), .QN(r837_n149) );
  NAND2X0 r837_U149 ( .IN1(P2_N353), .IN2(r837_n154), .QN(r837_n150) );
  OR2X1 r837_U148 ( .IN2(P2_N353), .IN1(r837_n154), .Q(r837_n152) );
  NAND2X0 r837_U147 ( .IN1(r837_n152), .IN2(n18923), .QN(r837_n151) );
  NAND2X0 r837_U146 ( .IN1(r837_n150), .IN2(r837_n151), .QN(r837_n144) );
  NAND2X0 r837_U145 ( .IN1(r837_n149), .IN2(r837_n144), .QN(r837_n147) );
  OR2X1 r837_U144 ( .IN2(r837_n144), .IN1(r837_n149), .Q(r837_n148) );
  NAND2X0 r837_U143 ( .IN1(r837_n147), .IN2(r837_n148), .QN(n124) );
  NAND2X0 r837_U141 ( .IN1(P2_N351), .IN2(n18919), .QN(r837_n145) );
  OR2X1 r837_U140 ( .IN2(P2_N351), .IN1(n18919), .Q(r837_n146) );
  NAND2X0 r837_U139 ( .IN1(r837_n145), .IN2(r837_n146), .QN(r837_n139) );
  NAND2X0 r837_U138 ( .IN1(P2_N352), .IN2(r837_n144), .QN(r837_n140) );
  OR2X1 r837_U137 ( .IN2(P2_N352), .IN1(r837_n144), .Q(r837_n142) );
  NAND2X0 r837_U136 ( .IN1(r837_n142), .IN2(n18921), .QN(r837_n141) );
  NAND2X0 r837_U135 ( .IN1(r837_n140), .IN2(r837_n141), .QN(r837_n134) );
  NAND2X0 r837_U134 ( .IN1(r837_n139), .IN2(r837_n134), .QN(r837_n137) );
  OR2X1 r837_U133 ( .IN2(r837_n134), .IN1(r837_n139), .Q(r837_n138) );
  NAND2X0 r837_U132 ( .IN1(r837_n137), .IN2(r837_n138), .QN(n123) );
  NAND2X0 r837_U130 ( .IN1(P2_N350), .IN2(n18917), .QN(r837_n135) );
  OR2X1 r837_U129 ( .IN2(P2_N350), .IN1(n18917), .Q(r837_n136) );
  NAND2X0 r837_U128 ( .IN1(r837_n135), .IN2(r837_n136), .QN(r837_n129) );
  NAND2X0 r837_U127 ( .IN1(P2_N351), .IN2(r837_n134), .QN(r837_n130) );
  OR2X1 r837_U126 ( .IN2(P2_N351), .IN1(r837_n134), .Q(r837_n132) );
  NAND2X0 r837_U125 ( .IN1(r837_n132), .IN2(n18919), .QN(r837_n131) );
  NAND2X0 r837_U124 ( .IN1(r837_n130), .IN2(r837_n131), .QN(r837_n124) );
  NAND2X0 r837_U123 ( .IN1(r837_n129), .IN2(r837_n124), .QN(r837_n127) );
  OR2X1 r837_U122 ( .IN2(r837_n124), .IN1(r837_n129), .Q(r837_n128) );
  NAND2X0 r837_U121 ( .IN1(r837_n127), .IN2(r837_n128), .QN(n122) );
  NAND2X0 r837_U119 ( .IN1(P2_N349), .IN2(n18915), .QN(r837_n125) );
  OR2X1 r837_U118 ( .IN2(P2_N349), .IN1(n18915), .Q(r837_n126) );
  NAND2X0 r837_U117 ( .IN1(r837_n125), .IN2(r837_n126), .QN(r837_n119) );
  NAND2X0 r837_U116 ( .IN1(P2_N350), .IN2(r837_n124), .QN(r837_n120) );
  OR2X1 r837_U115 ( .IN2(P2_N350), .IN1(r837_n124), .Q(r837_n122) );
  NAND2X0 r837_U114 ( .IN1(r837_n122), .IN2(n18917), .QN(r837_n121) );
  NAND2X0 r837_U113 ( .IN1(r837_n120), .IN2(r837_n121), .QN(r837_n114) );
  NAND2X0 r837_U112 ( .IN1(r837_n119), .IN2(r837_n114), .QN(r837_n117) );
  OR2X1 r837_U111 ( .IN2(r837_n114), .IN1(r837_n119), .Q(r837_n118) );
  NAND2X0 r837_U110 ( .IN1(r837_n117), .IN2(r837_n118), .QN(n121) );
  NAND2X0 r837_U108 ( .IN1(P2_N348), .IN2(n18913), .QN(r837_n115) );
  OR2X1 r837_U107 ( .IN2(P2_N348), .IN1(n18913), .Q(r837_n116) );
  NAND2X0 r837_U106 ( .IN1(r837_n115), .IN2(r837_n116), .QN(r837_n109) );
  NAND2X0 r837_U105 ( .IN1(P2_N349), .IN2(r837_n114), .QN(r837_n110) );
  OR2X1 r837_U104 ( .IN2(P2_N349), .IN1(r837_n114), .Q(r837_n112) );
  NAND2X0 r837_U103 ( .IN1(r837_n112), .IN2(n18915), .QN(r837_n111) );
  NAND2X0 r837_U102 ( .IN1(r837_n110), .IN2(r837_n111), .QN(r837_n104) );
  NAND2X0 r837_U101 ( .IN1(r837_n109), .IN2(r837_n104), .QN(r837_n107) );
  OR2X1 r837_U100 ( .IN2(r837_n104), .IN1(r837_n109), .Q(r837_n108) );
  NAND2X0 r837_U99 ( .IN1(r837_n107), .IN2(r837_n108), .QN(n120) );
  NAND2X0 r837_U97 ( .IN1(P2_N347), .IN2(n18911), .QN(r837_n105) );
  OR2X1 r837_U96 ( .IN2(P2_N347), .IN1(n18911), .Q(r837_n106) );
  NAND2X0 r837_U95 ( .IN1(r837_n105), .IN2(r837_n106), .QN(r837_n99) );
  NAND2X0 r837_U94 ( .IN1(P2_N348), .IN2(r837_n104), .QN(r837_n100) );
  OR2X1 r837_U93 ( .IN2(P2_N348), .IN1(r837_n104), .Q(r837_n102) );
  NAND2X0 r837_U92 ( .IN1(r837_n102), .IN2(n18913), .QN(r837_n101) );
  NAND2X0 r837_U91 ( .IN1(r837_n100), .IN2(r837_n101), .QN(r837_n94) );
  NAND2X0 r837_U90 ( .IN1(r837_n99), .IN2(r837_n94), .QN(r837_n97) );
  OR2X1 r837_U89 ( .IN2(r837_n94), .IN1(r837_n99), .Q(r837_n98) );
  NAND2X0 r837_U88 ( .IN1(r837_n97), .IN2(r837_n98), .QN(n119) );
  NAND2X0 r837_U86 ( .IN1(P2_N346), .IN2(n18909), .QN(r837_n95) );
  OR2X1 r837_U85 ( .IN2(P2_N346), .IN1(n18909), .Q(r837_n96) );
  NAND2X0 r837_U84 ( .IN1(r837_n95), .IN2(r837_n96), .QN(r837_n89) );
  NAND2X0 r837_U83 ( .IN1(P2_N347), .IN2(r837_n94), .QN(r837_n90) );
  OR2X1 r837_U82 ( .IN2(P2_N347), .IN1(r837_n94), .Q(r837_n92) );
  NAND2X0 r837_U81 ( .IN1(r837_n92), .IN2(n18911), .QN(r837_n91) );
  NAND2X0 r837_U80 ( .IN1(r837_n90), .IN2(r837_n91), .QN(r837_n84) );
  NAND2X0 r837_U79 ( .IN1(r837_n89), .IN2(r837_n84), .QN(r837_n87) );
  OR2X1 r837_U78 ( .IN2(r837_n84), .IN1(r837_n89), .Q(r837_n88) );
  NAND2X0 r837_U77 ( .IN1(r837_n87), .IN2(r837_n88), .QN(n118) );
  NAND2X0 r837_U75 ( .IN1(P2_N345), .IN2(n18907), .QN(r837_n85) );
  OR2X1 r837_U74 ( .IN2(P2_N345), .IN1(n18907), .Q(r837_n86) );
  NAND2X0 r837_U73 ( .IN1(r837_n85), .IN2(r837_n86), .QN(r837_n79) );
  NAND2X0 r837_U72 ( .IN1(P2_N346), .IN2(r837_n84), .QN(r837_n80) );
  OR2X1 r837_U71 ( .IN2(P2_N346), .IN1(r837_n84), .Q(r837_n82) );
  NAND2X0 r837_U70 ( .IN1(r837_n82), .IN2(n18909), .QN(r837_n81) );
  NAND2X0 r837_U69 ( .IN1(r837_n80), .IN2(r837_n81), .QN(r837_n73) );
  NAND2X0 r837_U68 ( .IN1(r837_n79), .IN2(r837_n73), .QN(r837_n77) );
  OR2X1 r837_U67 ( .IN2(r837_n73), .IN1(r837_n79), .Q(r837_n78) );
  NAND2X0 r837_U66 ( .IN1(r837_n77), .IN2(r837_n78), .QN(n117) );
  INVX0 r837_U211 ( .ZN(r837_n191), .INP(n9838) );
  NOR2X0 r837_U210 ( .QN(r837_n187), .IN1(r837_n191), .IN2(P2_N363) );
  INVX0 r837_U209 ( .ZN(r837_n60), .INP(r837_n187) );
  NAND2X0 r837_U208 ( .IN1(P2_N363), .IN2(r837_n191), .QN(r837_n190) );
  NAND2X0 r837_U207 ( .IN1(r837_n60), .IN2(r837_n190), .QN(n135) );
  NAND2X0 r837_U205 ( .IN1(P2_N353), .IN2(n18923), .QN(r837_n188) );
  OR2X1 r837_U204 ( .IN2(P2_N353), .IN1(n18923), .Q(r837_n189) );
  NAND2X0 r837_U203 ( .IN1(r837_n188), .IN2(r837_n189), .QN(r837_n159) );
  NAND2X0 r837_U202 ( .IN1(P2_N362), .IN2(r837_n60), .QN(r837_n184) );
  NAND2X0 r837_U200 ( .IN1(r837_n187), .IN2(n6733), .QN(r837_n186) );
  NAND2X0 r837_U198 ( .IN1(r837_n186), .IN2(n18939), .QN(r837_n185) );
  NAND2X0 r837_U197 ( .IN1(r837_n184), .IN2(r837_n185), .QN(r837_n53) );
  NAND2X0 r837_U196 ( .IN1(P2_N361), .IN2(r837_n53), .QN(r837_n181) );
  OR2X1 r837_U195 ( .IN2(P2_N361), .IN1(r837_n53), .Q(r837_n183) );
  NAND2X0 r837_U193 ( .IN1(r837_n183), .IN2(n18937), .QN(r837_n182) );
  NAND2X0 r837_U192 ( .IN1(r837_n181), .IN2(r837_n182), .QN(r837_n46) );
  NAND2X0 r837_U191 ( .IN1(P2_N360), .IN2(r837_n46), .QN(r837_n178) );
  OR2X1 r837_U190 ( .IN2(P2_N360), .IN1(r837_n46), .Q(r837_n180) );
  NAND2X0 r837_U188 ( .IN1(r837_n180), .IN2(n18935), .QN(r837_n179) );
  NAND2X0 r837_U187 ( .IN1(r837_n178), .IN2(r837_n179), .QN(r837_n39) );
  NAND2X0 r837_U186 ( .IN1(P2_N359), .IN2(r837_n39), .QN(r837_n175) );
  OR2X1 r837_U185 ( .IN2(P2_N359), .IN1(r837_n39), .Q(r837_n177) );
  NAND2X0 r837_U183 ( .IN1(r837_n177), .IN2(n18933), .QN(r837_n176) );
  NAND2X0 r837_U182 ( .IN1(r837_n175), .IN2(r837_n176), .QN(r837_n32) );
  NAND2X0 r837_U181 ( .IN1(P2_N358), .IN2(r837_n32), .QN(r837_n172) );
  OR2X1 r837_U180 ( .IN2(P2_N358), .IN1(r837_n32), .Q(r837_n174) );
  NAND2X0 r837_U178 ( .IN1(r837_n174), .IN2(n18931), .QN(r837_n173) );
  NAND2X0 r837_U177 ( .IN1(r837_n172), .IN2(r837_n173), .QN(r837_n25) );
  NAND2X0 r837_U176 ( .IN1(P2_N357), .IN2(r837_n25), .QN(r837_n169) );
  OR2X1 r837_U175 ( .IN2(P2_N357), .IN1(r837_n25), .Q(r837_n171) );
  NAND2X0 r837_U173 ( .IN1(r837_n171), .IN2(n18929), .QN(r837_n170) );
  NAND2X0 r837_U172 ( .IN1(r837_n169), .IN2(r837_n170), .QN(r837_n18) );
  NAND2X0 r837_U171 ( .IN1(P2_N356), .IN2(r837_n18), .QN(r837_n166) );
  OR2X1 r837_U170 ( .IN2(P2_N356), .IN1(r837_n18), .Q(r837_n168) );
  NAND2X0 r837_U168 ( .IN1(r837_n168), .IN2(n18927), .QN(r837_n167) );
  NAND2X0 r837_U167 ( .IN1(r837_n166), .IN2(r837_n167), .QN(r837_n11) );
  NAND2X0 r837_U166 ( .IN1(P2_N355), .IN2(r837_n11), .QN(r837_n163) );
  OR2X1 r837_U165 ( .IN2(P2_N355), .IN1(r837_n11), .Q(r837_n165) );
  INVX0 r837_U164 ( .ZN(r837_n14), .INP(n10250) );
  NAND2X0 r837_U163 ( .IN1(r837_n165), .IN2(r837_n14), .QN(r837_n164) );
  NAND2X0 r837_U162 ( .IN1(r837_n163), .IN2(r837_n164), .QN(r837_n4) );
  NAND2X0 r837_U161 ( .IN1(P2_N354), .IN2(r837_n4), .QN(r837_n160) );
  OR2X1 r837_U160 ( .IN2(P2_N354), .IN1(r837_n4), .Q(r837_n162) );
  NAND2X0 r837_U158 ( .IN1(r837_n162), .IN2(n18925), .QN(r837_n161) );
  OR2X1 r838_U89 ( .IN2(r838_n94), .IN1(r838_n99), .Q(r838_n98) );
  NAND2X0 r838_U88 ( .IN1(r838_n97), .IN2(r838_n98), .QN(n98) );
  NAND2X0 r838_U86 ( .IN1(P2_N346), .IN2(n18965), .QN(r838_n95) );
  OR2X1 r838_U85 ( .IN2(P2_N346), .IN1(n18965), .Q(r838_n96) );
  NAND2X0 r838_U84 ( .IN1(r838_n95), .IN2(r838_n96), .QN(r838_n89) );
  NAND2X0 r838_U83 ( .IN1(P2_N347), .IN2(r838_n94), .QN(r838_n90) );
  OR2X1 r838_U82 ( .IN2(P2_N347), .IN1(r838_n94), .Q(r838_n92) );
  NAND2X0 r838_U81 ( .IN1(r838_n92), .IN2(n18967), .QN(r838_n91) );
  NAND2X0 r838_U80 ( .IN1(r838_n90), .IN2(r838_n91), .QN(r838_n84) );
  NAND2X0 r838_U79 ( .IN1(r838_n89), .IN2(r838_n84), .QN(r838_n87) );
  OR2X1 r838_U78 ( .IN2(r838_n84), .IN1(r838_n89), .Q(r838_n88) );
  NAND2X0 r838_U77 ( .IN1(r838_n87), .IN2(r838_n88), .QN(n97) );
  NAND2X0 r838_U75 ( .IN1(P2_N345), .IN2(n18963), .QN(r838_n85) );
  OR2X1 r838_U74 ( .IN2(P2_N345), .IN1(n18963), .Q(r838_n86) );
  NAND2X0 r838_U73 ( .IN1(r838_n85), .IN2(r838_n86), .QN(r838_n79) );
  NAND2X0 r838_U72 ( .IN1(P2_N346), .IN2(r838_n84), .QN(r838_n80) );
  OR2X1 r838_U71 ( .IN2(P2_N346), .IN1(r838_n84), .Q(r838_n82) );
  NAND2X0 r838_U70 ( .IN1(r838_n82), .IN2(n18965), .QN(r838_n81) );
  NAND2X0 r838_U69 ( .IN1(r838_n80), .IN2(r838_n81), .QN(r838_n73) );
  NAND2X0 r838_U68 ( .IN1(r838_n79), .IN2(r838_n73), .QN(r838_n77) );
  OR2X1 r838_U67 ( .IN2(r838_n73), .IN1(r838_n79), .Q(r838_n78) );
  NAND2X0 r838_U66 ( .IN1(r838_n77), .IN2(r838_n78), .QN(n96) );
  OR2X1 r838_U64 ( .IN2(n10117), .IN1(n6771), .Q(r838_n74) );
  NAND2X0 r838_U63 ( .IN1(n10117), .IN2(n6771), .QN(r838_n75) );
  NAND2X0 r838_U62 ( .IN1(r838_n74), .IN2(r838_n75), .QN(r838_n68) );
  NAND2X0 r838_U61 ( .IN1(P2_N345), .IN2(r838_n73), .QN(r838_n69) );
  OR2X1 r838_U60 ( .IN2(P2_N345), .IN1(r838_n73), .Q(r838_n71) );
  NAND2X0 r838_U59 ( .IN1(r838_n71), .IN2(n18963), .QN(r838_n70) );
  NAND2X0 r838_U58 ( .IN1(r838_n69), .IN2(r838_n70), .QN(r838_n67) );
  NAND2X0 r838_U57 ( .IN1(r838_n68), .IN2(r838_n67), .QN(r838_n65) );
  OR2X1 r838_U56 ( .IN2(r838_n68), .IN1(r838_n67), .Q(r838_n66) );
  NAND2X0 r838_U55 ( .IN1(r838_n65), .IN2(r838_n66), .QN(n95) );
  NAND2X0 r838_U54 ( .IN1(P2_N362), .IN2(n18997), .QN(r838_n61) );
  NAND2X0 r838_U53 ( .IN1(n6720), .IN2(n6733), .QN(r838_n62) );
  NAND2X0 r838_U52 ( .IN1(r838_n61), .IN2(r838_n62), .QN(r838_n59) );
  NAND2X0 r838_U51 ( .IN1(r838_n59), .IN2(r838_n60), .QN(r838_n57) );
  OR2X1 r838_U50 ( .IN2(r838_n60), .IN1(r838_n59), .Q(r838_n58) );
  NAND2X0 r838_U49 ( .IN1(r838_n57), .IN2(r838_n58), .QN(n113) );
  NAND2X0 r838_U48 ( .IN1(P2_N361), .IN2(n18995), .QN(r838_n54) );
  OR2X1 r838_U47 ( .IN2(P2_N361), .IN1(n18995), .Q(r838_n55) );
  NAND2X0 r838_U46 ( .IN1(r838_n54), .IN2(r838_n55), .QN(r838_n52) );
  NAND2X0 r838_U45 ( .IN1(r838_n52), .IN2(r838_n53), .QN(r838_n50) );
  OR2X1 r838_U44 ( .IN2(r838_n53), .IN1(r838_n52), .Q(r838_n51) );
  NAND2X0 r838_U43 ( .IN1(r838_n50), .IN2(r838_n51), .QN(n112) );
  NAND2X0 r838_U42 ( .IN1(P2_N360), .IN2(n18993), .QN(r838_n47) );
  OR2X1 r838_U41 ( .IN2(P2_N360), .IN1(n18993), .Q(r838_n48) );
  NAND2X0 r838_U40 ( .IN1(r838_n47), .IN2(r838_n48), .QN(r838_n45) );
  NAND2X0 r838_U39 ( .IN1(r838_n45), .IN2(r838_n46), .QN(r838_n43) );
  OR2X1 r838_U38 ( .IN2(r838_n46), .IN1(r838_n45), .Q(r838_n44) );
  NAND2X0 r838_U37 ( .IN1(r838_n43), .IN2(r838_n44), .QN(n111) );
  NAND2X0 r838_U36 ( .IN1(P2_N359), .IN2(n18991), .QN(r838_n40) );
  OR2X1 r838_U35 ( .IN2(P2_N359), .IN1(n18991), .Q(r838_n41) );
  NAND2X0 r838_U34 ( .IN1(r838_n40), .IN2(r838_n41), .QN(r838_n38) );
  NAND2X0 r838_U33 ( .IN1(r838_n38), .IN2(r838_n39), .QN(r838_n36) );
  OR2X1 r838_U32 ( .IN2(r838_n39), .IN1(r838_n38), .Q(r838_n37) );
  NAND2X0 r838_U31 ( .IN1(r838_n36), .IN2(r838_n37), .QN(n110) );
  NAND2X0 r838_U30 ( .IN1(P2_N358), .IN2(n18989), .QN(r838_n33) );
  OR2X1 r838_U29 ( .IN2(P2_N358), .IN1(n18989), .Q(r838_n34) );
  NAND2X0 r838_U28 ( .IN1(r838_n33), .IN2(r838_n34), .QN(r838_n31) );
  NAND2X0 r838_U27 ( .IN1(r838_n31), .IN2(r838_n32), .QN(r838_n29) );
  OR2X1 r838_U26 ( .IN2(r838_n32), .IN1(r838_n31), .Q(r838_n30) );
  NAND2X0 r838_U25 ( .IN1(r838_n29), .IN2(r838_n30), .QN(n109) );
  NAND2X0 r838_U24 ( .IN1(P2_N357), .IN2(n18987), .QN(r838_n26) );
  OR2X1 r838_U23 ( .IN2(P2_N357), .IN1(n18987), .Q(r838_n27) );
  NAND2X0 r838_U22 ( .IN1(r838_n26), .IN2(r838_n27), .QN(r838_n24) );
  NAND2X0 r838_U21 ( .IN1(r838_n24), .IN2(r838_n25), .QN(r838_n22) );
  OR2X1 r838_U20 ( .IN2(r838_n25), .IN1(r838_n24), .Q(r838_n23) );
  NAND2X0 r838_U19 ( .IN1(r838_n22), .IN2(r838_n23), .QN(n108) );
  NAND2X0 r838_U18 ( .IN1(P2_N356), .IN2(n18985), .QN(r838_n19) );
  OR2X1 r838_U17 ( .IN2(P2_N356), .IN1(n18985), .Q(r838_n20) );
  NAND2X0 r838_U16 ( .IN1(r838_n19), .IN2(r838_n20), .QN(r838_n17) );
  NAND2X0 r838_U15 ( .IN1(r838_n17), .IN2(r838_n18), .QN(r838_n15) );
  OR2X1 r838_U14 ( .IN2(r838_n18), .IN1(r838_n17), .Q(r838_n16) );
  NAND2X0 r838_U13 ( .IN1(r838_n15), .IN2(r838_n16), .QN(n107) );
  NAND2X0 r838_U12 ( .IN1(P2_N355), .IN2(n18983), .QN(r838_n12) );
  OR2X1 r838_U11 ( .IN2(P2_N355), .IN1(n18983), .Q(r838_n13) );
  NAND2X0 r838_U10 ( .IN1(r838_n12), .IN2(r838_n13), .QN(r838_n10) );
  NAND2X0 r838_U9 ( .IN1(r838_n10), .IN2(r838_n11), .QN(r838_n8) );
  OR2X1 r838_U8 ( .IN2(r838_n11), .IN1(r838_n10), .Q(r838_n9) );
  NAND2X0 r838_U7 ( .IN1(r838_n8), .IN2(r838_n9), .QN(n106) );
  NAND2X0 r838_U6 ( .IN1(P2_N354), .IN2(n18981), .QN(r838_n5) );
  OR2X1 r838_U5 ( .IN2(P2_N354), .IN1(n18981), .Q(r838_n6) );
  NAND2X0 r838_U4 ( .IN1(r838_n5), .IN2(r838_n6), .QN(r838_n3) );
  NAND2X0 r838_U3 ( .IN1(r838_n3), .IN2(r838_n4), .QN(r838_n1) );
  OR2X1 r838_U2 ( .IN2(r838_n4), .IN1(r838_n3), .Q(r838_n2) );
  NAND2X0 r838_U1 ( .IN1(r838_n1), .IN2(r838_n2), .QN(n105) );
  NAND2X0 r838_U182 ( .IN1(r838_n175), .IN2(r838_n176), .QN(r838_n32) );
  NAND2X0 r838_U181 ( .IN1(P2_N358), .IN2(r838_n32), .QN(r838_n172) );
  OR2X1 r838_U180 ( .IN2(P2_N358), .IN1(r838_n32), .Q(r838_n174) );
  NAND2X0 r838_U178 ( .IN1(r838_n174), .IN2(n18989), .QN(r838_n173) );
  NAND2X0 r838_U177 ( .IN1(r838_n172), .IN2(r838_n173), .QN(r838_n25) );
  NAND2X0 r838_U176 ( .IN1(P2_N357), .IN2(r838_n25), .QN(r838_n169) );
  OR2X1 r838_U175 ( .IN2(P2_N357), .IN1(r838_n25), .Q(r838_n171) );
  NAND2X0 r838_U173 ( .IN1(r838_n171), .IN2(n18987), .QN(r838_n170) );
  NAND2X0 r838_U172 ( .IN1(r838_n169), .IN2(r838_n170), .QN(r838_n18) );
  NAND2X0 r838_U171 ( .IN1(P2_N356), .IN2(r838_n18), .QN(r838_n166) );
  OR2X1 r838_U170 ( .IN2(P2_N356), .IN1(r838_n18), .Q(r838_n168) );
  NAND2X0 r838_U168 ( .IN1(r838_n168), .IN2(n18985), .QN(r838_n167) );
  NAND2X0 r838_U167 ( .IN1(r838_n166), .IN2(r838_n167), .QN(r838_n11) );
  NAND2X0 r838_U166 ( .IN1(P2_N355), .IN2(r838_n11), .QN(r838_n163) );
  OR2X1 r838_U165 ( .IN2(P2_N355), .IN1(r838_n11), .Q(r838_n165) );
  NAND2X0 r838_U163 ( .IN1(r838_n165), .IN2(n18983), .QN(r838_n164) );
  NAND2X0 r838_U162 ( .IN1(r838_n163), .IN2(r838_n164), .QN(r838_n4) );
  NAND2X0 r838_U161 ( .IN1(P2_N354), .IN2(r838_n4), .QN(r838_n160) );
  OR2X1 r838_U160 ( .IN2(P2_N354), .IN1(r838_n4), .Q(r838_n162) );
  NAND2X0 r838_U158 ( .IN1(r838_n162), .IN2(n18981), .QN(r838_n161) );
  NAND2X0 r838_U157 ( .IN1(r838_n160), .IN2(r838_n161), .QN(r838_n154) );
  NAND2X0 r838_U156 ( .IN1(r838_n159), .IN2(r838_n154), .QN(r838_n157) );
  OR2X1 r838_U155 ( .IN2(r838_n154), .IN1(r838_n159), .Q(r838_n158) );
  NAND2X0 r838_U154 ( .IN1(r838_n157), .IN2(r838_n158), .QN(n104) );
  NAND2X0 r838_U152 ( .IN1(P2_N352), .IN2(n18977), .QN(r838_n155) );
  OR2X1 r838_U151 ( .IN2(P2_N352), .IN1(n18977), .Q(r838_n156) );
  NAND2X0 r838_U150 ( .IN1(r838_n155), .IN2(r838_n156), .QN(r838_n149) );
  NAND2X0 r838_U149 ( .IN1(P2_N353), .IN2(r838_n154), .QN(r838_n150) );
  OR2X1 r838_U148 ( .IN2(P2_N353), .IN1(r838_n154), .Q(r838_n152) );
  NAND2X0 r838_U147 ( .IN1(r838_n152), .IN2(n18979), .QN(r838_n151) );
  NAND2X0 r838_U146 ( .IN1(r838_n150), .IN2(r838_n151), .QN(r838_n144) );
  NAND2X0 r838_U145 ( .IN1(r838_n149), .IN2(r838_n144), .QN(r838_n147) );
  OR2X1 r838_U144 ( .IN2(r838_n144), .IN1(r838_n149), .Q(r838_n148) );
  NAND2X0 r838_U143 ( .IN1(r838_n147), .IN2(r838_n148), .QN(n103) );
  NAND2X0 r838_U141 ( .IN1(P2_N351), .IN2(n18975), .QN(r838_n145) );
  OR2X1 r838_U140 ( .IN2(P2_N351), .IN1(n18975), .Q(r838_n146) );
  NAND2X0 r838_U139 ( .IN1(r838_n145), .IN2(r838_n146), .QN(r838_n139) );
  NAND2X0 r838_U138 ( .IN1(P2_N352), .IN2(r838_n144), .QN(r838_n140) );
  OR2X1 r838_U137 ( .IN2(P2_N352), .IN1(r838_n144), .Q(r838_n142) );
  NAND2X0 r838_U136 ( .IN1(r838_n142), .IN2(n18977), .QN(r838_n141) );
  NAND2X0 r838_U135 ( .IN1(r838_n140), .IN2(r838_n141), .QN(r838_n134) );
  NAND2X0 r838_U134 ( .IN1(r838_n139), .IN2(r838_n134), .QN(r838_n137) );
  OR2X1 r838_U133 ( .IN2(r838_n134), .IN1(r838_n139), .Q(r838_n138) );
  NAND2X0 r838_U132 ( .IN1(r838_n137), .IN2(r838_n138), .QN(n102) );
  NAND2X0 r838_U130 ( .IN1(P2_N350), .IN2(n18973), .QN(r838_n135) );
  OR2X1 r838_U129 ( .IN2(P2_N350), .IN1(n18973), .Q(r838_n136) );
  NAND2X0 r838_U128 ( .IN1(r838_n135), .IN2(r838_n136), .QN(r838_n129) );
  NAND2X0 r838_U127 ( .IN1(P2_N351), .IN2(r838_n134), .QN(r838_n130) );
  OR2X1 r838_U126 ( .IN2(P2_N351), .IN1(r838_n134), .Q(r838_n132) );
  NAND2X0 r838_U125 ( .IN1(r838_n132), .IN2(n18975), .QN(r838_n131) );
  NAND2X0 r838_U124 ( .IN1(r838_n130), .IN2(r838_n131), .QN(r838_n124) );
  NAND2X0 r838_U123 ( .IN1(r838_n129), .IN2(r838_n124), .QN(r838_n127) );
  OR2X1 r838_U122 ( .IN2(r838_n124), .IN1(r838_n129), .Q(r838_n128) );
  NAND2X0 r838_U121 ( .IN1(r838_n127), .IN2(r838_n128), .QN(n101) );
  NAND2X0 r838_U119 ( .IN1(P2_N349), .IN2(n18971), .QN(r838_n125) );
  OR2X1 r838_U118 ( .IN2(P2_N349), .IN1(n18971), .Q(r838_n126) );
  NAND2X0 r838_U117 ( .IN1(r838_n125), .IN2(r838_n126), .QN(r838_n119) );
  NAND2X0 r838_U116 ( .IN1(P2_N350), .IN2(r838_n124), .QN(r838_n120) );
  OR2X1 r838_U115 ( .IN2(P2_N350), .IN1(r838_n124), .Q(r838_n122) );
  NAND2X0 r838_U114 ( .IN1(r838_n122), .IN2(n18973), .QN(r838_n121) );
  NAND2X0 r838_U113 ( .IN1(r838_n120), .IN2(r838_n121), .QN(r838_n114) );
  NAND2X0 r838_U112 ( .IN1(r838_n119), .IN2(r838_n114), .QN(r838_n117) );
  OR2X1 r838_U111 ( .IN2(r838_n114), .IN1(r838_n119), .Q(r838_n118) );
  NAND2X0 r838_U110 ( .IN1(r838_n117), .IN2(r838_n118), .QN(n100) );
  NAND2X0 r838_U108 ( .IN1(P2_N348), .IN2(n18969), .QN(r838_n115) );
  OR2X1 r838_U107 ( .IN2(P2_N348), .IN1(n18969), .Q(r838_n116) );
  NAND2X0 r838_U106 ( .IN1(r838_n115), .IN2(r838_n116), .QN(r838_n109) );
  NAND2X0 r838_U105 ( .IN1(P2_N349), .IN2(r838_n114), .QN(r838_n110) );
  OR2X1 r838_U104 ( .IN2(P2_N349), .IN1(r838_n114), .Q(r838_n112) );
  NAND2X0 r838_U103 ( .IN1(r838_n112), .IN2(n18971), .QN(r838_n111) );
  NAND2X0 r838_U102 ( .IN1(r838_n110), .IN2(r838_n111), .QN(r838_n104) );
  NAND2X0 r838_U101 ( .IN1(r838_n109), .IN2(r838_n104), .QN(r838_n107) );
  OR2X1 r838_U100 ( .IN2(r838_n104), .IN1(r838_n109), .Q(r838_n108) );
  NAND2X0 r838_U99 ( .IN1(r838_n107), .IN2(r838_n108), .QN(n99) );
  NAND2X0 r838_U97 ( .IN1(P2_N347), .IN2(n18967), .QN(r838_n105) );
  OR2X1 r838_U96 ( .IN2(P2_N347), .IN1(n18967), .Q(r838_n106) );
  NAND2X0 r838_U95 ( .IN1(r838_n105), .IN2(r838_n106), .QN(r838_n99) );
  NAND2X0 r838_U94 ( .IN1(P2_N348), .IN2(r838_n104), .QN(r838_n100) );
  OR2X1 r838_U93 ( .IN2(P2_N348), .IN1(r838_n104), .Q(r838_n102) );
  NAND2X0 r838_U92 ( .IN1(r838_n102), .IN2(n18969), .QN(r838_n101) );
  NAND2X0 r838_U91 ( .IN1(r838_n100), .IN2(r838_n101), .QN(r838_n94) );
  NAND2X0 r838_U90 ( .IN1(r838_n99), .IN2(r838_n94), .QN(r838_n97) );
  INVX0 r838_U211 ( .ZN(r838_n191), .INP(n9843) );
  NOR2X0 r838_U210 ( .QN(r838_n187), .IN1(r838_n191), .IN2(P2_N363) );
  INVX0 r838_U209 ( .ZN(r838_n60), .INP(r838_n187) );
  NAND2X0 r838_U208 ( .IN1(P2_N363), .IN2(r838_n191), .QN(r838_n190) );
  NAND2X0 r838_U207 ( .IN1(r838_n60), .IN2(r838_n190), .QN(n114) );
  NAND2X0 r838_U205 ( .IN1(P2_N353), .IN2(n18979), .QN(r838_n188) );
  OR2X1 r838_U204 ( .IN2(P2_N353), .IN1(n18979), .Q(r838_n189) );
  NAND2X0 r838_U203 ( .IN1(r838_n188), .IN2(r838_n189), .QN(r838_n159) );
  NAND2X0 r838_U202 ( .IN1(P2_N362), .IN2(r838_n60), .QN(r838_n184) );
  NAND2X0 r838_U200 ( .IN1(r838_n187), .IN2(n6733), .QN(r838_n186) );
  NAND2X0 r838_U198 ( .IN1(r838_n186), .IN2(n18997), .QN(r838_n185) );
  NAND2X0 r838_U197 ( .IN1(r838_n184), .IN2(r838_n185), .QN(r838_n53) );
  NAND2X0 r838_U196 ( .IN1(P2_N361), .IN2(r838_n53), .QN(r838_n181) );
  OR2X1 r838_U195 ( .IN2(P2_N361), .IN1(r838_n53), .Q(r838_n183) );
  NAND2X0 r838_U193 ( .IN1(r838_n183), .IN2(n18995), .QN(r838_n182) );
  NAND2X0 r838_U192 ( .IN1(r838_n181), .IN2(r838_n182), .QN(r838_n46) );
  NAND2X0 r838_U191 ( .IN1(P2_N360), .IN2(r838_n46), .QN(r838_n178) );
  OR2X1 r838_U190 ( .IN2(P2_N360), .IN1(r838_n46), .Q(r838_n180) );
  NAND2X0 r838_U188 ( .IN1(r838_n180), .IN2(n18993), .QN(r838_n179) );
  NAND2X0 r838_U187 ( .IN1(r838_n178), .IN2(r838_n179), .QN(r838_n39) );
  NAND2X0 r838_U186 ( .IN1(P2_N359), .IN2(r838_n39), .QN(r838_n175) );
  OR2X1 r838_U185 ( .IN2(P2_N359), .IN1(r838_n39), .Q(r838_n177) );
  NAND2X0 r838_U183 ( .IN1(r838_n177), .IN2(n18991), .QN(r838_n176) );
  OR2X1 P2_sub_632_U77 ( .IN2(n9545), .IN1(P2_sub_632_n9), .Q(P2_sub_632_n7)
         );
  OR2X1 P2_sub_632_U76 ( .IN2(n9541), .IN1(P2_sub_632_n7), .Q(P2_sub_632_n5)
         );
  OR2X1 P2_sub_632_U75 ( .IN2(n9537), .IN1(P2_sub_632_n5), .Q(P2_sub_632_n53)
         );
  NAND2X0 P2_sub_632_U74 ( .IN1(n9537), .IN2(P2_sub_632_n5), 
        .QN(P2_sub_632_n54) );
  NAND2X0 P2_sub_632_U73 ( .IN1(P2_sub_632_n53), .IN2(P2_sub_632_n54), 
        .QN(P2_N374) );
  OR2X1 P2_sub_632_U72 ( .IN2(n9533), .IN1(P2_sub_632_n53), .Q(P2_sub_632_n51)
         );
  NAND2X0 P2_sub_632_U71 ( .IN1(n9533), .IN2(P2_sub_632_n53), 
        .QN(P2_sub_632_n52) );
  NAND2X0 P2_sub_632_U70 ( .IN1(P2_sub_632_n51), .IN2(P2_sub_632_n52), 
        .QN(P2_N375) );
  OR2X1 P2_sub_632_U69 ( .IN2(n9529), .IN1(P2_sub_632_n51), .Q(P2_sub_632_n49)
         );
  NAND2X0 P2_sub_632_U68 ( .IN1(n9529), .IN2(P2_sub_632_n51), 
        .QN(P2_sub_632_n50) );
  NAND2X0 P2_sub_632_U67 ( .IN1(P2_sub_632_n49), .IN2(P2_sub_632_n50), 
        .QN(P2_N376) );
  OR2X1 P2_sub_632_U66 ( .IN2(n9525), .IN1(P2_sub_632_n49), .Q(P2_sub_632_n47)
         );
  NAND2X0 P2_sub_632_U65 ( .IN1(n9525), .IN2(P2_sub_632_n49), 
        .QN(P2_sub_632_n48) );
  NAND2X0 P2_sub_632_U64 ( .IN1(P2_sub_632_n47), .IN2(P2_sub_632_n48), 
        .QN(P2_N377) );
  OR2X1 P2_sub_632_U63 ( .IN2(n9521), .IN1(P2_sub_632_n47), .Q(P2_sub_632_n45)
         );
  NAND2X0 P2_sub_632_U62 ( .IN1(n9521), .IN2(P2_sub_632_n47), 
        .QN(P2_sub_632_n46) );
  NAND2X0 P2_sub_632_U61 ( .IN1(P2_sub_632_n45), .IN2(P2_sub_632_n46), 
        .QN(P2_N378) );
  OR2X1 P2_sub_632_U60 ( .IN2(n9517), .IN1(P2_sub_632_n45), .Q(P2_sub_632_n43)
         );
  NAND2X0 P2_sub_632_U59 ( .IN1(n9517), .IN2(P2_sub_632_n45), 
        .QN(P2_sub_632_n44) );
  NAND2X0 P2_sub_632_U58 ( .IN1(P2_sub_632_n43), .IN2(P2_sub_632_n44), 
        .QN(P2_N379) );
  OR2X1 P2_sub_632_U57 ( .IN2(n9513), .IN1(P2_sub_632_n43), .Q(P2_sub_632_n41)
         );
  NAND2X0 P2_sub_632_U56 ( .IN1(n9513), .IN2(P2_sub_632_n43), 
        .QN(P2_sub_632_n42) );
  NAND2X0 P2_sub_632_U55 ( .IN1(P2_sub_632_n41), .IN2(P2_sub_632_n42), 
        .QN(P2_N380) );
  OR2X1 P2_sub_632_U54 ( .IN2(n9509), .IN1(P2_sub_632_n41), .Q(P2_sub_632_n39)
         );
  NAND2X0 P2_sub_632_U53 ( .IN1(n9509), .IN2(P2_sub_632_n41), 
        .QN(P2_sub_632_n40) );
  NAND2X0 P2_sub_632_U52 ( .IN1(P2_sub_632_n39), .IN2(P2_sub_632_n40), 
        .QN(P2_N381) );
  OR2X1 P2_sub_632_U51 ( .IN2(n9505), .IN1(P2_sub_632_n39), .Q(P2_sub_632_n37)
         );
  NAND2X0 P2_sub_632_U50 ( .IN1(n9505), .IN2(P2_sub_632_n39), 
        .QN(P2_sub_632_n38) );
  NAND2X0 P2_sub_632_U49 ( .IN1(P2_sub_632_n37), .IN2(P2_sub_632_n38), 
        .QN(P2_N382) );
  OR2X1 P2_sub_632_U48 ( .IN2(n9501), .IN1(P2_sub_632_n37), .Q(P2_sub_632_n35)
         );
  NAND2X0 P2_sub_632_U47 ( .IN1(n9501), .IN2(P2_sub_632_n37), 
        .QN(P2_sub_632_n36) );
  NAND2X0 P2_sub_632_U46 ( .IN1(P2_sub_632_n35), .IN2(P2_sub_632_n36), 
        .QN(P2_N383) );
  OR2X1 P2_sub_632_U45 ( .IN2(n9381), .IN1(P2_sub_632_n35), .Q(P2_sub_632_n33)
         );
  NAND2X0 P2_sub_632_U44 ( .IN1(n9381), .IN2(P2_sub_632_n35), 
        .QN(P2_sub_632_n34) );
  NAND2X0 P2_sub_632_U43 ( .IN1(P2_sub_632_n33), .IN2(P2_sub_632_n34), 
        .QN(P2_N384) );
  OR2X1 P2_sub_632_U42 ( .IN2(n9377), .IN1(P2_sub_632_n33), .Q(P2_sub_632_n31)
         );
  NAND2X0 P2_sub_632_U41 ( .IN1(n9377), .IN2(P2_sub_632_n33), 
        .QN(P2_sub_632_n32) );
  NAND2X0 P2_sub_632_U40 ( .IN1(P2_sub_632_n31), .IN2(P2_sub_632_n32), 
        .QN(P2_N385) );
  OR2X1 P2_sub_632_U39 ( .IN2(n9373), .IN1(P2_sub_632_n31), .Q(P2_sub_632_n29)
         );
  NAND2X0 P2_sub_632_U38 ( .IN1(n9373), .IN2(P2_sub_632_n31), 
        .QN(P2_sub_632_n30) );
  NAND2X0 P2_sub_632_U37 ( .IN1(P2_sub_632_n29), .IN2(P2_sub_632_n30), 
        .QN(P2_N386) );
  OR2X1 P2_sub_632_U36 ( .IN2(n9369), .IN1(P2_sub_632_n29), .Q(P2_sub_632_n27)
         );
  NAND2X0 P2_sub_632_U35 ( .IN1(n9369), .IN2(P2_sub_632_n29), 
        .QN(P2_sub_632_n28) );
  NAND2X0 P2_sub_632_U34 ( .IN1(P2_sub_632_n27), .IN2(P2_sub_632_n28), 
        .QN(P2_N387) );
  OR2X1 P2_sub_632_U33 ( .IN2(n9365), .IN1(P2_sub_632_n27), .Q(P2_sub_632_n25)
         );
  NAND2X0 P2_sub_632_U32 ( .IN1(n9365), .IN2(P2_sub_632_n27), 
        .QN(P2_sub_632_n26) );
  NAND2X0 P2_sub_632_U31 ( .IN1(P2_sub_632_n25), .IN2(P2_sub_632_n26), 
        .QN(P2_N388) );
  OR2X1 P2_sub_632_U30 ( .IN2(n9361), .IN1(P2_sub_632_n25), .Q(P2_sub_632_n23)
         );
  NAND2X0 P2_sub_632_U29 ( .IN1(n9361), .IN2(P2_sub_632_n25), 
        .QN(P2_sub_632_n24) );
  NAND2X0 P2_sub_632_U28 ( .IN1(P2_sub_632_n23), .IN2(P2_sub_632_n24), 
        .QN(P2_N389) );
  OR2X1 P2_sub_632_U27 ( .IN2(n9357), .IN1(P2_sub_632_n23), .Q(P2_sub_632_n21)
         );
  NAND2X0 P2_sub_632_U26 ( .IN1(n9357), .IN2(P2_sub_632_n23), 
        .QN(P2_sub_632_n22) );
  NAND2X0 P2_sub_632_U25 ( .IN1(P2_sub_632_n21), .IN2(P2_sub_632_n22), 
        .QN(P2_N390) );
  OR2X1 P2_sub_632_U24 ( .IN2(n9353), .IN1(P2_sub_632_n21), .Q(P2_sub_632_n19)
         );
  NAND2X0 P2_sub_632_U23 ( .IN1(n9353), .IN2(P2_sub_632_n21), 
        .QN(P2_sub_632_n20) );
  NAND2X0 P2_sub_632_U22 ( .IN1(P2_sub_632_n19), .IN2(P2_sub_632_n20), 
        .QN(P2_N391) );
  NOR2X0 P2_sub_632_U21 ( .QN(P2_N394), .IN1(P2_sub_632_n19), .IN2(n9349) );
  INVX0 P2_sub_632_U20 ( .ZN(P2_sub_632_n17), .INP(P2_N394) );
  NAND2X0 P2_sub_632_U19 ( .IN1(n9349), .IN2(P2_sub_632_n19), 
        .QN(P2_sub_632_n18) );
  NAND2X0 P2_sub_632_U18 ( .IN1(P2_sub_632_n17), .IN2(P2_sub_632_n18), 
        .QN(P2_N392) );
  NAND2X0 P2_sub_632_U16 ( .IN1(n9397), .IN2(n6684), .QN(P2_sub_632_n16) );
  NAND2X0 P2_sub_632_U15 ( .IN1(P2_sub_632_n15), .IN2(P2_sub_632_n16), 
        .QN(P2_N368) );
  NAND2X0 P2_sub_632_U14 ( .IN1(n9557), .IN2(P2_sub_632_n15), 
        .QN(P2_sub_632_n14) );
  NAND2X0 P2_sub_632_U13 ( .IN1(P2_sub_632_n13), .IN2(P2_sub_632_n14), 
        .QN(P2_N369) );
  NAND2X0 P2_sub_632_U12 ( .IN1(n9553), .IN2(P2_sub_632_n13), 
        .QN(P2_sub_632_n12) );
  NAND2X0 P2_sub_632_U11 ( .IN1(P2_sub_632_n11), .IN2(P2_sub_632_n12), 
        .QN(P2_N370) );
  NAND2X0 P2_sub_632_U10 ( .IN1(n9549), .IN2(P2_sub_632_n11), 
        .QN(P2_sub_632_n10) );
  NAND2X0 P2_sub_632_U9 ( .IN1(P2_sub_632_n9), .IN2(P2_sub_632_n10), 
        .QN(P2_N371) );
  NAND2X0 P2_sub_632_U8 ( .IN1(n9545), .IN2(P2_sub_632_n9), .QN(P2_sub_632_n8)
         );
  NAND2X0 P2_sub_632_U7 ( .IN1(P2_sub_632_n7), .IN2(P2_sub_632_n8), 
        .QN(P2_N372) );
  NAND2X0 P2_sub_632_U6 ( .IN1(n9541), .IN2(P2_sub_632_n7), .QN(P2_sub_632_n6)
         );
  NAND2X0 P2_sub_632_U5 ( .IN1(P2_sub_632_n5), .IN2(P2_sub_632_n6), 
        .QN(P2_N373) );
  NBUFFX2 P2_sub_632_U1 ( .INP(P2_N394), .Z(P2_N393) );
  OR2X1 P2_sub_632_U81 ( .IN2(n6684), .IN1(n9397), .Q(P2_sub_632_n15) );
  OR2X1 P2_sub_632_U80 ( .IN2(n9557), .IN1(P2_sub_632_n15), .Q(P2_sub_632_n13)
         );
  OR2X1 P2_sub_632_U79 ( .IN2(n9553), .IN1(P2_sub_632_n13), .Q(P2_sub_632_n11)
         );
  OR2X1 P2_sub_632_U78 ( .IN2(n9549), .IN1(P2_sub_632_n11), .Q(P2_sub_632_n9)
         );
  NAND2X0 add_1108_U335 ( .IN1(add_1108_n184), .IN2(add_1108_n181), 
        .QN(add_1108_n307) );
  OR2X1 add_1108_U336 ( .IN2(add_1108_n181), .IN1(add_1108_n184), 
        .Q(add_1108_n305) );
  NAND2X0 add_1108_U337 ( .IN1(si_0_), .IN2(n9385), .QN(add_1108_n181) );
  INVX0 add_1108_U338 ( .ZN(add_1108_n184), .INP(n9333) );
  NAND2X0 add_1108_U339 ( .IN1(add_1108_n308), .IN2(add_1108_n309), .QN(N39)
         );
  NAND2X0 add_1108_U340 ( .IN1(si_0_), .IN2(add_1108_n310), .QN(add_1108_n309)
         );
  OR2X1 add_1108_U341 ( .IN2(si_0_), .IN1(add_1108_n310), .Q(add_1108_n308) );
  INVX0 add_1108_U342 ( .ZN(add_1108_n310), .INP(n9385) );
  OR2X1 add_1108_U327 ( .IN2(n9895), .IN1(add_1108_n45), .Q(add_1108_n301) );
  NAND2X0 add_1108_U328 ( .IN1(n9895), .IN2(add_1108_n45), .QN(add_1108_n299)
         );
  NAND2X0 add_1108_U329 ( .IN1(add_1108_n302), .IN2(add_1108_n303), 
        .QN(add_1108_n45) );
  NAND2X0 add_1108_U330 ( .IN1(si_2_), .IN2(add_1108_n304), .QN(add_1108_n303)
         );
  OR2X1 add_1108_U331 ( .IN2(n9899), .IN1(add_1108_n73), .Q(add_1108_n304) );
  NAND2X0 add_1108_U332 ( .IN1(n9899), .IN2(add_1108_n73), .QN(add_1108_n302)
         );
  NAND2X0 add_1108_U333 ( .IN1(add_1108_n305), .IN2(add_1108_n306), 
        .QN(add_1108_n73) );
  NAND2X0 add_1108_U334 ( .IN1(si_1_), .IN2(add_1108_n307), .QN(add_1108_n306)
         );
  OR2X1 add_1108_U319 ( .IN2(n9887), .IN1(add_1108_n31), .Q(add_1108_n295) );
  NAND2X0 add_1108_U320 ( .IN1(n9887), .IN2(add_1108_n31), .QN(add_1108_n293)
         );
  NAND2X0 add_1108_U321 ( .IN1(add_1108_n296), .IN2(add_1108_n297), 
        .QN(add_1108_n31) );
  NAND2X0 add_1108_U322 ( .IN1(si_4_), .IN2(add_1108_n298), .QN(add_1108_n297)
         );
  OR2X1 add_1108_U323 ( .IN2(n9891), .IN1(add_1108_n38), .Q(add_1108_n298) );
  NAND2X0 add_1108_U324 ( .IN1(n9891), .IN2(add_1108_n38), .QN(add_1108_n296)
         );
  NAND2X0 add_1108_U325 ( .IN1(add_1108_n299), .IN2(add_1108_n300), 
        .QN(add_1108_n38) );
  NAND2X0 add_1108_U326 ( .IN1(si_3_), .IN2(add_1108_n301), .QN(add_1108_n300)
         );
  OR2X1 add_1108_U311 ( .IN2(n9879), .IN1(add_1108_n17), .Q(add_1108_n289) );
  NAND2X0 add_1108_U312 ( .IN1(n9879), .IN2(add_1108_n17), .QN(add_1108_n287)
         );
  NAND2X0 add_1108_U313 ( .IN1(add_1108_n290), .IN2(add_1108_n291), 
        .QN(add_1108_n17) );
  NAND2X0 add_1108_U314 ( .IN1(si_6_), .IN2(add_1108_n292), .QN(add_1108_n291)
         );
  OR2X1 add_1108_U315 ( .IN2(n9883), .IN1(add_1108_n24), .Q(add_1108_n292) );
  NAND2X0 add_1108_U316 ( .IN1(n9883), .IN2(add_1108_n24), .QN(add_1108_n290)
         );
  NAND2X0 add_1108_U317 ( .IN1(add_1108_n293), .IN2(add_1108_n294), 
        .QN(add_1108_n24) );
  NAND2X0 add_1108_U318 ( .IN1(si_5_), .IN2(add_1108_n295), .QN(add_1108_n294)
         );
  OR2X1 add_1108_U303 ( .IN2(n9871), .IN1(add_1108_n3), .Q(add_1108_n283) );
  NAND2X0 add_1108_U304 ( .IN1(n9871), .IN2(add_1108_n3), .QN(add_1108_n281)
         );
  NAND2X0 add_1108_U305 ( .IN1(add_1108_n284), .IN2(add_1108_n285), 
        .QN(add_1108_n3) );
  NAND2X0 add_1108_U306 ( .IN1(si_8_), .IN2(add_1108_n286), .QN(add_1108_n285)
         );
  OR2X1 add_1108_U307 ( .IN2(n9875), .IN1(add_1108_n10), .Q(add_1108_n286) );
  NAND2X0 add_1108_U308 ( .IN1(n9875), .IN2(add_1108_n10), .QN(add_1108_n284)
         );
  NAND2X0 add_1108_U309 ( .IN1(add_1108_n287), .IN2(add_1108_n288), 
        .QN(add_1108_n10) );
  NAND2X0 add_1108_U310 ( .IN1(si_7_), .IN2(add_1108_n289), .QN(add_1108_n288)
         );
  AND2X1 add_1108_U295 ( .IN1(add_1108_n274), .IN2(add_1108_n277), 
        .Q(add_1108_n276) );
  NOR2X0 add_1108_U296 ( .QN(add_1108_n275), .IN1(add_1108_n274), 
        .IN2(add_1108_n277) );
  NAND2X0 add_1108_U297 ( .IN1(add_1108_n278), .IN2(add_1108_n279), 
        .QN(add_1108_n277) );
  NAND2X0 add_1108_U298 ( .IN1(si_10_), .IN2(add_1108_n280), 
        .QN(add_1108_n279) );
  OR2X1 add_1108_U299 ( .IN2(si_10_), .IN1(add_1108_n280), .Q(add_1108_n278)
         );
  INVX0 add_1108_U300 ( .ZN(add_1108_n280), .INP(n10007) );
  NAND2X0 add_1108_U301 ( .IN1(add_1108_n281), .IN2(add_1108_n282), 
        .QN(add_1108_n274) );
  NAND2X0 add_1108_U302 ( .IN1(si_9_), .IN2(add_1108_n283), .QN(add_1108_n282)
         );
  NAND2X0 add_1108_U287 ( .IN1(si_11_), .IN2(add_1108_n270), 
        .QN(add_1108_n269) );
  OR2X1 add_1108_U288 ( .IN2(si_11_), .IN1(add_1108_n270), .Q(add_1108_n268)
         );
  INVX0 add_1108_U289 ( .ZN(add_1108_n270), .INP(n10003) );
  NAND2X0 add_1108_U290 ( .IN1(add_1108_n271), .IN2(add_1108_n272), 
        .QN(add_1108_n264) );
  NAND2X0 add_1108_U291 ( .IN1(si_10_), .IN2(add_1108_n273), 
        .QN(add_1108_n272) );
  OR2X1 add_1108_U292 ( .IN2(n10007), .IN1(add_1108_n274), .Q(add_1108_n273)
         );
  NAND2X0 add_1108_U293 ( .IN1(n10007), .IN2(add_1108_n274), 
        .QN(add_1108_n271) );
  NOR2X0 add_1108_U294 ( .QN(N49), .IN1(add_1108_n275), .IN2(add_1108_n276) );
  NAND2X0 add_1108_U279 ( .IN1(add_1108_n261), .IN2(add_1108_n262), 
        .QN(add_1108_n254) );
  NAND2X0 add_1108_U280 ( .IN1(si_11_), .IN2(add_1108_n263), 
        .QN(add_1108_n262) );
  OR2X1 add_1108_U281 ( .IN2(n10003), .IN1(add_1108_n264), .Q(add_1108_n263)
         );
  NAND2X0 add_1108_U282 ( .IN1(n10003), .IN2(add_1108_n264), 
        .QN(add_1108_n261) );
  NOR2X0 add_1108_U283 ( .QN(N50), .IN1(add_1108_n265), .IN2(add_1108_n266) );
  AND2X1 add_1108_U284 ( .IN1(add_1108_n264), .IN2(add_1108_n267), 
        .Q(add_1108_n266) );
  NOR2X0 add_1108_U285 ( .QN(add_1108_n265), .IN1(add_1108_n264), 
        .IN2(add_1108_n267) );
  NAND2X0 add_1108_U286 ( .IN1(add_1108_n268), .IN2(add_1108_n269), 
        .QN(add_1108_n267) );
  NAND2X0 add_1108_U271 ( .IN1(n9999), .IN2(add_1108_n254), .QN(add_1108_n251)
         );
  NOR2X0 add_1108_U272 ( .QN(N51), .IN1(add_1108_n255), .IN2(add_1108_n256) );
  AND2X1 add_1108_U273 ( .IN1(add_1108_n254), .IN2(add_1108_n257), 
        .Q(add_1108_n256) );
  NOR2X0 add_1108_U274 ( .QN(add_1108_n255), .IN1(add_1108_n254), 
        .IN2(add_1108_n257) );
  NAND2X0 add_1108_U275 ( .IN1(add_1108_n258), .IN2(add_1108_n259), 
        .QN(add_1108_n257) );
  NAND2X0 add_1108_U276 ( .IN1(si_12_), .IN2(add_1108_n260), 
        .QN(add_1108_n259) );
  OR2X1 add_1108_U277 ( .IN2(si_12_), .IN1(add_1108_n260), .Q(add_1108_n258)
         );
  INVX0 add_1108_U278 ( .ZN(add_1108_n260), .INP(n9999) );
  NOR2X0 add_1108_U263 ( .QN(add_1108_n245), .IN1(add_1108_n244), 
        .IN2(add_1108_n247) );
  NAND2X0 add_1108_U264 ( .IN1(add_1108_n248), .IN2(add_1108_n249), 
        .QN(add_1108_n247) );
  NAND2X0 add_1108_U265 ( .IN1(si_13_), .IN2(add_1108_n250), 
        .QN(add_1108_n249) );
  OR2X1 add_1108_U266 ( .IN2(si_13_), .IN1(add_1108_n250), .Q(add_1108_n248)
         );
  INVX0 add_1108_U267 ( .ZN(add_1108_n250), .INP(n9995) );
  NAND2X0 add_1108_U268 ( .IN1(add_1108_n251), .IN2(add_1108_n252), 
        .QN(add_1108_n244) );
  NAND2X0 add_1108_U269 ( .IN1(si_12_), .IN2(add_1108_n253), 
        .QN(add_1108_n252) );
  OR2X1 add_1108_U270 ( .IN2(n9999), .IN1(add_1108_n254), .Q(add_1108_n253) );
  OR2X1 add_1108_U255 ( .IN2(si_14_), .IN1(add_1108_n240), .Q(add_1108_n238)
         );
  INVX0 add_1108_U256 ( .ZN(add_1108_n240), .INP(n9991) );
  NAND2X0 add_1108_U257 ( .IN1(add_1108_n241), .IN2(add_1108_n242), 
        .QN(add_1108_n234) );
  NAND2X0 add_1108_U258 ( .IN1(si_13_), .IN2(add_1108_n243), 
        .QN(add_1108_n242) );
  OR2X1 add_1108_U259 ( .IN2(n9995), .IN1(add_1108_n244), .Q(add_1108_n243) );
  NAND2X0 add_1108_U260 ( .IN1(n9995), .IN2(add_1108_n244), .QN(add_1108_n241)
         );
  NOR2X0 add_1108_U261 ( .QN(N52), .IN1(add_1108_n245), .IN2(add_1108_n246) );
  AND2X1 add_1108_U262 ( .IN1(add_1108_n244), .IN2(add_1108_n247), 
        .Q(add_1108_n246) );
  NAND2X0 add_1108_U247 ( .IN1(si_14_), .IN2(add_1108_n233), 
        .QN(add_1108_n232) );
  OR2X1 add_1108_U248 ( .IN2(n9991), .IN1(add_1108_n234), .Q(add_1108_n233) );
  NAND2X0 add_1108_U249 ( .IN1(n9991), .IN2(add_1108_n234), .QN(add_1108_n231)
         );
  NOR2X0 add_1108_U250 ( .QN(N53), .IN1(add_1108_n235), .IN2(add_1108_n236) );
  AND2X1 add_1108_U251 ( .IN1(add_1108_n234), .IN2(add_1108_n237), 
        .Q(add_1108_n236) );
  NOR2X0 add_1108_U252 ( .QN(add_1108_n235), .IN1(add_1108_n234), 
        .IN2(add_1108_n237) );
  NAND2X0 add_1108_U253 ( .IN1(add_1108_n238), .IN2(add_1108_n239), 
        .QN(add_1108_n237) );
  NAND2X0 add_1108_U254 ( .IN1(si_14_), .IN2(add_1108_n240), 
        .QN(add_1108_n239) );
  NOR2X0 add_1108_U239 ( .QN(N54), .IN1(add_1108_n225), .IN2(add_1108_n226) );
  AND2X1 add_1108_U240 ( .IN1(add_1108_n224), .IN2(add_1108_n227), 
        .Q(add_1108_n226) );
  NOR2X0 add_1108_U241 ( .QN(add_1108_n225), .IN1(add_1108_n224), 
        .IN2(add_1108_n227) );
  NAND2X0 add_1108_U242 ( .IN1(add_1108_n228), .IN2(add_1108_n229), 
        .QN(add_1108_n227) );
  NAND2X0 add_1108_U243 ( .IN1(si_15_), .IN2(add_1108_n230), 
        .QN(add_1108_n229) );
  OR2X1 add_1108_U244 ( .IN2(si_15_), .IN1(add_1108_n230), .Q(add_1108_n228)
         );
  INVX0 add_1108_U245 ( .ZN(add_1108_n230), .INP(n9987) );
  NAND2X0 add_1108_U246 ( .IN1(add_1108_n231), .IN2(add_1108_n232), 
        .QN(add_1108_n224) );
  NAND2X0 add_1108_U231 ( .IN1(add_1108_n218), .IN2(add_1108_n219), 
        .QN(add_1108_n217) );
  NAND2X0 add_1108_U232 ( .IN1(si_16_), .IN2(add_1108_n220), 
        .QN(add_1108_n219) );
  OR2X1 add_1108_U233 ( .IN2(si_16_), .IN1(add_1108_n220), .Q(add_1108_n218)
         );
  INVX0 add_1108_U234 ( .ZN(add_1108_n220), .INP(n9983) );
  NAND2X0 add_1108_U235 ( .IN1(add_1108_n221), .IN2(add_1108_n222), 
        .QN(add_1108_n214) );
  NAND2X0 add_1108_U236 ( .IN1(si_15_), .IN2(add_1108_n223), 
        .QN(add_1108_n222) );
  OR2X1 add_1108_U237 ( .IN2(n9987), .IN1(add_1108_n224), .Q(add_1108_n223) );
  NAND2X0 add_1108_U238 ( .IN1(n9987), .IN2(add_1108_n224), .QN(add_1108_n221)
         );
  INVX0 add_1108_U223 ( .ZN(add_1108_n210), .INP(n9979) );
  NAND2X0 add_1108_U224 ( .IN1(add_1108_n211), .IN2(add_1108_n212), 
        .QN(add_1108_n204) );
  NAND2X0 add_1108_U225 ( .IN1(si_16_), .IN2(add_1108_n213), 
        .QN(add_1108_n212) );
  OR2X1 add_1108_U226 ( .IN2(n9983), .IN1(add_1108_n214), .Q(add_1108_n213) );
  NAND2X0 add_1108_U227 ( .IN1(n9983), .IN2(add_1108_n214), .QN(add_1108_n211)
         );
  NOR2X0 add_1108_U228 ( .QN(N55), .IN1(add_1108_n215), .IN2(add_1108_n216) );
  AND2X1 add_1108_U229 ( .IN1(add_1108_n214), .IN2(add_1108_n217), 
        .Q(add_1108_n216) );
  NOR2X0 add_1108_U230 ( .QN(add_1108_n215), .IN1(add_1108_n214), 
        .IN2(add_1108_n217) );
  OR2X1 add_1108_U215 ( .IN2(n9979), .IN1(add_1108_n204), .Q(add_1108_n203) );
  NAND2X0 add_1108_U216 ( .IN1(n9979), .IN2(add_1108_n204), .QN(add_1108_n201)
         );
  NOR2X0 add_1108_U217 ( .QN(N56), .IN1(add_1108_n205), .IN2(add_1108_n206) );
  AND2X1 add_1108_U218 ( .IN1(add_1108_n204), .IN2(add_1108_n207), 
        .Q(add_1108_n206) );
  NOR2X0 add_1108_U219 ( .QN(add_1108_n205), .IN1(add_1108_n204), 
        .IN2(add_1108_n207) );
  NAND2X0 add_1108_U220 ( .IN1(add_1108_n208), .IN2(add_1108_n209), 
        .QN(add_1108_n207) );
  NAND2X0 add_1108_U221 ( .IN1(si_17_), .IN2(add_1108_n210), 
        .QN(add_1108_n209) );
  OR2X1 add_1108_U222 ( .IN2(si_17_), .IN1(add_1108_n210), .Q(add_1108_n208)
         );
  AND2X1 add_1108_U207 ( .IN1(add_1108_n194), .IN2(add_1108_n197), 
        .Q(add_1108_n196) );
  NOR2X0 add_1108_U208 ( .QN(add_1108_n195), .IN1(add_1108_n194), 
        .IN2(add_1108_n197) );
  NAND2X0 add_1108_U209 ( .IN1(add_1108_n198), .IN2(add_1108_n199), 
        .QN(add_1108_n197) );
  NAND2X0 add_1108_U210 ( .IN1(si_18_), .IN2(add_1108_n200), 
        .QN(add_1108_n199) );
  OR2X1 add_1108_U211 ( .IN2(si_18_), .IN1(add_1108_n200), .Q(add_1108_n198)
         );
  INVX0 add_1108_U212 ( .ZN(add_1108_n200), .INP(n9975) );
  NAND2X0 add_1108_U213 ( .IN1(add_1108_n201), .IN2(add_1108_n202), 
        .QN(add_1108_n194) );
  NAND2X0 add_1108_U214 ( .IN1(si_17_), .IN2(add_1108_n203), 
        .QN(add_1108_n202) );
  NAND2X0 add_1108_U199 ( .IN1(si_19_), .IN2(add_1108_n190), 
        .QN(add_1108_n189) );
  OR2X1 add_1108_U200 ( .IN2(si_19_), .IN1(add_1108_n190), .Q(add_1108_n188)
         );
  INVX0 add_1108_U201 ( .ZN(add_1108_n190), .INP(n9971) );
  NAND2X0 add_1108_U202 ( .IN1(add_1108_n191), .IN2(add_1108_n192), 
        .QN(add_1108_n177) );
  NAND2X0 add_1108_U203 ( .IN1(si_18_), .IN2(add_1108_n193), 
        .QN(add_1108_n192) );
  OR2X1 add_1108_U204 ( .IN2(n9975), .IN1(add_1108_n194), .Q(add_1108_n193) );
  NAND2X0 add_1108_U205 ( .IN1(n9975), .IN2(add_1108_n194), .QN(add_1108_n191)
         );
  NOR2X0 add_1108_U206 ( .QN(N57), .IN1(add_1108_n195), .IN2(add_1108_n196) );
  NAND2X0 add_1108_U191 ( .IN1(add_1108_n180), .IN2(add_1108_n181), 
        .QN(add_1108_n178) );
  NAND2X0 add_1108_U192 ( .IN1(add_1108_n182), .IN2(add_1108_n183), 
        .QN(add_1108_n180) );
  NAND2X0 add_1108_U193 ( .IN1(si_1_), .IN2(add_1108_n184), .QN(add_1108_n183)
         );
  OR2X1 add_1108_U194 ( .IN2(si_1_), .IN1(add_1108_n184), .Q(add_1108_n182) );
  NOR2X0 add_1108_U195 ( .QN(N58), .IN1(add_1108_n185), .IN2(add_1108_n186) );
  AND2X1 add_1108_U196 ( .IN1(add_1108_n177), .IN2(add_1108_n187), 
        .Q(add_1108_n186) );
  NOR2X0 add_1108_U197 ( .QN(add_1108_n185), .IN1(add_1108_n177), 
        .IN2(add_1108_n187) );
  NAND2X0 add_1108_U198 ( .IN1(add_1108_n188), .IN2(add_1108_n189), 
        .QN(add_1108_n187) );
  OR2X1 add_1108_U183 ( .IN2(si_20_), .IN1(add_1108_n173), .Q(add_1108_n171)
         );
  INVX0 add_1108_U184 ( .ZN(add_1108_n173), .INP(n9967) );
  NAND2X0 add_1108_U185 ( .IN1(add_1108_n174), .IN2(add_1108_n175), 
        .QN(add_1108_n167) );
  NAND2X0 add_1108_U186 ( .IN1(si_19_), .IN2(add_1108_n176), 
        .QN(add_1108_n175) );
  OR2X1 add_1108_U187 ( .IN2(n9971), .IN1(add_1108_n177), .Q(add_1108_n176) );
  NAND2X0 add_1108_U188 ( .IN1(n9971), .IN2(add_1108_n177), .QN(add_1108_n174)
         );
  NAND2X0 add_1108_U189 ( .IN1(add_1108_n178), .IN2(add_1108_n179), .QN(N40)
         );
  OR2X1 add_1108_U190 ( .IN2(add_1108_n181), .IN1(add_1108_n180), 
        .Q(add_1108_n179) );
  NAND2X0 add_1108_U175 ( .IN1(si_20_), .IN2(add_1108_n166), 
        .QN(add_1108_n165) );
  OR2X1 add_1108_U176 ( .IN2(n9967), .IN1(add_1108_n167), .Q(add_1108_n166) );
  NAND2X0 add_1108_U177 ( .IN1(n9967), .IN2(add_1108_n167), .QN(add_1108_n164)
         );
  NOR2X0 add_1108_U178 ( .QN(N59), .IN1(add_1108_n168), .IN2(add_1108_n169) );
  AND2X1 add_1108_U179 ( .IN1(add_1108_n167), .IN2(add_1108_n170), 
        .Q(add_1108_n169) );
  NOR2X0 add_1108_U180 ( .QN(add_1108_n168), .IN1(add_1108_n167), 
        .IN2(add_1108_n170) );
  NAND2X0 add_1108_U181 ( .IN1(add_1108_n171), .IN2(add_1108_n172), 
        .QN(add_1108_n170) );
  NAND2X0 add_1108_U182 ( .IN1(si_20_), .IN2(add_1108_n173), 
        .QN(add_1108_n172) );
  NOR2X0 add_1108_U167 ( .QN(N60), .IN1(add_1108_n158), .IN2(add_1108_n159) );
  AND2X1 add_1108_U168 ( .IN1(add_1108_n157), .IN2(add_1108_n160), 
        .Q(add_1108_n159) );
  NOR2X0 add_1108_U169 ( .QN(add_1108_n158), .IN1(add_1108_n157), 
        .IN2(add_1108_n160) );
  NAND2X0 add_1108_U170 ( .IN1(add_1108_n161), .IN2(add_1108_n162), 
        .QN(add_1108_n160) );
  NAND2X0 add_1108_U171 ( .IN1(si_21_), .IN2(add_1108_n163), 
        .QN(add_1108_n162) );
  OR2X1 add_1108_U172 ( .IN2(si_21_), .IN1(add_1108_n163), .Q(add_1108_n161)
         );
  INVX0 add_1108_U173 ( .ZN(add_1108_n163), .INP(n9963) );
  NAND2X0 add_1108_U174 ( .IN1(add_1108_n164), .IN2(add_1108_n165), 
        .QN(add_1108_n157) );
  NAND2X0 add_1108_U159 ( .IN1(add_1108_n151), .IN2(add_1108_n152), 
        .QN(add_1108_n150) );
  NAND2X0 add_1108_U160 ( .IN1(si_22_), .IN2(add_1108_n153), 
        .QN(add_1108_n152) );
  OR2X1 add_1108_U161 ( .IN2(si_22_), .IN1(add_1108_n153), .Q(add_1108_n151)
         );
  INVX0 add_1108_U162 ( .ZN(add_1108_n153), .INP(n9959) );
  NAND2X0 add_1108_U163 ( .IN1(add_1108_n154), .IN2(add_1108_n155), 
        .QN(add_1108_n147) );
  NAND2X0 add_1108_U164 ( .IN1(si_21_), .IN2(add_1108_n156), 
        .QN(add_1108_n155) );
  OR2X1 add_1108_U165 ( .IN2(n9963), .IN1(add_1108_n157), .Q(add_1108_n156) );
  NAND2X0 add_1108_U166 ( .IN1(n9963), .IN2(add_1108_n157), .QN(add_1108_n154)
         );
  INVX0 add_1108_U151 ( .ZN(add_1108_n143), .INP(n9955) );
  NAND2X0 add_1108_U152 ( .IN1(add_1108_n144), .IN2(add_1108_n145), 
        .QN(add_1108_n137) );
  NAND2X0 add_1108_U153 ( .IN1(si_22_), .IN2(add_1108_n146), 
        .QN(add_1108_n145) );
  OR2X1 add_1108_U154 ( .IN2(n9959), .IN1(add_1108_n147), .Q(add_1108_n146) );
  NAND2X0 add_1108_U155 ( .IN1(n9959), .IN2(add_1108_n147), .QN(add_1108_n144)
         );
  NOR2X0 add_1108_U156 ( .QN(N61), .IN1(add_1108_n148), .IN2(add_1108_n149) );
  AND2X1 add_1108_U157 ( .IN1(add_1108_n147), .IN2(add_1108_n150), 
        .Q(add_1108_n149) );
  NOR2X0 add_1108_U158 ( .QN(add_1108_n148), .IN1(add_1108_n147), 
        .IN2(add_1108_n150) );
  OR2X1 add_1108_U143 ( .IN2(n9955), .IN1(add_1108_n137), .Q(add_1108_n136) );
  NAND2X0 add_1108_U144 ( .IN1(n9955), .IN2(add_1108_n137), .QN(add_1108_n134)
         );
  NOR2X0 add_1108_U145 ( .QN(N62), .IN1(add_1108_n138), .IN2(add_1108_n139) );
  AND2X1 add_1108_U146 ( .IN1(add_1108_n137), .IN2(add_1108_n140), 
        .Q(add_1108_n139) );
  NOR2X0 add_1108_U147 ( .QN(add_1108_n138), .IN1(add_1108_n137), 
        .IN2(add_1108_n140) );
  NAND2X0 add_1108_U148 ( .IN1(add_1108_n141), .IN2(add_1108_n142), 
        .QN(add_1108_n140) );
  NAND2X0 add_1108_U149 ( .IN1(si_23_), .IN2(add_1108_n143), 
        .QN(add_1108_n142) );
  OR2X1 add_1108_U150 ( .IN2(si_23_), .IN1(add_1108_n143), .Q(add_1108_n141)
         );
  AND2X1 add_1108_U135 ( .IN1(add_1108_n127), .IN2(add_1108_n130), 
        .Q(add_1108_n129) );
  NOR2X0 add_1108_U136 ( .QN(add_1108_n128), .IN1(add_1108_n127), 
        .IN2(add_1108_n130) );
  NAND2X0 add_1108_U137 ( .IN1(add_1108_n131), .IN2(add_1108_n132), 
        .QN(add_1108_n130) );
  NAND2X0 add_1108_U138 ( .IN1(si_24_), .IN2(add_1108_n133), 
        .QN(add_1108_n132) );
  OR2X1 add_1108_U139 ( .IN2(si_24_), .IN1(add_1108_n133), .Q(add_1108_n131)
         );
  INVX0 add_1108_U140 ( .ZN(add_1108_n133), .INP(n9951) );
  NAND2X0 add_1108_U141 ( .IN1(add_1108_n134), .IN2(add_1108_n135), 
        .QN(add_1108_n127) );
  NAND2X0 add_1108_U142 ( .IN1(si_23_), .IN2(add_1108_n136), 
        .QN(add_1108_n135) );
  NAND2X0 add_1108_U127 ( .IN1(si_25_), .IN2(add_1108_n123), 
        .QN(add_1108_n122) );
  OR2X1 add_1108_U128 ( .IN2(si_25_), .IN1(add_1108_n123), .Q(add_1108_n121)
         );
  INVX0 add_1108_U129 ( .ZN(add_1108_n123), .INP(n9947) );
  NAND2X0 add_1108_U130 ( .IN1(add_1108_n124), .IN2(add_1108_n125), 
        .QN(add_1108_n117) );
  NAND2X0 add_1108_U131 ( .IN1(si_24_), .IN2(add_1108_n126), 
        .QN(add_1108_n125) );
  OR2X1 add_1108_U132 ( .IN2(n9951), .IN1(add_1108_n127), .Q(add_1108_n126) );
  NAND2X0 add_1108_U133 ( .IN1(n9951), .IN2(add_1108_n127), .QN(add_1108_n124)
         );
  NOR2X0 add_1108_U134 ( .QN(N63), .IN1(add_1108_n128), .IN2(add_1108_n129) );
  NAND2X0 add_1108_U119 ( .IN1(add_1108_n114), .IN2(add_1108_n115), 
        .QN(add_1108_n107) );
  NAND2X0 add_1108_U120 ( .IN1(si_25_), .IN2(add_1108_n116), 
        .QN(add_1108_n115) );
  OR2X1 add_1108_U121 ( .IN2(n9947), .IN1(add_1108_n117), .Q(add_1108_n116) );
  NAND2X0 add_1108_U122 ( .IN1(n9947), .IN2(add_1108_n117), .QN(add_1108_n114)
         );
  NOR2X0 add_1108_U123 ( .QN(N64), .IN1(add_1108_n118), .IN2(add_1108_n119) );
  AND2X1 add_1108_U124 ( .IN1(add_1108_n117), .IN2(add_1108_n120), 
        .Q(add_1108_n119) );
  NOR2X0 add_1108_U125 ( .QN(add_1108_n118), .IN1(add_1108_n117), 
        .IN2(add_1108_n120) );
  NAND2X0 add_1108_U126 ( .IN1(add_1108_n121), .IN2(add_1108_n122), 
        .QN(add_1108_n120) );
  NAND2X0 add_1108_U111 ( .IN1(n9943), .IN2(add_1108_n107), .QN(add_1108_n104)
         );
  NOR2X0 add_1108_U112 ( .QN(N65), .IN1(add_1108_n108), .IN2(add_1108_n109) );
  AND2X1 add_1108_U113 ( .IN1(add_1108_n107), .IN2(add_1108_n110), 
        .Q(add_1108_n109) );
  NOR2X0 add_1108_U114 ( .QN(add_1108_n108), .IN1(add_1108_n107), 
        .IN2(add_1108_n110) );
  NAND2X0 add_1108_U115 ( .IN1(add_1108_n111), .IN2(add_1108_n112), 
        .QN(add_1108_n110) );
  NAND2X0 add_1108_U116 ( .IN1(si_26_), .IN2(add_1108_n113), 
        .QN(add_1108_n112) );
  OR2X1 add_1108_U117 ( .IN2(si_26_), .IN1(add_1108_n113), .Q(add_1108_n111)
         );
  INVX0 add_1108_U118 ( .ZN(add_1108_n113), .INP(n9943) );
  NOR2X0 add_1108_U103 ( .QN(add_1108_n98), .IN1(add_1108_n97), 
        .IN2(add_1108_n100) );
  NAND2X0 add_1108_U104 ( .IN1(add_1108_n101), .IN2(add_1108_n102), 
        .QN(add_1108_n100) );
  NAND2X0 add_1108_U105 ( .IN1(si_27_), .IN2(add_1108_n103), 
        .QN(add_1108_n102) );
  OR2X1 add_1108_U106 ( .IN2(si_27_), .IN1(add_1108_n103), .Q(add_1108_n101)
         );
  INVX0 add_1108_U107 ( .ZN(add_1108_n103), .INP(n9939) );
  NAND2X0 add_1108_U108 ( .IN1(add_1108_n104), .IN2(add_1108_n105), 
        .QN(add_1108_n97) );
  NAND2X0 add_1108_U109 ( .IN1(si_26_), .IN2(add_1108_n106), 
        .QN(add_1108_n105) );
  OR2X1 add_1108_U110 ( .IN2(n9943), .IN1(add_1108_n107), .Q(add_1108_n106) );
  OR2X1 add_1108_U95 ( .IN2(si_28_), .IN1(add_1108_n93), .Q(add_1108_n91) );
  INVX0 add_1108_U96 ( .ZN(add_1108_n93), .INP(n9935) );
  NAND2X0 add_1108_U97 ( .IN1(add_1108_n94), .IN2(add_1108_n95), 
        .QN(add_1108_n87) );
  NAND2X0 add_1108_U98 ( .IN1(si_27_), .IN2(add_1108_n96), .QN(add_1108_n95)
         );
  OR2X1 add_1108_U99 ( .IN2(n9939), .IN1(add_1108_n97), .Q(add_1108_n96) );
  NAND2X0 add_1108_U100 ( .IN1(n9939), .IN2(add_1108_n97), .QN(add_1108_n94)
         );
  NOR2X0 add_1108_U101 ( .QN(N66), .IN1(add_1108_n98), .IN2(add_1108_n99) );
  AND2X1 add_1108_U102 ( .IN1(add_1108_n97), .IN2(add_1108_n100), 
        .Q(add_1108_n99) );
  NAND2X0 add_1108_U87 ( .IN1(si_28_), .IN2(add_1108_n86), .QN(add_1108_n85)
         );
  OR2X1 add_1108_U88 ( .IN2(n9935), .IN1(add_1108_n87), .Q(add_1108_n86) );
  NAND2X0 add_1108_U89 ( .IN1(n9935), .IN2(add_1108_n87), .QN(add_1108_n84) );
  NOR2X0 add_1108_U90 ( .QN(N67), .IN1(add_1108_n88), .IN2(add_1108_n89) );
  AND2X1 add_1108_U91 ( .IN1(add_1108_n87), .IN2(add_1108_n90), 
        .Q(add_1108_n89) );
  NOR2X0 add_1108_U92 ( .QN(add_1108_n88), .IN1(add_1108_n87), 
        .IN2(add_1108_n90) );
  NAND2X0 add_1108_U93 ( .IN1(add_1108_n91), .IN2(add_1108_n92), 
        .QN(add_1108_n90) );
  NAND2X0 add_1108_U94 ( .IN1(si_28_), .IN2(add_1108_n93), .QN(add_1108_n92)
         );
  NOR2X0 add_1108_U79 ( .QN(N68), .IN1(add_1108_n78), .IN2(add_1108_n79) );
  AND2X1 add_1108_U80 ( .IN1(add_1108_n70), .IN2(add_1108_n80), 
        .Q(add_1108_n79) );
  NOR2X0 add_1108_U81 ( .QN(add_1108_n78), .IN1(add_1108_n70), 
        .IN2(add_1108_n80) );
  NAND2X0 add_1108_U82 ( .IN1(add_1108_n81), .IN2(add_1108_n82), 
        .QN(add_1108_n80) );
  NAND2X0 add_1108_U83 ( .IN1(si_29_), .IN2(add_1108_n83), .QN(add_1108_n82)
         );
  OR2X1 add_1108_U84 ( .IN2(si_29_), .IN1(add_1108_n83), .Q(add_1108_n81) );
  INVX0 add_1108_U85 ( .ZN(add_1108_n83), .INP(n10095) );
  NAND2X0 add_1108_U86 ( .IN1(add_1108_n84), .IN2(add_1108_n85), 
        .QN(add_1108_n70) );
  NAND2X0 add_1108_U71 ( .IN1(n10095), .IN2(add_1108_n70), .QN(add_1108_n67)
         );
  NOR2X0 add_1108_U72 ( .QN(N41), .IN1(add_1108_n71), .IN2(add_1108_n72) );
  AND2X1 add_1108_U73 ( .IN1(add_1108_n73), .IN2(add_1108_n74), 
        .Q(add_1108_n72) );
  NOR2X0 add_1108_U74 ( .QN(add_1108_n71), .IN1(add_1108_n73), 
        .IN2(add_1108_n74) );
  NAND2X0 add_1108_U75 ( .IN1(add_1108_n75), .IN2(add_1108_n76), 
        .QN(add_1108_n74) );
  NAND2X0 add_1108_U76 ( .IN1(si_2_), .IN2(add_1108_n77), .QN(add_1108_n76) );
  OR2X1 add_1108_U77 ( .IN2(si_2_), .IN1(add_1108_n77), .Q(add_1108_n75) );
  INVX0 add_1108_U78 ( .ZN(add_1108_n77), .INP(n9899) );
  NOR2X0 add_1108_U63 ( .QN(add_1108_n61), .IN1(add_1108_n57), 
        .IN2(add_1108_n63) );
  NAND2X0 add_1108_U64 ( .IN1(add_1108_n64), .IN2(add_1108_n65), 
        .QN(add_1108_n63) );
  NAND2X0 add_1108_U65 ( .IN1(si_30_), .IN2(add_1108_n66), .QN(add_1108_n65)
         );
  OR2X1 add_1108_U66 ( .IN2(si_30_), .IN1(add_1108_n66), .Q(add_1108_n64) );
  INVX0 add_1108_U67 ( .ZN(add_1108_n66), .INP(n10103) );
  NAND2X0 add_1108_U68 ( .IN1(add_1108_n67), .IN2(add_1108_n68), 
        .QN(add_1108_n57) );
  NAND2X0 add_1108_U69 ( .IN1(si_29_), .IN2(add_1108_n69), .QN(add_1108_n68)
         );
  OR2X1 add_1108_U70 ( .IN2(n10095), .IN1(add_1108_n70), .Q(add_1108_n69) );
  OR2X1 add_1108_U55 ( .IN2(n10103), .IN1(add_1108_n57), .Q(add_1108_n56) );
  NAND2X0 add_1108_U56 ( .IN1(n10103), .IN2(add_1108_n57), .QN(add_1108_n54)
         );
  NAND2X0 add_1108_U57 ( .IN1(add_1108_n58), .IN2(add_1108_n59), 
        .QN(add_1108_n53) );
  NAND2X0 add_1108_U58 ( .IN1(si_31_), .IN2(add_1108_n60), .QN(add_1108_n59)
         );
  OR2X1 add_1108_U59 ( .IN2(si_31_), .IN1(add_1108_n60), .Q(add_1108_n58) );
  INVX0 add_1108_U60 ( .ZN(add_1108_n60), .INP(n9345) );
  NOR2X0 add_1108_U61 ( .QN(N69), .IN1(add_1108_n61), .IN2(add_1108_n62) );
  AND2X1 add_1108_U62 ( .IN1(add_1108_n57), .IN2(add_1108_n63), 
        .Q(add_1108_n62) );
  NAND2X0 add_1108_U47 ( .IN1(si_3_), .IN2(add_1108_n49), .QN(add_1108_n48) );
  OR2X1 add_1108_U48 ( .IN2(si_3_), .IN1(add_1108_n49), .Q(add_1108_n47) );
  INVX0 add_1108_U49 ( .ZN(add_1108_n49), .INP(n9895) );
  NOR2X0 add_1108_U50 ( .QN(N70), .IN1(add_1108_n50), .IN2(add_1108_n51) );
  AND2X1 add_1108_U51 ( .IN1(add_1108_n52), .IN2(add_1108_n53), 
        .Q(add_1108_n51) );
  NOR2X0 add_1108_U52 ( .QN(add_1108_n50), .IN1(add_1108_n53), 
        .IN2(add_1108_n52) );
  NAND2X0 add_1108_U53 ( .IN1(add_1108_n54), .IN2(add_1108_n55), 
        .QN(add_1108_n52) );
  NAND2X0 add_1108_U54 ( .IN1(si_30_), .IN2(add_1108_n56), .QN(add_1108_n55)
         );
  NAND2X0 add_1108_U39 ( .IN1(add_1108_n40), .IN2(add_1108_n41), 
        .QN(add_1108_n39) );
  NAND2X0 add_1108_U40 ( .IN1(si_4_), .IN2(add_1108_n42), .QN(add_1108_n41) );
  OR2X1 add_1108_U41 ( .IN2(si_4_), .IN1(add_1108_n42), .Q(add_1108_n40) );
  INVX0 add_1108_U42 ( .ZN(add_1108_n42), .INP(n9891) );
  NOR2X0 add_1108_U43 ( .QN(N42), .IN1(add_1108_n43), .IN2(add_1108_n44) );
  AND2X1 add_1108_U44 ( .IN1(add_1108_n45), .IN2(add_1108_n46), 
        .Q(add_1108_n44) );
  NOR2X0 add_1108_U45 ( .QN(add_1108_n43), .IN1(add_1108_n45), 
        .IN2(add_1108_n46) );
  NAND2X0 add_1108_U46 ( .IN1(add_1108_n47), .IN2(add_1108_n48), 
        .QN(add_1108_n46) );
  NOR2X0 add_1108_U31 ( .QN(add_1108_n29), .IN1(add_1108_n31), 
        .IN2(add_1108_n32) );
  NAND2X0 add_1108_U32 ( .IN1(add_1108_n33), .IN2(add_1108_n34), 
        .QN(add_1108_n32) );
  NAND2X0 add_1108_U33 ( .IN1(si_5_), .IN2(add_1108_n35), .QN(add_1108_n34) );
  OR2X1 add_1108_U34 ( .IN2(si_5_), .IN1(add_1108_n35), .Q(add_1108_n33) );
  INVX0 add_1108_U35 ( .ZN(add_1108_n35), .INP(n9887) );
  NOR2X0 add_1108_U36 ( .QN(N43), .IN1(add_1108_n36), .IN2(add_1108_n37) );
  AND2X1 add_1108_U37 ( .IN1(add_1108_n38), .IN2(add_1108_n39), 
        .Q(add_1108_n37) );
  NOR2X0 add_1108_U38 ( .QN(add_1108_n36), .IN1(add_1108_n38), 
        .IN2(add_1108_n39) );
  AND2X1 add_1108_U23 ( .IN1(add_1108_n24), .IN2(add_1108_n25), 
        .Q(add_1108_n23) );
  NOR2X0 add_1108_U24 ( .QN(add_1108_n22), .IN1(add_1108_n24), 
        .IN2(add_1108_n25) );
  NAND2X0 add_1108_U25 ( .IN1(add_1108_n26), .IN2(add_1108_n27), 
        .QN(add_1108_n25) );
  NAND2X0 add_1108_U26 ( .IN1(si_6_), .IN2(add_1108_n28), .QN(add_1108_n27) );
  OR2X1 add_1108_U27 ( .IN2(si_6_), .IN1(add_1108_n28), .Q(add_1108_n26) );
  INVX0 add_1108_U28 ( .ZN(add_1108_n28), .INP(n9883) );
  NOR2X0 add_1108_U29 ( .QN(N44), .IN1(add_1108_n29), .IN2(add_1108_n30) );
  AND2X1 add_1108_U30 ( .IN1(add_1108_n31), .IN2(add_1108_n32), 
        .Q(add_1108_n30) );
  NOR2X0 add_1108_U15 ( .QN(N46), .IN1(add_1108_n15), .IN2(add_1108_n16) );
  AND2X1 add_1108_U16 ( .IN1(add_1108_n17), .IN2(add_1108_n18), 
        .Q(add_1108_n16) );
  NOR2X0 add_1108_U17 ( .QN(add_1108_n15), .IN1(add_1108_n17), 
        .IN2(add_1108_n18) );
  NAND2X0 add_1108_U18 ( .IN1(add_1108_n19), .IN2(add_1108_n20), 
        .QN(add_1108_n18) );
  NAND2X0 add_1108_U19 ( .IN1(si_7_), .IN2(add_1108_n21), .QN(add_1108_n20) );
  OR2X1 add_1108_U20 ( .IN2(si_7_), .IN1(add_1108_n21), .Q(add_1108_n19) );
  INVX0 add_1108_U21 ( .ZN(add_1108_n21), .INP(n9879) );
  NOR2X0 add_1108_U22 ( .QN(N45), .IN1(add_1108_n22), .IN2(add_1108_n23) );
  INVX0 add_1108_U7 ( .ZN(add_1108_n7), .INP(n9871) );
  NOR2X0 add_1108_U8 ( .QN(N47), .IN1(add_1108_n8), .IN2(add_1108_n9) );
  AND2X1 add_1108_U9 ( .IN1(add_1108_n10), .IN2(add_1108_n11), .Q(add_1108_n9)
         );
  NOR2X0 add_1108_U10 ( .QN(add_1108_n8), .IN1(add_1108_n10), 
        .IN2(add_1108_n11) );
  NAND2X0 add_1108_U11 ( .IN1(add_1108_n12), .IN2(add_1108_n13), 
        .QN(add_1108_n11) );
  NAND2X0 add_1108_U12 ( .IN1(si_8_), .IN2(add_1108_n14), .QN(add_1108_n13) );
  OR2X1 add_1108_U13 ( .IN2(si_8_), .IN1(add_1108_n14), .Q(add_1108_n12) );
  INVX0 add_1108_U14 ( .ZN(add_1108_n14), .INP(n9875) );
  NOR2X0 add_1108_U1 ( .QN(N48), .IN1(add_1108_n1), .IN2(add_1108_n2) );
  AND2X1 add_1108_U2 ( .IN1(add_1108_n3), .IN2(add_1108_n4), .Q(add_1108_n2)
         );
  NOR2X0 add_1108_U3 ( .QN(add_1108_n1), .IN1(add_1108_n3), .IN2(add_1108_n4)
         );
  NAND2X0 add_1108_U4 ( .IN1(add_1108_n5), .IN2(add_1108_n6), .QN(add_1108_n4)
         );
  NAND2X0 add_1108_U5 ( .IN1(si_9_), .IN2(add_1108_n7), .QN(add_1108_n6) );
  OR2X1 add_1108_U6 ( .IN2(si_9_), .IN1(add_1108_n7), .Q(add_1108_n5) );
  NAND2X0 r839_U89 ( .IN1(r839_n97), .IN2(r839_n98), .QN(r839_n91) );
  NAND2X0 r839_U88 ( .IN1(P2_N5096), .IN2(r839_n96), .QN(r839_n92) );
  OR2X1 r839_U87 ( .IN2(P2_N5096), .IN1(r839_n96), .Q(r839_n94) );
  NAND2X0 r839_U86 ( .IN1(r839_n94), .IN2(r839_n95), .QN(r839_n93) );
  NAND2X0 r839_U85 ( .IN1(r839_n92), .IN2(r839_n93), .QN(r839_n86) );
  NAND2X0 r839_U84 ( .IN1(r839_n91), .IN2(r839_n86), .QN(r839_n89) );
  OR2X1 r839_U83 ( .IN2(r839_n86), .IN1(r839_n91), .Q(r839_n90) );
  NAND2X0 r839_U82 ( .IN1(r839_n89), .IN2(r839_n90), .QN(P2_N1664) );
  INVX0 r839_U81 ( .ZN(r839_n75), .INP(P2_N1513) );
  NAND2X0 r839_U80 ( .IN1(n7227), .IN2(r839_n75), .QN(r839_n87) );
  OR2X1 r839_U79 ( .IN2(n7227), .IN1(r839_n75), .Q(r839_n88) );
  NAND2X0 r839_U78 ( .IN1(r839_n87), .IN2(r839_n88), .QN(r839_n81) );
  NAND2X0 r839_U77 ( .IN1(P2_N5097), .IN2(r839_n86), .QN(r839_n82) );
  OR2X1 r839_U76 ( .IN2(P2_N5097), .IN1(r839_n86), .Q(r839_n84) );
  NAND2X0 r839_U75 ( .IN1(r839_n84), .IN2(r839_n85), .QN(r839_n83) );
  NAND2X0 r839_U74 ( .IN1(r839_n82), .IN2(r839_n83), .QN(r839_n76) );
  NAND2X0 r839_U73 ( .IN1(r839_n81), .IN2(r839_n76), .QN(r839_n79) );
  OR2X1 r839_U72 ( .IN2(r839_n76), .IN1(r839_n81), .Q(r839_n80) );
  NAND2X0 r839_U71 ( .IN1(r839_n79), .IN2(r839_n80), .QN(P2_N1665) );
  INVX0 r839_U70 ( .ZN(r839_n64), .INP(P2_N1514) );
  NAND2X0 r839_U69 ( .IN1(P2_N5099), .IN2(r839_n64), .QN(r839_n77) );
  OR2X1 r839_U68 ( .IN2(P2_N5099), .IN1(r839_n64), .Q(r839_n78) );
  NAND2X0 r839_U67 ( .IN1(r839_n77), .IN2(r839_n78), .QN(r839_n71) );
  NAND2X0 r839_U66 ( .IN1(n7227), .IN2(r839_n76), .QN(r839_n72) );
  OR2X1 r839_U65 ( .IN2(n7227), .IN1(r839_n76), .Q(r839_n74) );
  NAND2X0 r839_U64 ( .IN1(r839_n74), .IN2(r839_n75), .QN(r839_n73) );
  NAND2X0 r839_U63 ( .IN1(r839_n72), .IN2(r839_n73), .QN(r839_n65) );
  NAND2X0 r839_U62 ( .IN1(r839_n71), .IN2(r839_n65), .QN(r839_n69) );
  OR2X1 r839_U61 ( .IN2(r839_n65), .IN1(r839_n71), .Q(r839_n70) );
  NAND2X0 r839_U60 ( .IN1(r839_n69), .IN2(r839_n70), .QN(P2_N1666) );
  OR2X1 r839_U58 ( .IN2(P2_N1515), .IN1(n7266), .Q(r839_n66) );
  NAND2X0 r839_U57 ( .IN1(P2_N1515), .IN2(n7266), .QN(r839_n67) );
  NAND2X0 r839_U56 ( .IN1(r839_n66), .IN2(r839_n67), .QN(r839_n60) );
  NAND2X0 r839_U55 ( .IN1(P2_N5099), .IN2(r839_n65), .QN(r839_n61) );
  OR2X1 r839_U54 ( .IN2(P2_N5099), .IN1(r839_n65), .Q(r839_n63) );
  NAND2X0 r839_U53 ( .IN1(r839_n63), .IN2(r839_n64), .QN(r839_n62) );
  NAND2X0 r839_U52 ( .IN1(r839_n61), .IN2(r839_n62), .QN(r839_n59) );
  NAND2X0 r839_U51 ( .IN1(r839_n60), .IN2(r839_n59), .QN(r839_n57) );
  OR2X1 r839_U50 ( .IN2(r839_n60), .IN1(r839_n59), .Q(r839_n58) );
  NAND2X0 r839_U49 ( .IN1(r839_n57), .IN2(r839_n58), .QN(P2_N1667) );
  NAND2X0 r839_U48 ( .IN1(P2_N5073), .IN2(r839_n56), .QN(r839_n54) );
  OR2X1 r839_U47 ( .IN2(P2_N5073), .IN1(r839_n56), .Q(r839_n55) );
  NAND2X0 r839_U46 ( .IN1(r839_n54), .IN2(r839_n55), .QN(r839_n52) );
  NAND2X0 r839_U45 ( .IN1(r839_n52), .IN2(r839_n53), .QN(r839_n50) );
  OR2X1 r839_U44 ( .IN2(r839_n53), .IN1(r839_n52), .Q(r839_n51) );
  NAND2X0 r839_U43 ( .IN1(r839_n50), .IN2(r839_n51), .QN(P2_N1640) );
  NAND2X0 r839_U42 ( .IN1(P2_N5074), .IN2(r839_n49), .QN(r839_n47) );
  OR2X1 r839_U41 ( .IN2(P2_N5074), .IN1(r839_n49), .Q(r839_n48) );
  NAND2X0 r839_U40 ( .IN1(r839_n47), .IN2(r839_n48), .QN(r839_n45) );
  NAND2X0 r839_U39 ( .IN1(r839_n45), .IN2(r839_n46), .QN(r839_n43) );
  OR2X1 r839_U38 ( .IN2(r839_n46), .IN1(r839_n45), .Q(r839_n44) );
  NAND2X0 r839_U37 ( .IN1(r839_n43), .IN2(r839_n44), .QN(P2_N1641) );
  NAND2X0 r839_U36 ( .IN1(P2_N5075), .IN2(r839_n42), .QN(r839_n40) );
  OR2X1 r839_U35 ( .IN2(P2_N5075), .IN1(r839_n42), .Q(r839_n41) );
  NAND2X0 r839_U34 ( .IN1(r839_n40), .IN2(r839_n41), .QN(r839_n38) );
  NAND2X0 r839_U33 ( .IN1(r839_n38), .IN2(r839_n39), .QN(r839_n36) );
  OR2X1 r839_U32 ( .IN2(r839_n39), .IN1(r839_n38), .Q(r839_n37) );
  NAND2X0 r839_U31 ( .IN1(r839_n36), .IN2(r839_n37), .QN(P2_N1642) );
  NAND2X0 r839_U30 ( .IN1(P2_N5076), .IN2(r839_n35), .QN(r839_n33) );
  OR2X1 r839_U29 ( .IN2(P2_N5076), .IN1(r839_n35), .Q(r839_n34) );
  NAND2X0 r839_U28 ( .IN1(r839_n33), .IN2(r839_n34), .QN(r839_n31) );
  NAND2X0 r839_U27 ( .IN1(r839_n31), .IN2(r839_n32), .QN(r839_n29) );
  OR2X1 r839_U26 ( .IN2(r839_n32), .IN1(r839_n31), .Q(r839_n30) );
  NAND2X0 r839_U25 ( .IN1(r839_n29), .IN2(r839_n30), .QN(P2_N1643) );
  NAND2X0 r839_U24 ( .IN1(n7162), .IN2(r839_n28), .QN(r839_n26) );
  OR2X1 r839_U23 ( .IN2(n7162), .IN1(r839_n28), .Q(r839_n27) );
  NAND2X0 r839_U22 ( .IN1(r839_n26), .IN2(r839_n27), .QN(r839_n24) );
  NAND2X0 r839_U21 ( .IN1(r839_n24), .IN2(r839_n25), .QN(r839_n22) );
  OR2X1 r839_U20 ( .IN2(r839_n25), .IN1(r839_n24), .Q(r839_n23) );
  NAND2X0 r839_U19 ( .IN1(r839_n22), .IN2(r839_n23), .QN(P2_N1644) );
  NAND2X0 r839_U18 ( .IN1(n7158), .IN2(r839_n21), .QN(r839_n19) );
  OR2X1 r839_U17 ( .IN2(n7158), .IN1(r839_n21), .Q(r839_n20) );
  NAND2X0 r839_U16 ( .IN1(r839_n19), .IN2(r839_n20), .QN(r839_n17) );
  NAND2X0 r839_U15 ( .IN1(r839_n17), .IN2(r839_n18), .QN(r839_n15) );
  OR2X1 r839_U14 ( .IN2(r839_n18), .IN1(r839_n17), .Q(r839_n16) );
  NAND2X0 r839_U13 ( .IN1(r839_n15), .IN2(r839_n16), .QN(P2_N1645) );
  NAND2X0 r839_U12 ( .IN1(P2_N5079), .IN2(r839_n14), .QN(r839_n12) );
  OR2X1 r839_U11 ( .IN2(P2_N5079), .IN1(r839_n14), .Q(r839_n13) );
  NAND2X0 r839_U10 ( .IN1(r839_n12), .IN2(r839_n13), .QN(r839_n10) );
  NAND2X0 r839_U9 ( .IN1(r839_n10), .IN2(r839_n11), .QN(r839_n8) );
  OR2X1 r839_U8 ( .IN2(r839_n11), .IN1(r839_n10), .Q(r839_n9) );
  NAND2X0 r839_U7 ( .IN1(r839_n8), .IN2(r839_n9), .QN(P2_N1646) );
  NAND2X0 r839_U6 ( .IN1(n7151), .IN2(r839_n7), .QN(r839_n5) );
  OR2X1 r839_U5 ( .IN2(n7151), .IN1(r839_n7), .Q(r839_n6) );
  NAND2X0 r839_U4 ( .IN1(r839_n5), .IN2(r839_n6), .QN(r839_n3) );
  NAND2X0 r839_U3 ( .IN1(r839_n3), .IN2(r839_n4), .QN(r839_n1) );
  OR2X1 r839_U2 ( .IN2(r839_n4), .IN1(r839_n3), .Q(r839_n2) );
  NAND2X0 r839_U1 ( .IN1(r839_n1), .IN2(r839_n2), .QN(P2_N1647) );
  NAND2X0 r839_U182 ( .IN1(n7194), .IN2(r839_n184), .QN(r839_n180) );
  OR2X1 r839_U181 ( .IN2(n7194), .IN1(r839_n184), .Q(r839_n182) );
  NAND2X0 r839_U180 ( .IN1(r839_n182), .IN2(r839_n183), .QN(r839_n181) );
  NAND2X0 r839_U179 ( .IN1(r839_n180), .IN2(r839_n181), .QN(r839_n174) );
  NAND2X0 r839_U178 ( .IN1(r839_n179), .IN2(r839_n174), .QN(r839_n177) );
  OR2X1 r839_U177 ( .IN2(r839_n174), .IN1(r839_n179), .Q(r839_n178) );
  NAND2X0 r839_U176 ( .IN1(r839_n177), .IN2(r839_n178), .QN(P2_N1656) );
  INVX0 r839_U175 ( .ZN(r839_n155), .INP(P2_N1505) );
  NAND2X0 r839_U174 ( .IN1(P2_N5090), .IN2(r839_n155), .QN(r839_n175) );
  OR2X1 r839_U173 ( .IN2(P2_N5090), .IN1(r839_n155), .Q(r839_n176) );
  NAND2X0 r839_U172 ( .IN1(r839_n175), .IN2(r839_n176), .QN(r839_n169) );
  NAND2X0 r839_U171 ( .IN1(n7187), .IN2(r839_n174), .QN(r839_n170) );
  OR2X1 r839_U170 ( .IN2(n7187), .IN1(r839_n174), .Q(r839_n172) );
  NAND2X0 r839_U169 ( .IN1(r839_n172), .IN2(r839_n173), .QN(r839_n171) );
  NAND2X0 r839_U168 ( .IN1(r839_n170), .IN2(r839_n171), .QN(r839_n156) );
  NAND2X0 r839_U167 ( .IN1(r839_n169), .IN2(r839_n156), .QN(r839_n167) );
  OR2X1 r839_U166 ( .IN2(r839_n156), .IN1(r839_n169), .Q(r839_n168) );
  NAND2X0 r839_U165 ( .IN1(r839_n167), .IN2(r839_n168), .QN(P2_N1657) );
  NAND2X0 r839_U164 ( .IN1(P2_N5072), .IN2(r839_n166), .QN(r839_n163) );
  NAND2X0 r839_U163 ( .IN1(P2_N1487), .IN2(n7184), .QN(r839_n164) );
  NAND2X0 r839_U162 ( .IN1(r839_n163), .IN2(r839_n164), .QN(r839_n161) );
  NAND2X0 r839_U161 ( .IN1(r839_n161), .IN2(r839_n162), .QN(r839_n159) );
  OR2X1 r839_U160 ( .IN2(r839_n162), .IN1(r839_n161), .Q(r839_n160) );
  NAND2X0 r839_U159 ( .IN1(r839_n159), .IN2(r839_n160), .QN(P2_N1639) );
  INVX0 r839_U158 ( .ZN(r839_n145), .INP(P2_N1506) );
  NAND2X0 r839_U157 ( .IN1(P2_N5091), .IN2(r839_n145), .QN(r839_n157) );
  OR2X1 r839_U156 ( .IN2(P2_N5091), .IN1(r839_n145), .Q(r839_n158) );
  NAND2X0 r839_U155 ( .IN1(r839_n157), .IN2(r839_n158), .QN(r839_n151) );
  NAND2X0 r839_U154 ( .IN1(P2_N5090), .IN2(r839_n156), .QN(r839_n152) );
  OR2X1 r839_U153 ( .IN2(P2_N5090), .IN1(r839_n156), .Q(r839_n154) );
  NAND2X0 r839_U152 ( .IN1(r839_n154), .IN2(r839_n155), .QN(r839_n153) );
  NAND2X0 r839_U151 ( .IN1(r839_n152), .IN2(r839_n153), .QN(r839_n146) );
  NAND2X0 r839_U150 ( .IN1(r839_n151), .IN2(r839_n146), .QN(r839_n149) );
  OR2X1 r839_U149 ( .IN2(r839_n146), .IN1(r839_n151), .Q(r839_n150) );
  NAND2X0 r839_U148 ( .IN1(r839_n149), .IN2(r839_n150), .QN(P2_N1658) );
  INVX0 r839_U147 ( .ZN(r839_n135), .INP(P2_N1507) );
  NAND2X0 r839_U146 ( .IN1(n7252), .IN2(r839_n135), .QN(r839_n147) );
  OR2X1 r839_U145 ( .IN2(n7252), .IN1(r839_n135), .Q(r839_n148) );
  NAND2X0 r839_U144 ( .IN1(r839_n147), .IN2(r839_n148), .QN(r839_n141) );
  NAND2X0 r839_U143 ( .IN1(P2_N5091), .IN2(r839_n146), .QN(r839_n142) );
  OR2X1 r839_U142 ( .IN2(P2_N5091), .IN1(r839_n146), .Q(r839_n144) );
  NAND2X0 r839_U141 ( .IN1(r839_n144), .IN2(r839_n145), .QN(r839_n143) );
  NAND2X0 r839_U140 ( .IN1(r839_n142), .IN2(r839_n143), .QN(r839_n136) );
  NAND2X0 r839_U139 ( .IN1(r839_n141), .IN2(r839_n136), .QN(r839_n139) );
  OR2X1 r839_U138 ( .IN2(r839_n136), .IN1(r839_n141), .Q(r839_n140) );
  NAND2X0 r839_U137 ( .IN1(r839_n139), .IN2(r839_n140), .QN(P2_N1659) );
  INVX0 r839_U136 ( .ZN(r839_n125), .INP(P2_N1508) );
  NAND2X0 r839_U135 ( .IN1(n7247), .IN2(r839_n125), .QN(r839_n137) );
  OR2X1 r839_U134 ( .IN2(n7247), .IN1(r839_n125), .Q(r839_n138) );
  NAND2X0 r839_U133 ( .IN1(r839_n137), .IN2(r839_n138), .QN(r839_n131) );
  NAND2X0 r839_U132 ( .IN1(n7252), .IN2(r839_n136), .QN(r839_n132) );
  OR2X1 r839_U131 ( .IN2(n7252), .IN1(r839_n136), .Q(r839_n134) );
  NAND2X0 r839_U130 ( .IN1(r839_n134), .IN2(r839_n135), .QN(r839_n133) );
  NAND2X0 r839_U129 ( .IN1(r839_n132), .IN2(r839_n133), .QN(r839_n126) );
  NAND2X0 r839_U128 ( .IN1(r839_n131), .IN2(r839_n126), .QN(r839_n129) );
  OR2X1 r839_U127 ( .IN2(r839_n126), .IN1(r839_n131), .Q(r839_n130) );
  NAND2X0 r839_U126 ( .IN1(r839_n129), .IN2(r839_n130), .QN(P2_N1660) );
  INVX0 r839_U125 ( .ZN(r839_n115), .INP(P2_N1509) );
  NAND2X0 r839_U124 ( .IN1(n7242), .IN2(r839_n115), .QN(r839_n127) );
  OR2X1 r839_U123 ( .IN2(n7242), .IN1(r839_n115), .Q(r839_n128) );
  NAND2X0 r839_U122 ( .IN1(r839_n127), .IN2(r839_n128), .QN(r839_n121) );
  NAND2X0 r839_U121 ( .IN1(n7247), .IN2(r839_n126), .QN(r839_n122) );
  OR2X1 r839_U120 ( .IN2(n7247), .IN1(r839_n126), .Q(r839_n124) );
  NAND2X0 r839_U119 ( .IN1(r839_n124), .IN2(r839_n125), .QN(r839_n123) );
  NAND2X0 r839_U118 ( .IN1(r839_n122), .IN2(r839_n123), .QN(r839_n116) );
  NAND2X0 r839_U117 ( .IN1(r839_n121), .IN2(r839_n116), .QN(r839_n119) );
  OR2X1 r839_U116 ( .IN2(r839_n116), .IN1(r839_n121), .Q(r839_n120) );
  NAND2X0 r839_U115 ( .IN1(r839_n119), .IN2(r839_n120), .QN(P2_N1661) );
  INVX0 r839_U114 ( .ZN(r839_n105), .INP(P2_N1510) );
  NAND2X0 r839_U113 ( .IN1(n7238), .IN2(r839_n105), .QN(r839_n117) );
  OR2X1 r839_U112 ( .IN2(n7238), .IN1(r839_n105), .Q(r839_n118) );
  NAND2X0 r839_U111 ( .IN1(r839_n117), .IN2(r839_n118), .QN(r839_n111) );
  NAND2X0 r839_U110 ( .IN1(n7242), .IN2(r839_n116), .QN(r839_n112) );
  OR2X1 r839_U109 ( .IN2(n7242), .IN1(r839_n116), .Q(r839_n114) );
  NAND2X0 r839_U108 ( .IN1(r839_n114), .IN2(r839_n115), .QN(r839_n113) );
  NAND2X0 r839_U107 ( .IN1(r839_n112), .IN2(r839_n113), .QN(r839_n106) );
  NAND2X0 r839_U106 ( .IN1(r839_n111), .IN2(r839_n106), .QN(r839_n109) );
  OR2X1 r839_U105 ( .IN2(r839_n106), .IN1(r839_n111), .Q(r839_n110) );
  NAND2X0 r839_U104 ( .IN1(r839_n109), .IN2(r839_n110), .QN(P2_N1662) );
  INVX0 r839_U103 ( .ZN(r839_n95), .INP(P2_N1511) );
  NAND2X0 r839_U102 ( .IN1(P2_N5096), .IN2(r839_n95), .QN(r839_n107) );
  OR2X1 r839_U101 ( .IN2(P2_N5096), .IN1(r839_n95), .Q(r839_n108) );
  NAND2X0 r839_U100 ( .IN1(r839_n107), .IN2(r839_n108), .QN(r839_n101) );
  NAND2X0 r839_U99 ( .IN1(n7238), .IN2(r839_n106), .QN(r839_n102) );
  OR2X1 r839_U98 ( .IN2(n7238), .IN1(r839_n106), .Q(r839_n104) );
  NAND2X0 r839_U97 ( .IN1(r839_n104), .IN2(r839_n105), .QN(r839_n103) );
  NAND2X0 r839_U96 ( .IN1(r839_n102), .IN2(r839_n103), .QN(r839_n96) );
  NAND2X0 r839_U95 ( .IN1(r839_n101), .IN2(r839_n96), .QN(r839_n99) );
  OR2X1 r839_U94 ( .IN2(r839_n96), .IN1(r839_n101), .Q(r839_n100) );
  NAND2X0 r839_U93 ( .IN1(r839_n99), .IN2(r839_n100), .QN(P2_N1663) );
  INVX0 r839_U92 ( .ZN(r839_n85), .INP(P2_N1512) );
  NAND2X0 r839_U91 ( .IN1(P2_N5097), .IN2(r839_n85), .QN(r839_n97) );
  OR2X1 r839_U90 ( .IN2(P2_N5097), .IN1(r839_n85), .Q(r839_n98) );
  OR2X1 r839_U275 ( .IN2(P2_N5079), .IN1(r839_n11), .Q(r839_n265) );
  INVX0 r839_U274 ( .ZN(r839_n14), .INP(P2_N1494) );
  NAND2X0 r839_U273 ( .IN1(r839_n265), .IN2(r839_n14), .QN(r839_n264) );
  NAND2X0 r839_U272 ( .IN1(r839_n263), .IN2(r839_n264), .QN(r839_n4) );
  NAND2X0 r839_U271 ( .IN1(n7151), .IN2(r839_n4), .QN(r839_n260) );
  OR2X1 r839_U270 ( .IN2(n7151), .IN1(r839_n4), .Q(r839_n262) );
  INVX0 r839_U269 ( .ZN(r839_n7), .INP(P2_N1495) );
  NAND2X0 r839_U268 ( .IN1(r839_n262), .IN2(r839_n7), .QN(r839_n261) );
  NAND2X0 r839_U267 ( .IN1(r839_n260), .IN2(r839_n261), .QN(r839_n254) );
  NAND2X0 r839_U266 ( .IN1(r839_n259), .IN2(r839_n254), .QN(r839_n257) );
  OR2X1 r839_U265 ( .IN2(r839_n254), .IN1(r839_n259), .Q(r839_n258) );
  NAND2X0 r839_U264 ( .IN1(r839_n257), .IN2(r839_n258), .QN(P2_N1648) );
  INVX0 r839_U263 ( .ZN(r839_n243), .INP(P2_N1497) );
  NAND2X0 r839_U262 ( .IN1(P2_N5082), .IN2(r839_n243), .QN(r839_n255) );
  OR2X1 r839_U261 ( .IN2(P2_N5082), .IN1(r839_n243), .Q(r839_n256) );
  NAND2X0 r839_U260 ( .IN1(r839_n255), .IN2(r839_n256), .QN(r839_n249) );
  NAND2X0 r839_U259 ( .IN1(P2_N5081), .IN2(r839_n254), .QN(r839_n250) );
  OR2X1 r839_U258 ( .IN2(P2_N5081), .IN1(r839_n254), .Q(r839_n252) );
  NAND2X0 r839_U257 ( .IN1(r839_n252), .IN2(r839_n253), .QN(r839_n251) );
  NAND2X0 r839_U256 ( .IN1(r839_n250), .IN2(r839_n251), .QN(r839_n244) );
  NAND2X0 r839_U255 ( .IN1(r839_n249), .IN2(r839_n244), .QN(r839_n247) );
  OR2X1 r839_U254 ( .IN2(r839_n244), .IN1(r839_n249), .Q(r839_n248) );
  NAND2X0 r839_U253 ( .IN1(r839_n247), .IN2(r839_n248), .QN(P2_N1649) );
  INVX0 r839_U252 ( .ZN(r839_n233), .INP(P2_N1498) );
  NAND2X0 r839_U251 ( .IN1(n7210), .IN2(r839_n233), .QN(r839_n245) );
  OR2X1 r839_U250 ( .IN2(n7210), .IN1(r839_n233), .Q(r839_n246) );
  NAND2X0 r839_U249 ( .IN1(r839_n245), .IN2(r839_n246), .QN(r839_n239) );
  NAND2X0 r839_U248 ( .IN1(P2_N5082), .IN2(r839_n244), .QN(r839_n240) );
  OR2X1 r839_U247 ( .IN2(P2_N5082), .IN1(r839_n244), .Q(r839_n242) );
  NAND2X0 r839_U246 ( .IN1(r839_n242), .IN2(r839_n243), .QN(r839_n241) );
  NAND2X0 r839_U245 ( .IN1(r839_n240), .IN2(r839_n241), .QN(r839_n234) );
  NAND2X0 r839_U244 ( .IN1(r839_n239), .IN2(r839_n234), .QN(r839_n237) );
  OR2X1 r839_U243 ( .IN2(r839_n234), .IN1(r839_n239), .Q(r839_n238) );
  NAND2X0 r839_U242 ( .IN1(r839_n237), .IN2(r839_n238), .QN(P2_N1650) );
  INVX0 r839_U241 ( .ZN(r839_n223), .INP(P2_N1499) );
  NAND2X0 r839_U240 ( .IN1(P2_N5084), .IN2(r839_n223), .QN(r839_n235) );
  OR2X1 r839_U239 ( .IN2(P2_N5084), .IN1(r839_n223), .Q(r839_n236) );
  NAND2X0 r839_U238 ( .IN1(r839_n235), .IN2(r839_n236), .QN(r839_n229) );
  NAND2X0 r839_U237 ( .IN1(n7210), .IN2(r839_n234), .QN(r839_n230) );
  OR2X1 r839_U236 ( .IN2(n7210), .IN1(r839_n234), .Q(r839_n232) );
  NAND2X0 r839_U235 ( .IN1(r839_n232), .IN2(r839_n233), .QN(r839_n231) );
  NAND2X0 r839_U234 ( .IN1(r839_n230), .IN2(r839_n231), .QN(r839_n224) );
  NAND2X0 r839_U233 ( .IN1(r839_n229), .IN2(r839_n224), .QN(r839_n227) );
  OR2X1 r839_U232 ( .IN2(r839_n224), .IN1(r839_n229), .Q(r839_n228) );
  NAND2X0 r839_U231 ( .IN1(r839_n227), .IN2(r839_n228), .QN(P2_N1651) );
  INVX0 r839_U230 ( .ZN(r839_n213), .INP(P2_N1500) );
  NAND2X0 r839_U229 ( .IN1(P2_N5085), .IN2(r839_n213), .QN(r839_n225) );
  OR2X1 r839_U228 ( .IN2(P2_N5085), .IN1(r839_n213), .Q(r839_n226) );
  NAND2X0 r839_U227 ( .IN1(r839_n225), .IN2(r839_n226), .QN(r839_n219) );
  NAND2X0 r839_U226 ( .IN1(P2_N5084), .IN2(r839_n224), .QN(r839_n220) );
  OR2X1 r839_U225 ( .IN2(P2_N5084), .IN1(r839_n224), .Q(r839_n222) );
  NAND2X0 r839_U224 ( .IN1(r839_n222), .IN2(r839_n223), .QN(r839_n221) );
  NAND2X0 r839_U223 ( .IN1(r839_n220), .IN2(r839_n221), .QN(r839_n214) );
  NAND2X0 r839_U222 ( .IN1(r839_n219), .IN2(r839_n214), .QN(r839_n217) );
  OR2X1 r839_U221 ( .IN2(r839_n214), .IN1(r839_n219), .Q(r839_n218) );
  NAND2X0 r839_U220 ( .IN1(r839_n217), .IN2(r839_n218), .QN(P2_N1652) );
  INVX0 r839_U219 ( .ZN(r839_n203), .INP(P2_N1501) );
  NAND2X0 r839_U218 ( .IN1(P2_N5086), .IN2(r839_n203), .QN(r839_n215) );
  OR2X1 r839_U217 ( .IN2(P2_N5086), .IN1(r839_n203), .Q(r839_n216) );
  NAND2X0 r839_U216 ( .IN1(r839_n215), .IN2(r839_n216), .QN(r839_n209) );
  NAND2X0 r839_U215 ( .IN1(P2_N5085), .IN2(r839_n214), .QN(r839_n210) );
  OR2X1 r839_U214 ( .IN2(P2_N5085), .IN1(r839_n214), .Q(r839_n212) );
  NAND2X0 r839_U213 ( .IN1(r839_n212), .IN2(r839_n213), .QN(r839_n211) );
  NAND2X0 r839_U212 ( .IN1(r839_n210), .IN2(r839_n211), .QN(r839_n204) );
  NAND2X0 r839_U211 ( .IN1(r839_n209), .IN2(r839_n204), .QN(r839_n207) );
  OR2X1 r839_U210 ( .IN2(r839_n204), .IN1(r839_n209), .Q(r839_n208) );
  NAND2X0 r839_U209 ( .IN1(r839_n207), .IN2(r839_n208), .QN(P2_N1653) );
  INVX0 r839_U208 ( .ZN(r839_n193), .INP(P2_N1502) );
  NAND2X0 r839_U207 ( .IN1(n7198), .IN2(r839_n193), .QN(r839_n205) );
  OR2X1 r839_U206 ( .IN2(n7198), .IN1(r839_n193), .Q(r839_n206) );
  NAND2X0 r839_U205 ( .IN1(r839_n205), .IN2(r839_n206), .QN(r839_n199) );
  NAND2X0 r839_U204 ( .IN1(P2_N5086), .IN2(r839_n204), .QN(r839_n200) );
  OR2X1 r839_U203 ( .IN2(P2_N5086), .IN1(r839_n204), .Q(r839_n202) );
  NAND2X0 r839_U202 ( .IN1(r839_n202), .IN2(r839_n203), .QN(r839_n201) );
  NAND2X0 r839_U201 ( .IN1(r839_n200), .IN2(r839_n201), .QN(r839_n194) );
  NAND2X0 r839_U200 ( .IN1(r839_n199), .IN2(r839_n194), .QN(r839_n197) );
  OR2X1 r839_U199 ( .IN2(r839_n194), .IN1(r839_n199), .Q(r839_n198) );
  NAND2X0 r839_U198 ( .IN1(r839_n197), .IN2(r839_n198), .QN(P2_N1654) );
  INVX0 r839_U197 ( .ZN(r839_n183), .INP(P2_N1503) );
  NAND2X0 r839_U196 ( .IN1(n7194), .IN2(r839_n183), .QN(r839_n195) );
  OR2X1 r839_U195 ( .IN2(n7194), .IN1(r839_n183), .Q(r839_n196) );
  NAND2X0 r839_U194 ( .IN1(r839_n195), .IN2(r839_n196), .QN(r839_n189) );
  NAND2X0 r839_U193 ( .IN1(n7198), .IN2(r839_n194), .QN(r839_n190) );
  OR2X1 r839_U192 ( .IN2(n7198), .IN1(r839_n194), .Q(r839_n192) );
  NAND2X0 r839_U191 ( .IN1(r839_n192), .IN2(r839_n193), .QN(r839_n191) );
  NAND2X0 r839_U190 ( .IN1(r839_n190), .IN2(r839_n191), .QN(r839_n184) );
  NAND2X0 r839_U189 ( .IN1(r839_n189), .IN2(r839_n184), .QN(r839_n187) );
  OR2X1 r839_U188 ( .IN2(r839_n184), .IN1(r839_n189), .Q(r839_n188) );
  NAND2X0 r839_U187 ( .IN1(r839_n187), .IN2(r839_n188), .QN(P2_N1655) );
  INVX0 r839_U186 ( .ZN(r839_n173), .INP(P2_N1504) );
  NAND2X0 r839_U185 ( .IN1(n7187), .IN2(r839_n173), .QN(r839_n185) );
  OR2X1 r839_U184 ( .IN2(n7187), .IN1(r839_n173), .Q(r839_n186) );
  NAND2X0 r839_U183 ( .IN1(r839_n185), .IN2(r839_n186), .QN(r839_n179) );
  INVX0 r839_U321 ( .ZN(r839_n291), .INP(P2_N1486) );
  NOR2X0 r839_U320 ( .QN(r839_n287), .IN1(r839_n291), .IN2(n7035) );
  INVX0 r839_U319 ( .ZN(r839_n162), .INP(r839_n287) );
  NAND2X0 r839_U318 ( .IN1(n7035), .IN2(r839_n291), .QN(r839_n290) );
  NAND2X0 r839_U317 ( .IN1(r839_n162), .IN2(r839_n290), .QN(P2_N1638) );
  INVX0 r839_U316 ( .ZN(r839_n253), .INP(P2_N1496) );
  NAND2X0 r839_U315 ( .IN1(P2_N5081), .IN2(r839_n253), .QN(r839_n288) );
  OR2X1 r839_U314 ( .IN2(P2_N5081), .IN1(r839_n253), .Q(r839_n289) );
  NAND2X0 r839_U313 ( .IN1(r839_n288), .IN2(r839_n289), .QN(r839_n259) );
  NAND2X0 r839_U312 ( .IN1(P2_N5072), .IN2(r839_n162), .QN(r839_n284) );
  NAND2X0 r839_U310 ( .IN1(r839_n287), .IN2(n7184), .QN(r839_n286) );
  INVX0 r839_U309 ( .ZN(r839_n166), .INP(P2_N1487) );
  NAND2X0 r839_U308 ( .IN1(r839_n286), .IN2(r839_n166), .QN(r839_n285) );
  NAND2X0 r839_U307 ( .IN1(r839_n284), .IN2(r839_n285), .QN(r839_n53) );
  NAND2X0 r839_U306 ( .IN1(n7181), .IN2(r839_n53), .QN(r839_n281) );
  OR2X1 r839_U305 ( .IN2(P2_N5073), .IN1(r839_n53), .Q(r839_n283) );
  INVX0 r839_U304 ( .ZN(r839_n56), .INP(P2_N1488) );
  NAND2X0 r839_U303 ( .IN1(r839_n283), .IN2(r839_n56), .QN(r839_n282) );
  NAND2X0 r839_U302 ( .IN1(r839_n281), .IN2(r839_n282), .QN(r839_n46) );
  NAND2X0 r839_U301 ( .IN1(P2_N5074), .IN2(r839_n46), .QN(r839_n278) );
  OR2X1 r839_U300 ( .IN2(P2_N5074), .IN1(r839_n46), .Q(r839_n280) );
  INVX0 r839_U299 ( .ZN(r839_n49), .INP(P2_N1489) );
  NAND2X0 r839_U298 ( .IN1(r839_n280), .IN2(r839_n49), .QN(r839_n279) );
  NAND2X0 r839_U297 ( .IN1(r839_n278), .IN2(r839_n279), .QN(r839_n39) );
  NAND2X0 r839_U296 ( .IN1(P2_N5075), .IN2(r839_n39), .QN(r839_n275) );
  OR2X1 r839_U295 ( .IN2(P2_N5075), .IN1(r839_n39), .Q(r839_n277) );
  INVX0 r839_U294 ( .ZN(r839_n42), .INP(P2_N1490) );
  NAND2X0 r839_U293 ( .IN1(r839_n277), .IN2(r839_n42), .QN(r839_n276) );
  NAND2X0 r839_U292 ( .IN1(r839_n275), .IN2(r839_n276), .QN(r839_n32) );
  NAND2X0 r839_U291 ( .IN1(P2_N5076), .IN2(r839_n32), .QN(r839_n272) );
  OR2X1 r839_U290 ( .IN2(P2_N5076), .IN1(r839_n32), .Q(r839_n274) );
  INVX0 r839_U289 ( .ZN(r839_n35), .INP(P2_N1491) );
  NAND2X0 r839_U288 ( .IN1(r839_n274), .IN2(r839_n35), .QN(r839_n273) );
  NAND2X0 r839_U287 ( .IN1(r839_n272), .IN2(r839_n273), .QN(r839_n25) );
  NAND2X0 r839_U286 ( .IN1(n7162), .IN2(r839_n25), .QN(r839_n269) );
  OR2X1 r839_U285 ( .IN2(n7162), .IN1(r839_n25), .Q(r839_n271) );
  INVX0 r839_U284 ( .ZN(r839_n28), .INP(P2_N1492) );
  NAND2X0 r839_U283 ( .IN1(r839_n271), .IN2(r839_n28), .QN(r839_n270) );
  NAND2X0 r839_U282 ( .IN1(r839_n269), .IN2(r839_n270), .QN(r839_n18) );
  NAND2X0 r839_U281 ( .IN1(n7158), .IN2(r839_n18), .QN(r839_n266) );
  OR2X1 r839_U280 ( .IN2(n7158), .IN1(r839_n18), .Q(r839_n268) );
  INVX0 r839_U279 ( .ZN(r839_n21), .INP(P2_N1493) );
  NAND2X0 r839_U278 ( .IN1(r839_n268), .IN2(r839_n21), .QN(r839_n267) );
  NAND2X0 r839_U277 ( .IN1(r839_n266), .IN2(r839_n267), .QN(r839_n11) );
  NAND2X0 r839_U276 ( .IN1(P2_N5079), .IN2(r839_n11), .QN(r839_n263) );
  OR2X1 r841_U38 ( .IN2(r841_n46), .IN1(r841_n45), .Q(r841_n44) );
  NAND2X0 r841_U37 ( .IN1(r841_n43), .IN2(r841_n44), .QN(P2_N2014) );
  NAND2X0 r841_U36 ( .IN1(n7173), .IN2(r841_n42), .QN(r841_n40) );
  OR2X1 r841_U35 ( .IN2(n7173), .IN1(r841_n42), .Q(r841_n41) );
  NAND2X0 r841_U34 ( .IN1(r841_n40), .IN2(r841_n41), .QN(r841_n38) );
  NAND2X0 r841_U33 ( .IN1(r841_n38), .IN2(r841_n39), .QN(r841_n36) );
  OR2X1 r841_U32 ( .IN2(r841_n39), .IN1(r841_n38), .Q(r841_n37) );
  NAND2X0 r841_U31 ( .IN1(r841_n36), .IN2(r841_n37), .QN(P2_N2015) );
  NAND2X0 r841_U30 ( .IN1(n7165), .IN2(r841_n35), .QN(r841_n33) );
  OR2X1 r841_U29 ( .IN2(n7165), .IN1(r841_n35), .Q(r841_n34) );
  NAND2X0 r841_U28 ( .IN1(r841_n33), .IN2(r841_n34), .QN(r841_n31) );
  NAND2X0 r841_U27 ( .IN1(r841_n31), .IN2(r841_n32), .QN(r841_n29) );
  OR2X1 r841_U26 ( .IN2(r841_n32), .IN1(r841_n31), .Q(r841_n30) );
  NAND2X0 r841_U25 ( .IN1(r841_n29), .IN2(r841_n30), .QN(P2_N2016) );
  NAND2X0 r841_U24 ( .IN1(n7162), .IN2(r841_n28), .QN(r841_n26) );
  OR2X1 r841_U23 ( .IN2(n7162), .IN1(r841_n28), .Q(r841_n27) );
  NAND2X0 r841_U22 ( .IN1(r841_n26), .IN2(r841_n27), .QN(r841_n24) );
  NAND2X0 r841_U21 ( .IN1(r841_n24), .IN2(r841_n25), .QN(r841_n22) );
  OR2X1 r841_U20 ( .IN2(r841_n25), .IN1(r841_n24), .Q(r841_n23) );
  NAND2X0 r841_U19 ( .IN1(r841_n22), .IN2(r841_n23), .QN(P2_N2017) );
  NAND2X0 r841_U18 ( .IN1(n7158), .IN2(r841_n21), .QN(r841_n19) );
  OR2X1 r841_U17 ( .IN2(n7158), .IN1(r841_n21), .Q(r841_n20) );
  NAND2X0 r841_U16 ( .IN1(r841_n19), .IN2(r841_n20), .QN(r841_n17) );
  NAND2X0 r841_U15 ( .IN1(r841_n17), .IN2(r841_n18), .QN(r841_n15) );
  OR2X1 r841_U14 ( .IN2(r841_n18), .IN1(r841_n17), .Q(r841_n16) );
  NAND2X0 r841_U13 ( .IN1(r841_n15), .IN2(r841_n16), .QN(P2_N2018) );
  NAND2X0 r841_U12 ( .IN1(n7154), .IN2(r841_n14), .QN(r841_n12) );
  OR2X1 r841_U11 ( .IN2(n7154), .IN1(r841_n14), .Q(r841_n13) );
  NAND2X0 r841_U10 ( .IN1(r841_n12), .IN2(r841_n13), .QN(r841_n10) );
  NAND2X0 r841_U9 ( .IN1(r841_n10), .IN2(r841_n11), .QN(r841_n8) );
  OR2X1 r841_U8 ( .IN2(r841_n11), .IN1(r841_n10), .Q(r841_n9) );
  NAND2X0 r841_U7 ( .IN1(r841_n8), .IN2(r841_n9), .QN(P2_N2019) );
  NAND2X0 r841_U6 ( .IN1(P2_N5080), .IN2(r841_n7), .QN(r841_n5) );
  OR2X1 r841_U5 ( .IN2(P2_N5080), .IN1(r841_n7), .Q(r841_n6) );
  NAND2X0 r841_U4 ( .IN1(r841_n5), .IN2(r841_n6), .QN(r841_n3) );
  NAND2X0 r841_U3 ( .IN1(r841_n3), .IN2(r841_n4), .QN(r841_n1) );
  OR2X1 r841_U2 ( .IN2(r841_n4), .IN1(r841_n3), .Q(r841_n2) );
  NAND2X0 r841_U1 ( .IN1(r841_n1), .IN2(r841_n2), .QN(P2_N2020) );
  OR2X1 r841_U131 ( .IN2(n7252), .IN1(r841_n136), .Q(r841_n134) );
  NAND2X0 r841_U130 ( .IN1(r841_n134), .IN2(r841_n135), .QN(r841_n133) );
  NAND2X0 r841_U129 ( .IN1(r841_n132), .IN2(r841_n133), .QN(r841_n126) );
  NAND2X0 r841_U128 ( .IN1(r841_n131), .IN2(r841_n126), .QN(r841_n129) );
  OR2X1 r841_U127 ( .IN2(r841_n126), .IN1(r841_n131), .Q(r841_n130) );
  NAND2X0 r841_U126 ( .IN1(r841_n129), .IN2(r841_n130), .QN(P2_N2033) );
  INVX0 r841_U125 ( .ZN(r841_n115), .INP(P2_N1882) );
  NAND2X0 r841_U124 ( .IN1(n7242), .IN2(r841_n115), .QN(r841_n127) );
  OR2X1 r841_U123 ( .IN2(n7242), .IN1(r841_n115), .Q(r841_n128) );
  NAND2X0 r841_U122 ( .IN1(r841_n127), .IN2(r841_n128), .QN(r841_n121) );
  NAND2X0 r841_U121 ( .IN1(n7247), .IN2(r841_n126), .QN(r841_n122) );
  OR2X1 r841_U120 ( .IN2(n7247), .IN1(r841_n126), .Q(r841_n124) );
  NAND2X0 r841_U119 ( .IN1(r841_n124), .IN2(r841_n125), .QN(r841_n123) );
  NAND2X0 r841_U118 ( .IN1(r841_n122), .IN2(r841_n123), .QN(r841_n116) );
  NAND2X0 r841_U117 ( .IN1(r841_n121), .IN2(r841_n116), .QN(r841_n119) );
  OR2X1 r841_U116 ( .IN2(r841_n116), .IN1(r841_n121), .Q(r841_n120) );
  NAND2X0 r841_U115 ( .IN1(r841_n119), .IN2(r841_n120), .QN(P2_N2034) );
  INVX0 r841_U114 ( .ZN(r841_n105), .INP(P2_N1883) );
  NAND2X0 r841_U113 ( .IN1(n7238), .IN2(r841_n105), .QN(r841_n117) );
  OR2X1 r841_U112 ( .IN2(n7238), .IN1(r841_n105), .Q(r841_n118) );
  NAND2X0 r841_U111 ( .IN1(r841_n117), .IN2(r841_n118), .QN(r841_n111) );
  NAND2X0 r841_U110 ( .IN1(n7242), .IN2(r841_n116), .QN(r841_n112) );
  OR2X1 r841_U109 ( .IN2(n7242), .IN1(r841_n116), .Q(r841_n114) );
  NAND2X0 r841_U108 ( .IN1(r841_n114), .IN2(r841_n115), .QN(r841_n113) );
  NAND2X0 r841_U107 ( .IN1(r841_n112), .IN2(r841_n113), .QN(r841_n106) );
  NAND2X0 r841_U106 ( .IN1(r841_n111), .IN2(r841_n106), .QN(r841_n109) );
  OR2X1 r841_U105 ( .IN2(r841_n106), .IN1(r841_n111), .Q(r841_n110) );
  NAND2X0 r841_U104 ( .IN1(r841_n109), .IN2(r841_n110), .QN(P2_N2035) );
  INVX0 r841_U103 ( .ZN(r841_n95), .INP(P2_N1884) );
  NAND2X0 r841_U102 ( .IN1(P2_N5096), .IN2(r841_n95), .QN(r841_n107) );
  OR2X1 r841_U101 ( .IN2(P2_N5096), .IN1(r841_n95), .Q(r841_n108) );
  NAND2X0 r841_U100 ( .IN1(r841_n107), .IN2(r841_n108), .QN(r841_n101) );
  NAND2X0 r841_U99 ( .IN1(n7238), .IN2(r841_n106), .QN(r841_n102) );
  OR2X1 r841_U98 ( .IN2(n7238), .IN1(r841_n106), .Q(r841_n104) );
  NAND2X0 r841_U97 ( .IN1(r841_n104), .IN2(r841_n105), .QN(r841_n103) );
  NAND2X0 r841_U96 ( .IN1(r841_n102), .IN2(r841_n103), .QN(r841_n96) );
  NAND2X0 r841_U95 ( .IN1(r841_n101), .IN2(r841_n96), .QN(r841_n99) );
  OR2X1 r841_U94 ( .IN2(r841_n96), .IN1(r841_n101), .Q(r841_n100) );
  NAND2X0 r841_U93 ( .IN1(r841_n99), .IN2(r841_n100), .QN(P2_N2036) );
  INVX0 r841_U92 ( .ZN(r841_n85), .INP(P2_N1885) );
  NAND2X0 r841_U91 ( .IN1(P2_N5097), .IN2(r841_n85), .QN(r841_n97) );
  OR2X1 r841_U90 ( .IN2(P2_N5097), .IN1(r841_n85), .Q(r841_n98) );
  NAND2X0 r841_U89 ( .IN1(r841_n97), .IN2(r841_n98), .QN(r841_n91) );
  NAND2X0 r841_U88 ( .IN1(P2_N5096), .IN2(r841_n96), .QN(r841_n92) );
  OR2X1 r841_U87 ( .IN2(P2_N5096), .IN1(r841_n96), .Q(r841_n94) );
  NAND2X0 r841_U86 ( .IN1(r841_n94), .IN2(r841_n95), .QN(r841_n93) );
  NAND2X0 r841_U85 ( .IN1(r841_n92), .IN2(r841_n93), .QN(r841_n86) );
  NAND2X0 r841_U84 ( .IN1(r841_n91), .IN2(r841_n86), .QN(r841_n89) );
  OR2X1 r841_U83 ( .IN2(r841_n86), .IN1(r841_n91), .Q(r841_n90) );
  NAND2X0 r841_U82 ( .IN1(r841_n89), .IN2(r841_n90), .QN(P2_N2037) );
  INVX0 r841_U81 ( .ZN(r841_n75), .INP(P2_N1886) );
  NAND2X0 r841_U80 ( .IN1(n7227), .IN2(r841_n75), .QN(r841_n87) );
  OR2X1 r841_U79 ( .IN2(n7227), .IN1(r841_n75), .Q(r841_n88) );
  NAND2X0 r841_U78 ( .IN1(r841_n87), .IN2(r841_n88), .QN(r841_n81) );
  NAND2X0 r841_U77 ( .IN1(P2_N5097), .IN2(r841_n86), .QN(r841_n82) );
  OR2X1 r841_U76 ( .IN2(P2_N5097), .IN1(r841_n86), .Q(r841_n84) );
  NAND2X0 r841_U75 ( .IN1(r841_n84), .IN2(r841_n85), .QN(r841_n83) );
  NAND2X0 r841_U74 ( .IN1(r841_n82), .IN2(r841_n83), .QN(r841_n76) );
  NAND2X0 r841_U73 ( .IN1(r841_n81), .IN2(r841_n76), .QN(r841_n79) );
  OR2X1 r841_U72 ( .IN2(r841_n76), .IN1(r841_n81), .Q(r841_n80) );
  NAND2X0 r841_U71 ( .IN1(r841_n79), .IN2(r841_n80), .QN(P2_N2038) );
  INVX0 r841_U70 ( .ZN(r841_n64), .INP(P2_N1887) );
  NAND2X0 r841_U69 ( .IN1(P2_N5099), .IN2(r841_n64), .QN(r841_n77) );
  OR2X1 r841_U68 ( .IN2(P2_N5099), .IN1(r841_n64), .Q(r841_n78) );
  NAND2X0 r841_U67 ( .IN1(r841_n77), .IN2(r841_n78), .QN(r841_n71) );
  NAND2X0 r841_U66 ( .IN1(n7227), .IN2(r841_n76), .QN(r841_n72) );
  OR2X1 r841_U65 ( .IN2(n7227), .IN1(r841_n76), .Q(r841_n74) );
  NAND2X0 r841_U64 ( .IN1(r841_n74), .IN2(r841_n75), .QN(r841_n73) );
  NAND2X0 r841_U63 ( .IN1(r841_n72), .IN2(r841_n73), .QN(r841_n65) );
  NAND2X0 r841_U62 ( .IN1(r841_n71), .IN2(r841_n65), .QN(r841_n69) );
  OR2X1 r841_U61 ( .IN2(r841_n65), .IN1(r841_n71), .Q(r841_n70) );
  NAND2X0 r841_U60 ( .IN1(r841_n69), .IN2(r841_n70), .QN(P2_N2039) );
  OR2X1 r841_U58 ( .IN2(P2_N1888), .IN1(n7266), .Q(r841_n66) );
  NAND2X0 r841_U57 ( .IN1(P2_N1888), .IN2(n7266), .QN(r841_n67) );
  NAND2X0 r841_U56 ( .IN1(r841_n66), .IN2(r841_n67), .QN(r841_n60) );
  NAND2X0 r841_U55 ( .IN1(P2_N5099), .IN2(r841_n65), .QN(r841_n61) );
  OR2X1 r841_U54 ( .IN2(P2_N5099), .IN1(r841_n65), .Q(r841_n63) );
  NAND2X0 r841_U53 ( .IN1(r841_n63), .IN2(r841_n64), .QN(r841_n62) );
  NAND2X0 r841_U52 ( .IN1(r841_n61), .IN2(r841_n62), .QN(r841_n59) );
  NAND2X0 r841_U51 ( .IN1(r841_n60), .IN2(r841_n59), .QN(r841_n57) );
  OR2X1 r841_U50 ( .IN2(r841_n60), .IN1(r841_n59), .Q(r841_n58) );
  NAND2X0 r841_U49 ( .IN1(r841_n57), .IN2(r841_n58), .QN(P2_N2040) );
  NAND2X0 r841_U48 ( .IN1(n7181), .IN2(r841_n56), .QN(r841_n54) );
  OR2X1 r841_U47 ( .IN2(n7181), .IN1(r841_n56), .Q(r841_n55) );
  NAND2X0 r841_U46 ( .IN1(r841_n54), .IN2(r841_n55), .QN(r841_n52) );
  NAND2X0 r841_U45 ( .IN1(r841_n52), .IN2(r841_n53), .QN(r841_n50) );
  OR2X1 r841_U44 ( .IN2(r841_n53), .IN1(r841_n52), .Q(r841_n51) );
  NAND2X0 r841_U43 ( .IN1(r841_n50), .IN2(r841_n51), .QN(P2_N2013) );
  NAND2X0 r841_U42 ( .IN1(n7177), .IN2(r841_n49), .QN(r841_n47) );
  OR2X1 r841_U41 ( .IN2(n7177), .IN1(r841_n49), .Q(r841_n48) );
  NAND2X0 r841_U40 ( .IN1(r841_n47), .IN2(r841_n48), .QN(r841_n45) );
  NAND2X0 r841_U39 ( .IN1(r841_n45), .IN2(r841_n46), .QN(r841_n43) );
  NAND2X0 r841_U224 ( .IN1(r841_n222), .IN2(r841_n223), .QN(r841_n221) );
  NAND2X0 r841_U223 ( .IN1(r841_n220), .IN2(r841_n221), .QN(r841_n214) );
  NAND2X0 r841_U222 ( .IN1(r841_n219), .IN2(r841_n214), .QN(r841_n217) );
  OR2X1 r841_U221 ( .IN2(r841_n214), .IN1(r841_n219), .Q(r841_n218) );
  NAND2X0 r841_U220 ( .IN1(r841_n217), .IN2(r841_n218), .QN(P2_N2025) );
  INVX0 r841_U219 ( .ZN(r841_n203), .INP(P2_N1874) );
  NAND2X0 r841_U218 ( .IN1(n7202), .IN2(r841_n203), .QN(r841_n215) );
  OR2X1 r841_U217 ( .IN2(n7202), .IN1(r841_n203), .Q(r841_n216) );
  NAND2X0 r841_U216 ( .IN1(r841_n215), .IN2(r841_n216), .QN(r841_n209) );
  NAND2X0 r841_U215 ( .IN1(P2_N5085), .IN2(r841_n214), .QN(r841_n210) );
  OR2X1 r841_U214 ( .IN2(P2_N5085), .IN1(r841_n214), .Q(r841_n212) );
  NAND2X0 r841_U213 ( .IN1(r841_n212), .IN2(r841_n213), .QN(r841_n211) );
  NAND2X0 r841_U212 ( .IN1(r841_n210), .IN2(r841_n211), .QN(r841_n204) );
  NAND2X0 r841_U211 ( .IN1(r841_n209), .IN2(r841_n204), .QN(r841_n207) );
  OR2X1 r841_U210 ( .IN2(r841_n204), .IN1(r841_n209), .Q(r841_n208) );
  NAND2X0 r841_U209 ( .IN1(r841_n207), .IN2(r841_n208), .QN(P2_N2026) );
  INVX0 r841_U208 ( .ZN(r841_n193), .INP(P2_N1875) );
  NAND2X0 r841_U207 ( .IN1(P2_N5087), .IN2(r841_n193), .QN(r841_n205) );
  OR2X1 r841_U206 ( .IN2(P2_N5087), .IN1(r841_n193), .Q(r841_n206) );
  NAND2X0 r841_U205 ( .IN1(r841_n205), .IN2(r841_n206), .QN(r841_n199) );
  NAND2X0 r841_U204 ( .IN1(n7202), .IN2(r841_n204), .QN(r841_n200) );
  OR2X1 r841_U203 ( .IN2(n7202), .IN1(r841_n204), .Q(r841_n202) );
  NAND2X0 r841_U202 ( .IN1(r841_n202), .IN2(r841_n203), .QN(r841_n201) );
  NAND2X0 r841_U201 ( .IN1(r841_n200), .IN2(r841_n201), .QN(r841_n194) );
  NAND2X0 r841_U200 ( .IN1(r841_n199), .IN2(r841_n194), .QN(r841_n197) );
  OR2X1 r841_U199 ( .IN2(r841_n194), .IN1(r841_n199), .Q(r841_n198) );
  NAND2X0 r841_U198 ( .IN1(r841_n197), .IN2(r841_n198), .QN(P2_N2027) );
  INVX0 r841_U197 ( .ZN(r841_n183), .INP(P2_N1876) );
  NAND2X0 r841_U196 ( .IN1(P2_N5088), .IN2(r841_n183), .QN(r841_n195) );
  OR2X1 r841_U195 ( .IN2(P2_N5088), .IN1(r841_n183), .Q(r841_n196) );
  NAND2X0 r841_U194 ( .IN1(r841_n195), .IN2(r841_n196), .QN(r841_n189) );
  NAND2X0 r841_U193 ( .IN1(P2_N5087), .IN2(r841_n194), .QN(r841_n190) );
  OR2X1 r841_U192 ( .IN2(P2_N5087), .IN1(r841_n194), .Q(r841_n192) );
  NAND2X0 r841_U191 ( .IN1(r841_n192), .IN2(r841_n193), .QN(r841_n191) );
  NAND2X0 r841_U190 ( .IN1(r841_n190), .IN2(r841_n191), .QN(r841_n184) );
  NAND2X0 r841_U189 ( .IN1(r841_n189), .IN2(r841_n184), .QN(r841_n187) );
  OR2X1 r841_U188 ( .IN2(r841_n184), .IN1(r841_n189), .Q(r841_n188) );
  NAND2X0 r841_U187 ( .IN1(r841_n187), .IN2(r841_n188), .QN(P2_N2028) );
  INVX0 r841_U186 ( .ZN(r841_n173), .INP(P2_N1877) );
  NAND2X0 r841_U185 ( .IN1(P2_N5089), .IN2(r841_n173), .QN(r841_n185) );
  OR2X1 r841_U184 ( .IN2(P2_N5089), .IN1(r841_n173), .Q(r841_n186) );
  NAND2X0 r841_U183 ( .IN1(r841_n185), .IN2(r841_n186), .QN(r841_n179) );
  NAND2X0 r841_U182 ( .IN1(P2_N5088), .IN2(r841_n184), .QN(r841_n180) );
  OR2X1 r841_U181 ( .IN2(P2_N5088), .IN1(r841_n184), .Q(r841_n182) );
  NAND2X0 r841_U180 ( .IN1(r841_n182), .IN2(r841_n183), .QN(r841_n181) );
  NAND2X0 r841_U179 ( .IN1(r841_n180), .IN2(r841_n181), .QN(r841_n174) );
  NAND2X0 r841_U178 ( .IN1(r841_n179), .IN2(r841_n174), .QN(r841_n177) );
  OR2X1 r841_U177 ( .IN2(r841_n174), .IN1(r841_n179), .Q(r841_n178) );
  NAND2X0 r841_U176 ( .IN1(r841_n177), .IN2(r841_n178), .QN(P2_N2029) );
  INVX0 r841_U175 ( .ZN(r841_n155), .INP(P2_N1878) );
  NAND2X0 r841_U174 ( .IN1(n7263), .IN2(r841_n155), .QN(r841_n175) );
  OR2X1 r841_U173 ( .IN2(n7263), .IN1(r841_n155), .Q(r841_n176) );
  NAND2X0 r841_U172 ( .IN1(r841_n175), .IN2(r841_n176), .QN(r841_n169) );
  NAND2X0 r841_U171 ( .IN1(P2_N5089), .IN2(r841_n174), .QN(r841_n170) );
  OR2X1 r841_U170 ( .IN2(P2_N5089), .IN1(r841_n174), .Q(r841_n172) );
  NAND2X0 r841_U169 ( .IN1(r841_n172), .IN2(r841_n173), .QN(r841_n171) );
  NAND2X0 r841_U168 ( .IN1(r841_n170), .IN2(r841_n171), .QN(r841_n156) );
  NAND2X0 r841_U167 ( .IN1(r841_n169), .IN2(r841_n156), .QN(r841_n167) );
  OR2X1 r841_U166 ( .IN2(r841_n156), .IN1(r841_n169), .Q(r841_n168) );
  NAND2X0 r841_U165 ( .IN1(r841_n167), .IN2(r841_n168), .QN(P2_N2030) );
  NAND2X0 r841_U164 ( .IN1(P2_N5072), .IN2(r841_n166), .QN(r841_n163) );
  NAND2X0 r841_U163 ( .IN1(P2_N1860), .IN2(n7186), .QN(r841_n164) );
  NAND2X0 r841_U162 ( .IN1(r841_n163), .IN2(r841_n164), .QN(r841_n161) );
  NAND2X0 r841_U161 ( .IN1(r841_n161), .IN2(r841_n162), .QN(r841_n159) );
  OR2X1 r841_U160 ( .IN2(r841_n162), .IN1(r841_n161), .Q(r841_n160) );
  NAND2X0 r841_U159 ( .IN1(r841_n159), .IN2(r841_n160), .QN(P2_N2012) );
  INVX0 r841_U158 ( .ZN(r841_n145), .INP(P2_N1879) );
  NAND2X0 r841_U157 ( .IN1(n7259), .IN2(r841_n145), .QN(r841_n157) );
  OR2X1 r841_U156 ( .IN2(n7259), .IN1(r841_n145), .Q(r841_n158) );
  NAND2X0 r841_U155 ( .IN1(r841_n157), .IN2(r841_n158), .QN(r841_n151) );
  NAND2X0 r841_U154 ( .IN1(n7263), .IN2(r841_n156), .QN(r841_n152) );
  OR2X1 r841_U153 ( .IN2(n7263), .IN1(r841_n156), .Q(r841_n154) );
  NAND2X0 r841_U152 ( .IN1(r841_n154), .IN2(r841_n155), .QN(r841_n153) );
  NAND2X0 r841_U151 ( .IN1(r841_n152), .IN2(r841_n153), .QN(r841_n146) );
  NAND2X0 r841_U150 ( .IN1(r841_n151), .IN2(r841_n146), .QN(r841_n149) );
  OR2X1 r841_U149 ( .IN2(r841_n146), .IN1(r841_n151), .Q(r841_n150) );
  NAND2X0 r841_U148 ( .IN1(r841_n149), .IN2(r841_n150), .QN(P2_N2031) );
  INVX0 r841_U147 ( .ZN(r841_n135), .INP(P2_N1880) );
  NAND2X0 r841_U146 ( .IN1(n7252), .IN2(r841_n135), .QN(r841_n147) );
  OR2X1 r841_U145 ( .IN2(n7252), .IN1(r841_n135), .Q(r841_n148) );
  NAND2X0 r841_U144 ( .IN1(r841_n147), .IN2(r841_n148), .QN(r841_n141) );
  NAND2X0 r841_U143 ( .IN1(n7259), .IN2(r841_n146), .QN(r841_n142) );
  OR2X1 r841_U142 ( .IN2(n7259), .IN1(r841_n146), .Q(r841_n144) );
  NAND2X0 r841_U141 ( .IN1(r841_n144), .IN2(r841_n145), .QN(r841_n143) );
  NAND2X0 r841_U140 ( .IN1(r841_n142), .IN2(r841_n143), .QN(r841_n136) );
  NAND2X0 r841_U139 ( .IN1(r841_n141), .IN2(r841_n136), .QN(r841_n139) );
  OR2X1 r841_U138 ( .IN2(r841_n136), .IN1(r841_n141), .Q(r841_n140) );
  NAND2X0 r841_U137 ( .IN1(r841_n139), .IN2(r841_n140), .QN(P2_N2032) );
  INVX0 r841_U136 ( .ZN(r841_n125), .INP(P2_N1881) );
  NAND2X0 r841_U135 ( .IN1(n7247), .IN2(r841_n125), .QN(r841_n137) );
  OR2X1 r841_U134 ( .IN2(n7247), .IN1(r841_n125), .Q(r841_n138) );
  NAND2X0 r841_U133 ( .IN1(r841_n137), .IN2(r841_n138), .QN(r841_n131) );
  NAND2X0 r841_U132 ( .IN1(n7252), .IN2(r841_n136), .QN(r841_n132) );
  NAND2X0 r841_U317 ( .IN1(r841_n162), .IN2(r841_n290), .QN(P2_N2011) );
  INVX0 r841_U316 ( .ZN(r841_n253), .INP(P2_N1869) );
  NAND2X0 r841_U315 ( .IN1(P2_N5081), .IN2(r841_n253), .QN(r841_n288) );
  OR2X1 r841_U314 ( .IN2(P2_N5081), .IN1(r841_n253), .Q(r841_n289) );
  NAND2X0 r841_U313 ( .IN1(r841_n288), .IN2(r841_n289), .QN(r841_n259) );
  NAND2X0 r841_U312 ( .IN1(P2_N5072), .IN2(r841_n162), .QN(r841_n284) );
  NAND2X0 r841_U310 ( .IN1(r841_n287), .IN2(n7186), .QN(r841_n286) );
  INVX0 r841_U309 ( .ZN(r841_n166), .INP(P2_N1860) );
  NAND2X0 r841_U308 ( .IN1(r841_n286), .IN2(r841_n166), .QN(r841_n285) );
  NAND2X0 r841_U307 ( .IN1(r841_n284), .IN2(r841_n285), .QN(r841_n53) );
  NAND2X0 r841_U306 ( .IN1(n7181), .IN2(r841_n53), .QN(r841_n281) );
  OR2X1 r841_U305 ( .IN2(n7181), .IN1(r841_n53), .Q(r841_n283) );
  INVX0 r841_U304 ( .ZN(r841_n56), .INP(P2_N1861) );
  NAND2X0 r841_U303 ( .IN1(r841_n283), .IN2(r841_n56), .QN(r841_n282) );
  NAND2X0 r841_U302 ( .IN1(r841_n281), .IN2(r841_n282), .QN(r841_n46) );
  NAND2X0 r841_U301 ( .IN1(n7177), .IN2(r841_n46), .QN(r841_n278) );
  OR2X1 r841_U300 ( .IN2(n7177), .IN1(r841_n46), .Q(r841_n280) );
  INVX0 r841_U299 ( .ZN(r841_n49), .INP(P2_N1862) );
  NAND2X0 r841_U298 ( .IN1(r841_n280), .IN2(r841_n49), .QN(r841_n279) );
  NAND2X0 r841_U297 ( .IN1(r841_n278), .IN2(r841_n279), .QN(r841_n39) );
  NAND2X0 r841_U296 ( .IN1(n7173), .IN2(r841_n39), .QN(r841_n275) );
  OR2X1 r841_U295 ( .IN2(n7173), .IN1(r841_n39), .Q(r841_n277) );
  INVX0 r841_U294 ( .ZN(r841_n42), .INP(P2_N1863) );
  NAND2X0 r841_U293 ( .IN1(r841_n277), .IN2(r841_n42), .QN(r841_n276) );
  NAND2X0 r841_U292 ( .IN1(r841_n275), .IN2(r841_n276), .QN(r841_n32) );
  NAND2X0 r841_U291 ( .IN1(n7165), .IN2(r841_n32), .QN(r841_n272) );
  OR2X1 r841_U290 ( .IN2(n7165), .IN1(r841_n32), .Q(r841_n274) );
  INVX0 r841_U289 ( .ZN(r841_n35), .INP(P2_N1864) );
  NAND2X0 r841_U288 ( .IN1(r841_n274), .IN2(r841_n35), .QN(r841_n273) );
  NAND2X0 r841_U287 ( .IN1(r841_n272), .IN2(r841_n273), .QN(r841_n25) );
  NAND2X0 r841_U286 ( .IN1(n7162), .IN2(r841_n25), .QN(r841_n269) );
  OR2X1 r841_U285 ( .IN2(n7162), .IN1(r841_n25), .Q(r841_n271) );
  INVX0 r841_U284 ( .ZN(r841_n28), .INP(P2_N1865) );
  NAND2X0 r841_U283 ( .IN1(r841_n271), .IN2(r841_n28), .QN(r841_n270) );
  NAND2X0 r841_U282 ( .IN1(r841_n269), .IN2(r841_n270), .QN(r841_n18) );
  NAND2X0 r841_U281 ( .IN1(n7158), .IN2(r841_n18), .QN(r841_n266) );
  OR2X1 r841_U280 ( .IN2(n7158), .IN1(r841_n18), .Q(r841_n268) );
  INVX0 r841_U279 ( .ZN(r841_n21), .INP(P2_N1866) );
  NAND2X0 r841_U278 ( .IN1(r841_n268), .IN2(r841_n21), .QN(r841_n267) );
  NAND2X0 r841_U277 ( .IN1(r841_n266), .IN2(r841_n267), .QN(r841_n11) );
  NAND2X0 r841_U276 ( .IN1(n7154), .IN2(r841_n11), .QN(r841_n263) );
  OR2X1 r841_U275 ( .IN2(n7154), .IN1(r841_n11), .Q(r841_n265) );
  INVX0 r841_U274 ( .ZN(r841_n14), .INP(P2_N1867) );
  NAND2X0 r841_U273 ( .IN1(r841_n265), .IN2(r841_n14), .QN(r841_n264) );
  NAND2X0 r841_U272 ( .IN1(r841_n263), .IN2(r841_n264), .QN(r841_n4) );
  NAND2X0 r841_U271 ( .IN1(P2_N5080), .IN2(r841_n4), .QN(r841_n260) );
  OR2X1 r841_U270 ( .IN2(P2_N5080), .IN1(r841_n4), .Q(r841_n262) );
  INVX0 r841_U269 ( .ZN(r841_n7), .INP(P2_N1868) );
  NAND2X0 r841_U268 ( .IN1(r841_n262), .IN2(r841_n7), .QN(r841_n261) );
  NAND2X0 r841_U267 ( .IN1(r841_n260), .IN2(r841_n261), .QN(r841_n254) );
  NAND2X0 r841_U266 ( .IN1(r841_n259), .IN2(r841_n254), .QN(r841_n257) );
  OR2X1 r841_U265 ( .IN2(r841_n254), .IN1(r841_n259), .Q(r841_n258) );
  NAND2X0 r841_U264 ( .IN1(r841_n257), .IN2(r841_n258), .QN(P2_N2021) );
  INVX0 r841_U263 ( .ZN(r841_n243), .INP(P2_N1870) );
  NAND2X0 r841_U262 ( .IN1(n7216), .IN2(r841_n243), .QN(r841_n255) );
  OR2X1 r841_U261 ( .IN2(n7216), .IN1(r841_n243), .Q(r841_n256) );
  NAND2X0 r841_U260 ( .IN1(r841_n255), .IN2(r841_n256), .QN(r841_n249) );
  NAND2X0 r841_U259 ( .IN1(P2_N5081), .IN2(r841_n254), .QN(r841_n250) );
  OR2X1 r841_U258 ( .IN2(P2_N5081), .IN1(r841_n254), .Q(r841_n252) );
  NAND2X0 r841_U257 ( .IN1(r841_n252), .IN2(r841_n253), .QN(r841_n251) );
  NAND2X0 r841_U256 ( .IN1(r841_n250), .IN2(r841_n251), .QN(r841_n244) );
  NAND2X0 r841_U255 ( .IN1(r841_n249), .IN2(r841_n244), .QN(r841_n247) );
  OR2X1 r841_U254 ( .IN2(r841_n244), .IN1(r841_n249), .Q(r841_n248) );
  NAND2X0 r841_U253 ( .IN1(r841_n247), .IN2(r841_n248), .QN(P2_N2022) );
  INVX0 r841_U252 ( .ZN(r841_n233), .INP(P2_N1871) );
  NAND2X0 r841_U251 ( .IN1(n7210), .IN2(r841_n233), .QN(r841_n245) );
  OR2X1 r841_U250 ( .IN2(n7210), .IN1(r841_n233), .Q(r841_n246) );
  NAND2X0 r841_U249 ( .IN1(r841_n245), .IN2(r841_n246), .QN(r841_n239) );
  NAND2X0 r841_U248 ( .IN1(n7216), .IN2(r841_n244), .QN(r841_n240) );
  OR2X1 r841_U247 ( .IN2(n7216), .IN1(r841_n244), .Q(r841_n242) );
  NAND2X0 r841_U246 ( .IN1(r841_n242), .IN2(r841_n243), .QN(r841_n241) );
  NAND2X0 r841_U245 ( .IN1(r841_n240), .IN2(r841_n241), .QN(r841_n234) );
  NAND2X0 r841_U244 ( .IN1(r841_n239), .IN2(r841_n234), .QN(r841_n237) );
  OR2X1 r841_U243 ( .IN2(r841_n234), .IN1(r841_n239), .Q(r841_n238) );
  NAND2X0 r841_U242 ( .IN1(r841_n237), .IN2(r841_n238), .QN(P2_N2023) );
  INVX0 r841_U241 ( .ZN(r841_n223), .INP(P2_N1872) );
  NAND2X0 r841_U240 ( .IN1(P2_N5084), .IN2(r841_n223), .QN(r841_n235) );
  OR2X1 r841_U239 ( .IN2(P2_N5084), .IN1(r841_n223), .Q(r841_n236) );
  NAND2X0 r841_U238 ( .IN1(r841_n235), .IN2(r841_n236), .QN(r841_n229) );
  NAND2X0 r841_U237 ( .IN1(n7210), .IN2(r841_n234), .QN(r841_n230) );
  OR2X1 r841_U236 ( .IN2(n7210), .IN1(r841_n234), .Q(r841_n232) );
  NAND2X0 r841_U235 ( .IN1(r841_n232), .IN2(r841_n233), .QN(r841_n231) );
  NAND2X0 r841_U234 ( .IN1(r841_n230), .IN2(r841_n231), .QN(r841_n224) );
  NAND2X0 r841_U233 ( .IN1(r841_n229), .IN2(r841_n224), .QN(r841_n227) );
  OR2X1 r841_U232 ( .IN2(r841_n224), .IN1(r841_n229), .Q(r841_n228) );
  NAND2X0 r841_U231 ( .IN1(r841_n227), .IN2(r841_n228), .QN(P2_N2024) );
  INVX0 r841_U230 ( .ZN(r841_n213), .INP(P2_N1873) );
  NAND2X0 r841_U229 ( .IN1(P2_N5085), .IN2(r841_n213), .QN(r841_n225) );
  OR2X1 r841_U228 ( .IN2(P2_N5085), .IN1(r841_n213), .Q(r841_n226) );
  NAND2X0 r841_U227 ( .IN1(r841_n225), .IN2(r841_n226), .QN(r841_n219) );
  NAND2X0 r841_U226 ( .IN1(P2_N5084), .IN2(r841_n224), .QN(r841_n220) );
  OR2X1 r841_U225 ( .IN2(P2_N5084), .IN1(r841_n224), .Q(r841_n222) );
  INVX0 r841_U321 ( .ZN(r841_n291), .INP(P2_N1859) );
  NOR2X0 r841_U320 ( .QN(r841_n287), .IN1(r841_n291), .IN2(n7035) );
  INVX0 r841_U319 ( .ZN(r841_n162), .INP(r841_n287) );
  NAND2X0 r841_U318 ( .IN1(n7035), .IN2(r841_n291), .QN(r841_n290) );
  NOR2X0 r843_U79 ( .QN(P2_N2411), .IN1(r843_n78), .IN2(r843_n79) );
  NAND2X0 r843_U78 ( .IN1(n7227), .IN2(r843_n77), .QN(r843_n74) );
  OR2X1 r843_U77 ( .IN2(n7227), .IN1(r843_n77), .Q(r843_n76) );
  NAND2X0 r843_U76 ( .IN1(P2_N2259), .IN2(r843_n76), .QN(r843_n75) );
  NAND2X0 r843_U75 ( .IN1(r843_n74), .IN2(r843_n75), .QN(r843_n64) );
  OR2X1 r843_U73 ( .IN2(P2_N2260), .IN1(n7222), .Q(r843_n71) );
  NAND2X0 r843_U72 ( .IN1(P2_N2260), .IN2(n7222), .QN(r843_n72) );
  NAND2X0 r843_U71 ( .IN1(r843_n71), .IN2(r843_n72), .QN(r843_n70) );
  NOR2X0 r843_U70 ( .QN(r843_n68), .IN1(r843_n64), .IN2(r843_n70) );
  AND2X1 r843_U69 ( .IN1(r843_n64), .IN2(r843_n70), .Q(r843_n69) );
  NOR2X0 r843_U68 ( .QN(P2_N2412), .IN1(r843_n68), .IN2(r843_n69) );
  OR2X1 r843_U66 ( .IN2(P2_N2261), .IN1(n7266), .Q(r843_n65) );
  NAND2X0 r843_U65 ( .IN1(P2_N2261), .IN2(n7266), .QN(r843_n66) );
  NAND2X0 r843_U64 ( .IN1(r843_n65), .IN2(r843_n66), .QN(r843_n60) );
  NAND2X0 r843_U63 ( .IN1(P2_N5099), .IN2(r843_n64), .QN(r843_n61) );
  OR2X1 r843_U62 ( .IN2(P2_N5099), .IN1(r843_n64), .Q(r843_n63) );
  NAND2X0 r843_U61 ( .IN1(P2_N2260), .IN2(r843_n63), .QN(r843_n62) );
  NAND2X0 r843_U60 ( .IN1(r843_n61), .IN2(r843_n62), .QN(r843_n59) );
  NOR2X0 r843_U59 ( .QN(r843_n57), .IN1(r843_n60), .IN2(r843_n59) );
  AND2X1 r843_U58 ( .IN1(r843_n59), .IN2(r843_n60), .Q(r843_n58) );
  NOR2X0 r843_U57 ( .QN(P2_N2413), .IN1(r843_n57), .IN2(r843_n58) );
  OR2X1 r843_U55 ( .IN2(P2_N2234), .IN1(n7182), .Q(r843_n54) );
  NAND2X0 r843_U54 ( .IN1(P2_N2234), .IN2(n7182), .QN(r843_n55) );
  NAND2X0 r843_U53 ( .IN1(r843_n54), .IN2(r843_n55), .QN(r843_n53) );
  NOR2X0 r843_U52 ( .QN(r843_n50), .IN1(r843_n52), .IN2(r843_n53) );
  AND2X1 r843_U51 ( .IN1(r843_n52), .IN2(r843_n53), .Q(r843_n51) );
  NOR2X0 r843_U50 ( .QN(P2_N2386), .IN1(r843_n50), .IN2(r843_n51) );
  OR2X1 r843_U48 ( .IN2(P2_N2235), .IN1(n7178), .Q(r843_n47) );
  NAND2X0 r843_U47 ( .IN1(P2_N2235), .IN2(n7178), .QN(r843_n48) );
  NAND2X0 r843_U46 ( .IN1(r843_n47), .IN2(r843_n48), .QN(r843_n46) );
  NOR2X0 r843_U45 ( .QN(r843_n43), .IN1(r843_n45), .IN2(r843_n46) );
  AND2X1 r843_U44 ( .IN1(r843_n45), .IN2(r843_n46), .Q(r843_n44) );
  NOR2X0 r843_U43 ( .QN(P2_N2387), .IN1(r843_n43), .IN2(r843_n44) );
  OR2X1 r843_U41 ( .IN2(P2_N2236), .IN1(n7174), .Q(r843_n40) );
  NAND2X0 r843_U40 ( .IN1(P2_N2236), .IN2(n7174), .QN(r843_n41) );
  NAND2X0 r843_U39 ( .IN1(r843_n40), .IN2(r843_n41), .QN(r843_n39) );
  NOR2X0 r843_U38 ( .QN(r843_n36), .IN1(r843_n38), .IN2(r843_n39) );
  AND2X1 r843_U37 ( .IN1(r843_n38), .IN2(r843_n39), .Q(r843_n37) );
  NOR2X0 r843_U36 ( .QN(P2_N2388), .IN1(r843_n36), .IN2(r843_n37) );
  OR2X1 r843_U34 ( .IN2(P2_N2237), .IN1(n7166), .Q(r843_n33) );
  NAND2X0 r843_U33 ( .IN1(P2_N2237), .IN2(n7166), .QN(r843_n34) );
  NAND2X0 r843_U32 ( .IN1(r843_n33), .IN2(r843_n34), .QN(r843_n32) );
  NOR2X0 r843_U31 ( .QN(r843_n29), .IN1(r843_n31), .IN2(r843_n32) );
  AND2X1 r843_U30 ( .IN1(r843_n31), .IN2(r843_n32), .Q(r843_n30) );
  NOR2X0 r843_U29 ( .QN(P2_N2389), .IN1(r843_n29), .IN2(r843_n30) );
  OR2X1 r843_U27 ( .IN2(P2_N2238), .IN1(n7164), .Q(r843_n26) );
  NAND2X0 r843_U26 ( .IN1(P2_N2238), .IN2(n7164), .QN(r843_n27) );
  NAND2X0 r843_U25 ( .IN1(r843_n26), .IN2(r843_n27), .QN(r843_n25) );
  NOR2X0 r843_U24 ( .QN(r843_n22), .IN1(r843_n24), .IN2(r843_n25) );
  AND2X1 r843_U23 ( .IN1(r843_n24), .IN2(r843_n25), .Q(r843_n23) );
  NOR2X0 r843_U22 ( .QN(P2_N2390), .IN1(r843_n22), .IN2(r843_n23) );
  OR2X1 r843_U20 ( .IN2(P2_N2239), .IN1(n7157), .Q(r843_n19) );
  NAND2X0 r843_U19 ( .IN1(P2_N2239), .IN2(n7157), .QN(r843_n20) );
  NAND2X0 r843_U18 ( .IN1(r843_n19), .IN2(r843_n20), .QN(r843_n18) );
  NOR2X0 r843_U17 ( .QN(r843_n15), .IN1(r843_n17), .IN2(r843_n18) );
  AND2X1 r843_U16 ( .IN1(r843_n17), .IN2(r843_n18), .Q(r843_n16) );
  NOR2X0 r843_U15 ( .QN(P2_N2391), .IN1(r843_n15), .IN2(r843_n16) );
  OR2X1 r843_U13 ( .IN2(P2_N2240), .IN1(n7153), .Q(r843_n12) );
  NAND2X0 r843_U12 ( .IN1(P2_N2240), .IN2(n7153), .QN(r843_n13) );
  NAND2X0 r843_U11 ( .IN1(r843_n12), .IN2(r843_n13), .QN(r843_n11) );
  NOR2X0 r843_U10 ( .QN(r843_n8), .IN1(r843_n10), .IN2(r843_n11) );
  AND2X1 r843_U9 ( .IN1(r843_n10), .IN2(r843_n11), .Q(r843_n9) );
  NOR2X0 r843_U8 ( .QN(P2_N2392), .IN1(r843_n8), .IN2(r843_n9) );
  OR2X1 r843_U6 ( .IN2(P2_N2241), .IN1(n7149), .Q(r843_n5) );
  NAND2X0 r843_U5 ( .IN1(P2_N2241), .IN2(n7149), .QN(r843_n6) );
  NAND2X0 r843_U4 ( .IN1(r843_n5), .IN2(r843_n6), .QN(r843_n4) );
  NOR2X0 r843_U3 ( .QN(r843_n1), .IN1(r843_n3), .IN2(r843_n4) );
  AND2X1 r843_U2 ( .IN1(r843_n3), .IN2(r843_n4), .Q(r843_n2) );
  NOR2X0 r843_U1 ( .QN(P2_N2393), .IN1(r843_n1), .IN2(r843_n2) );
  OR2X1 r843_U172 ( .IN2(P2_N2233), .IN1(n7184), .Q(r843_n162) );
  NAND2X0 r843_U171 ( .IN1(P2_N2233), .IN2(n7184), .QN(r843_n163) );
  NAND2X0 r843_U170 ( .IN1(r843_n162), .IN2(r843_n163), .QN(r843_n160) );
  NAND2X0 r843_U169 ( .IN1(r843_n160), .IN2(r843_n161), .QN(r843_n158) );
  OR2X1 r843_U168 ( .IN2(r843_n161), .IN1(r843_n160), .Q(r843_n159) );
  NAND2X0 r843_U167 ( .IN1(r843_n158), .IN2(r843_n159), .QN(P2_N2385) );
  NAND2X0 r843_U166 ( .IN1(n7263), .IN2(r843_n157), .QN(r843_n154) );
  OR2X1 r843_U165 ( .IN2(n7263), .IN1(r843_n157), .Q(r843_n156) );
  NAND2X0 r843_U164 ( .IN1(P2_N2251), .IN2(r843_n156), .QN(r843_n155) );
  NAND2X0 r843_U163 ( .IN1(r843_n154), .IN2(r843_n155), .QN(r843_n147) );
  OR2X1 r843_U161 ( .IN2(P2_N2252), .IN1(n7260), .Q(r843_n151) );
  NAND2X0 r843_U160 ( .IN1(P2_N2252), .IN2(n7260), .QN(r843_n152) );
  NAND2X0 r843_U159 ( .IN1(r843_n151), .IN2(r843_n152), .QN(r843_n150) );
  NOR2X0 r843_U158 ( .QN(r843_n148), .IN1(r843_n147), .IN2(r843_n150) );
  AND2X1 r843_U157 ( .IN1(r843_n147), .IN2(r843_n150), .Q(r843_n149) );
  NOR2X0 r843_U156 ( .QN(P2_N2404), .IN1(r843_n148), .IN2(r843_n149) );
  NAND2X0 r843_U155 ( .IN1(n7259), .IN2(r843_n147), .QN(r843_n144) );
  OR2X1 r843_U154 ( .IN2(n7259), .IN1(r843_n147), .Q(r843_n146) );
  NAND2X0 r843_U153 ( .IN1(P2_N2252), .IN2(r843_n146), .QN(r843_n145) );
  NAND2X0 r843_U152 ( .IN1(r843_n144), .IN2(r843_n145), .QN(r843_n137) );
  OR2X1 r843_U150 ( .IN2(P2_N2253), .IN1(n7253), .Q(r843_n141) );
  NAND2X0 r843_U149 ( .IN1(P2_N2253), .IN2(n7253), .QN(r843_n142) );
  NAND2X0 r843_U148 ( .IN1(r843_n141), .IN2(r843_n142), .QN(r843_n140) );
  NOR2X0 r843_U147 ( .QN(r843_n138), .IN1(r843_n137), .IN2(r843_n140) );
  AND2X1 r843_U146 ( .IN1(r843_n137), .IN2(r843_n140), .Q(r843_n139) );
  NOR2X0 r843_U145 ( .QN(P2_N2405), .IN1(r843_n138), .IN2(r843_n139) );
  NAND2X0 r843_U144 ( .IN1(n7252), .IN2(r843_n137), .QN(r843_n134) );
  OR2X1 r843_U143 ( .IN2(n7252), .IN1(r843_n137), .Q(r843_n136) );
  NAND2X0 r843_U142 ( .IN1(P2_N2253), .IN2(r843_n136), .QN(r843_n135) );
  NAND2X0 r843_U141 ( .IN1(r843_n134), .IN2(r843_n135), .QN(r843_n127) );
  OR2X1 r843_U139 ( .IN2(P2_N2254), .IN1(n7248), .Q(r843_n131) );
  NAND2X0 r843_U138 ( .IN1(P2_N2254), .IN2(n7248), .QN(r843_n132) );
  NAND2X0 r843_U137 ( .IN1(r843_n131), .IN2(r843_n132), .QN(r843_n130) );
  NOR2X0 r843_U136 ( .QN(r843_n128), .IN1(r843_n127), .IN2(r843_n130) );
  AND2X1 r843_U135 ( .IN1(r843_n127), .IN2(r843_n130), .Q(r843_n129) );
  NOR2X0 r843_U134 ( .QN(P2_N2406), .IN1(r843_n128), .IN2(r843_n129) );
  NAND2X0 r843_U133 ( .IN1(P2_N5093), .IN2(r843_n127), .QN(r843_n124) );
  OR2X1 r843_U132 ( .IN2(P2_N5093), .IN1(r843_n127), .Q(r843_n126) );
  NAND2X0 r843_U131 ( .IN1(P2_N2254), .IN2(r843_n126), .QN(r843_n125) );
  NAND2X0 r843_U130 ( .IN1(r843_n124), .IN2(r843_n125), .QN(r843_n117) );
  OR2X1 r843_U128 ( .IN2(P2_N2255), .IN1(n7243), .Q(r843_n121) );
  NAND2X0 r843_U127 ( .IN1(P2_N2255), .IN2(n7243), .QN(r843_n122) );
  NAND2X0 r843_U126 ( .IN1(r843_n121), .IN2(r843_n122), .QN(r843_n120) );
  NOR2X0 r843_U125 ( .QN(r843_n118), .IN1(r843_n117), .IN2(r843_n120) );
  AND2X1 r843_U124 ( .IN1(r843_n117), .IN2(r843_n120), .Q(r843_n119) );
  NOR2X0 r843_U123 ( .QN(P2_N2407), .IN1(r843_n118), .IN2(r843_n119) );
  NAND2X0 r843_U122 ( .IN1(n7242), .IN2(r843_n117), .QN(r843_n114) );
  OR2X1 r843_U121 ( .IN2(n7242), .IN1(r843_n117), .Q(r843_n116) );
  NAND2X0 r843_U120 ( .IN1(P2_N2255), .IN2(r843_n116), .QN(r843_n115) );
  NAND2X0 r843_U119 ( .IN1(r843_n114), .IN2(r843_n115), .QN(r843_n107) );
  OR2X1 r843_U117 ( .IN2(P2_N2256), .IN1(n7239), .Q(r843_n111) );
  NAND2X0 r843_U116 ( .IN1(P2_N2256), .IN2(n7239), .QN(r843_n112) );
  NAND2X0 r843_U115 ( .IN1(r843_n111), .IN2(r843_n112), .QN(r843_n110) );
  NOR2X0 r843_U114 ( .QN(r843_n108), .IN1(r843_n107), .IN2(r843_n110) );
  AND2X1 r843_U113 ( .IN1(r843_n107), .IN2(r843_n110), .Q(r843_n109) );
  NOR2X0 r843_U112 ( .QN(P2_N2408), .IN1(r843_n108), .IN2(r843_n109) );
  NAND2X0 r843_U111 ( .IN1(n7238), .IN2(r843_n107), .QN(r843_n104) );
  OR2X1 r843_U110 ( .IN2(n7238), .IN1(r843_n107), .Q(r843_n106) );
  NAND2X0 r843_U109 ( .IN1(P2_N2256), .IN2(r843_n106), .QN(r843_n105) );
  NAND2X0 r843_U108 ( .IN1(r843_n104), .IN2(r843_n105), .QN(r843_n97) );
  OR2X1 r843_U106 ( .IN2(P2_N2257), .IN1(n7234), .Q(r843_n101) );
  NAND2X0 r843_U105 ( .IN1(P2_N2257), .IN2(n7234), .QN(r843_n102) );
  NAND2X0 r843_U104 ( .IN1(r843_n101), .IN2(r843_n102), .QN(r843_n100) );
  NOR2X0 r843_U103 ( .QN(r843_n98), .IN1(r843_n97), .IN2(r843_n100) );
  AND2X1 r843_U102 ( .IN1(r843_n97), .IN2(r843_n100), .Q(r843_n99) );
  NOR2X0 r843_U101 ( .QN(P2_N2409), .IN1(r843_n98), .IN2(r843_n99) );
  NAND2X0 r843_U100 ( .IN1(P2_N5096), .IN2(r843_n97), .QN(r843_n94) );
  OR2X1 r843_U99 ( .IN2(P2_N5096), .IN1(r843_n97), .Q(r843_n96) );
  NAND2X0 r843_U98 ( .IN1(P2_N2257), .IN2(r843_n96), .QN(r843_n95) );
  NAND2X0 r843_U97 ( .IN1(r843_n94), .IN2(r843_n95), .QN(r843_n87) );
  OR2X1 r843_U95 ( .IN2(P2_N2258), .IN1(n7229), .Q(r843_n91) );
  NAND2X0 r843_U94 ( .IN1(P2_N2258), .IN2(n7229), .QN(r843_n92) );
  NAND2X0 r843_U93 ( .IN1(r843_n91), .IN2(r843_n92), .QN(r843_n90) );
  NOR2X0 r843_U92 ( .QN(r843_n88), .IN1(r843_n87), .IN2(r843_n90) );
  AND2X1 r843_U91 ( .IN1(r843_n87), .IN2(r843_n90), .Q(r843_n89) );
  NOR2X0 r843_U90 ( .QN(P2_N2410), .IN1(r843_n88), .IN2(r843_n89) );
  NAND2X0 r843_U89 ( .IN1(P2_N5097), .IN2(r843_n87), .QN(r843_n84) );
  OR2X1 r843_U88 ( .IN2(P2_N5097), .IN1(r843_n87), .Q(r843_n86) );
  NAND2X0 r843_U87 ( .IN1(P2_N2258), .IN2(r843_n86), .QN(r843_n85) );
  NAND2X0 r843_U86 ( .IN1(r843_n84), .IN2(r843_n85), .QN(r843_n77) );
  OR2X1 r843_U84 ( .IN2(P2_N2259), .IN1(n7224), .Q(r843_n81) );
  NAND2X0 r843_U83 ( .IN1(P2_N2259), .IN2(n7224), .QN(r843_n82) );
  NAND2X0 r843_U82 ( .IN1(r843_n81), .IN2(r843_n82), .QN(r843_n80) );
  NOR2X0 r843_U81 ( .QN(r843_n78), .IN1(r843_n77), .IN2(r843_n80) );
  AND2X1 r843_U80 ( .IN1(r843_n77), .IN2(r843_n80), .Q(r843_n79) );
  NAND2X0 r843_U265 ( .IN1(P2_N2243), .IN2(n7214), .QN(r843_n249) );
  NAND2X0 r843_U264 ( .IN1(r843_n248), .IN2(r843_n249), .QN(r843_n247) );
  NOR2X0 r843_U263 ( .QN(r843_n245), .IN1(r843_n244), .IN2(r843_n247) );
  AND2X1 r843_U262 ( .IN1(r843_n244), .IN2(r843_n247), .Q(r843_n246) );
  NOR2X0 r843_U261 ( .QN(P2_N2395), .IN1(r843_n245), .IN2(r843_n246) );
  NAND2X0 r843_U260 ( .IN1(n7216), .IN2(r843_n244), .QN(r843_n241) );
  OR2X1 r843_U259 ( .IN2(n7216), .IN1(r843_n244), .Q(r843_n243) );
  NAND2X0 r843_U258 ( .IN1(P2_N2243), .IN2(r843_n243), .QN(r843_n242) );
  NAND2X0 r843_U257 ( .IN1(r843_n241), .IN2(r843_n242), .QN(r843_n234) );
  OR2X1 r843_U255 ( .IN2(P2_N2244), .IN1(n7211), .Q(r843_n238) );
  NAND2X0 r843_U254 ( .IN1(P2_N2244), .IN2(n7211), .QN(r843_n239) );
  NAND2X0 r843_U253 ( .IN1(r843_n238), .IN2(r843_n239), .QN(r843_n237) );
  NOR2X0 r843_U252 ( .QN(r843_n235), .IN1(r843_n234), .IN2(r843_n237) );
  AND2X1 r843_U251 ( .IN1(r843_n234), .IN2(r843_n237), .Q(r843_n236) );
  NOR2X0 r843_U250 ( .QN(P2_N2396), .IN1(r843_n235), .IN2(r843_n236) );
  NAND2X0 r843_U249 ( .IN1(n7210), .IN2(r843_n234), .QN(r843_n231) );
  OR2X1 r843_U248 ( .IN2(n7210), .IN1(r843_n234), .Q(r843_n233) );
  NAND2X0 r843_U247 ( .IN1(P2_N2244), .IN2(r843_n233), .QN(r843_n232) );
  NAND2X0 r843_U246 ( .IN1(r843_n231), .IN2(r843_n232), .QN(r843_n224) );
  OR2X1 r843_U244 ( .IN2(P2_N2245), .IN1(n7208), .Q(r843_n228) );
  NAND2X0 r843_U243 ( .IN1(P2_N2245), .IN2(n7208), .QN(r843_n229) );
  NAND2X0 r843_U242 ( .IN1(r843_n228), .IN2(r843_n229), .QN(r843_n227) );
  NOR2X0 r843_U241 ( .QN(r843_n225), .IN1(r843_n224), .IN2(r843_n227) );
  AND2X1 r843_U240 ( .IN1(r843_n224), .IN2(r843_n227), .Q(r843_n226) );
  NOR2X0 r843_U239 ( .QN(P2_N2397), .IN1(r843_n225), .IN2(r843_n226) );
  NAND2X0 r843_U238 ( .IN1(P2_N5084), .IN2(r843_n224), .QN(r843_n221) );
  OR2X1 r843_U237 ( .IN2(P2_N5084), .IN1(r843_n224), .Q(r843_n223) );
  NAND2X0 r843_U236 ( .IN1(P2_N2245), .IN2(r843_n223), .QN(r843_n222) );
  NAND2X0 r843_U235 ( .IN1(r843_n221), .IN2(r843_n222), .QN(r843_n214) );
  OR2X1 r843_U233 ( .IN2(P2_N2246), .IN1(n7205), .Q(r843_n218) );
  NAND2X0 r843_U232 ( .IN1(P2_N2246), .IN2(n7205), .QN(r843_n219) );
  NAND2X0 r843_U231 ( .IN1(r843_n218), .IN2(r843_n219), .QN(r843_n217) );
  NOR2X0 r843_U230 ( .QN(r843_n215), .IN1(r843_n214), .IN2(r843_n217) );
  AND2X1 r843_U229 ( .IN1(r843_n214), .IN2(r843_n217), .Q(r843_n216) );
  NOR2X0 r843_U228 ( .QN(P2_N2398), .IN1(r843_n215), .IN2(r843_n216) );
  NAND2X0 r843_U227 ( .IN1(P2_N5085), .IN2(r843_n214), .QN(r843_n211) );
  OR2X1 r843_U226 ( .IN2(P2_N5085), .IN1(r843_n214), .Q(r843_n213) );
  NAND2X0 r843_U225 ( .IN1(P2_N2246), .IN2(r843_n213), .QN(r843_n212) );
  NAND2X0 r843_U224 ( .IN1(r843_n211), .IN2(r843_n212), .QN(r843_n204) );
  OR2X1 r843_U222 ( .IN2(P2_N2247), .IN1(n7201), .Q(r843_n208) );
  NAND2X0 r843_U221 ( .IN1(P2_N2247), .IN2(n7201), .QN(r843_n209) );
  NAND2X0 r843_U220 ( .IN1(r843_n208), .IN2(r843_n209), .QN(r843_n207) );
  NOR2X0 r843_U219 ( .QN(r843_n205), .IN1(r843_n204), .IN2(r843_n207) );
  AND2X1 r843_U218 ( .IN1(r843_n204), .IN2(r843_n207), .Q(r843_n206) );
  NOR2X0 r843_U217 ( .QN(P2_N2399), .IN1(r843_n205), .IN2(r843_n206) );
  NAND2X0 r843_U216 ( .IN1(P2_N5086), .IN2(r843_n204), .QN(r843_n201) );
  OR2X1 r843_U215 ( .IN2(P2_N5086), .IN1(r843_n204), .Q(r843_n203) );
  NAND2X0 r843_U214 ( .IN1(P2_N2247), .IN2(r843_n203), .QN(r843_n202) );
  NAND2X0 r843_U213 ( .IN1(r843_n201), .IN2(r843_n202), .QN(r843_n194) );
  OR2X1 r843_U211 ( .IN2(P2_N2248), .IN1(n7197), .Q(r843_n198) );
  NAND2X0 r843_U210 ( .IN1(P2_N2248), .IN2(n7197), .QN(r843_n199) );
  NAND2X0 r843_U209 ( .IN1(r843_n198), .IN2(r843_n199), .QN(r843_n197) );
  NOR2X0 r843_U208 ( .QN(r843_n195), .IN1(r843_n194), .IN2(r843_n197) );
  AND2X1 r843_U207 ( .IN1(r843_n194), .IN2(r843_n197), .Q(r843_n196) );
  NOR2X0 r843_U206 ( .QN(P2_N2400), .IN1(r843_n195), .IN2(r843_n196) );
  NAND2X0 r843_U205 ( .IN1(P2_N5087), .IN2(r843_n194), .QN(r843_n191) );
  OR2X1 r843_U204 ( .IN2(P2_N5087), .IN1(r843_n194), .Q(r843_n193) );
  NAND2X0 r843_U203 ( .IN1(P2_N2248), .IN2(r843_n193), .QN(r843_n192) );
  NAND2X0 r843_U202 ( .IN1(r843_n191), .IN2(r843_n192), .QN(r843_n184) );
  OR2X1 r843_U200 ( .IN2(P2_N2249), .IN1(n7195), .Q(r843_n188) );
  NAND2X0 r843_U199 ( .IN1(P2_N2249), .IN2(n7195), .QN(r843_n189) );
  NAND2X0 r843_U198 ( .IN1(r843_n188), .IN2(r843_n189), .QN(r843_n187) );
  NOR2X0 r843_U197 ( .QN(r843_n185), .IN1(r843_n184), .IN2(r843_n187) );
  AND2X1 r843_U196 ( .IN1(r843_n184), .IN2(r843_n187), .Q(r843_n186) );
  NOR2X0 r843_U195 ( .QN(P2_N2401), .IN1(r843_n185), .IN2(r843_n186) );
  NAND2X0 r843_U194 ( .IN1(P2_N5088), .IN2(r843_n184), .QN(r843_n181) );
  OR2X1 r843_U193 ( .IN2(P2_N5088), .IN1(r843_n184), .Q(r843_n183) );
  NAND2X0 r843_U192 ( .IN1(P2_N2249), .IN2(r843_n183), .QN(r843_n182) );
  NAND2X0 r843_U191 ( .IN1(r843_n181), .IN2(r843_n182), .QN(r843_n174) );
  OR2X1 r843_U189 ( .IN2(P2_N2250), .IN1(n7188), .Q(r843_n178) );
  NAND2X0 r843_U188 ( .IN1(P2_N2250), .IN2(n7188), .QN(r843_n179) );
  NAND2X0 r843_U187 ( .IN1(r843_n178), .IN2(r843_n179), .QN(r843_n177) );
  NOR2X0 r843_U186 ( .QN(r843_n175), .IN1(r843_n174), .IN2(r843_n177) );
  AND2X1 r843_U185 ( .IN1(r843_n174), .IN2(r843_n177), .Q(r843_n176) );
  NOR2X0 r843_U184 ( .QN(P2_N2402), .IN1(r843_n175), .IN2(r843_n176) );
  NAND2X0 r843_U183 ( .IN1(P2_N5089), .IN2(r843_n174), .QN(r843_n171) );
  OR2X1 r843_U182 ( .IN2(P2_N5089), .IN1(r843_n174), .Q(r843_n173) );
  NAND2X0 r843_U181 ( .IN1(P2_N2250), .IN2(r843_n173), .QN(r843_n172) );
  NAND2X0 r843_U180 ( .IN1(r843_n171), .IN2(r843_n172), .QN(r843_n157) );
  OR2X1 r843_U178 ( .IN2(P2_N2251), .IN1(n7264), .Q(r843_n168) );
  NAND2X0 r843_U177 ( .IN1(P2_N2251), .IN2(n7264), .QN(r843_n169) );
  NAND2X0 r843_U176 ( .IN1(r843_n168), .IN2(r843_n169), .QN(r843_n167) );
  NOR2X0 r843_U175 ( .QN(r843_n165), .IN1(r843_n157), .IN2(r843_n167) );
  AND2X1 r843_U174 ( .IN1(r843_n157), .IN2(r843_n167), .Q(r843_n166) );
  NOR2X0 r843_U173 ( .QN(P2_N2403), .IN1(r843_n165), .IN2(r843_n166) );
  OR2X1 r843_U319 ( .IN2(P2_N2232), .IN1(n2919), .Q(r843_n288) );
  NAND2X0 r843_U318 ( .IN1(P2_N2232), .IN2(n2919), .QN(r843_n289) );
  NAND2X0 r843_U317 ( .IN1(r843_n288), .IN2(r843_n289), .QN(P2_N2384) );
  NAND2X0 r843_U315 ( .IN1(P2_N2232), .IN2(n7035), .QN(r843_n161) );
  OR2X1 r843_U314 ( .IN2(r843_n161), .IN1(n7184), .Q(r843_n285) );
  NAND2X0 r843_U313 ( .IN1(n7184), .IN2(r843_n161), .QN(r843_n287) );
  NAND2X0 r843_U312 ( .IN1(P2_N2233), .IN2(r843_n287), .QN(r843_n286) );
  NAND2X0 r843_U311 ( .IN1(r843_n285), .IN2(r843_n286), .QN(r843_n52) );
  NAND2X0 r843_U310 ( .IN1(P2_N5073), .IN2(r843_n52), .QN(r843_n282) );
  OR2X1 r843_U309 ( .IN2(P2_N5073), .IN1(r843_n52), .Q(r843_n284) );
  NAND2X0 r843_U308 ( .IN1(P2_N2234), .IN2(r843_n284), .QN(r843_n283) );
  NAND2X0 r843_U307 ( .IN1(r843_n282), .IN2(r843_n283), .QN(r843_n45) );
  NAND2X0 r843_U306 ( .IN1(P2_N5074), .IN2(r843_n45), .QN(r843_n279) );
  OR2X1 r843_U305 ( .IN2(P2_N5074), .IN1(r843_n45), .Q(r843_n281) );
  NAND2X0 r843_U304 ( .IN1(P2_N2235), .IN2(r843_n281), .QN(r843_n280) );
  NAND2X0 r843_U303 ( .IN1(r843_n279), .IN2(r843_n280), .QN(r843_n38) );
  NAND2X0 r843_U302 ( .IN1(P2_N5075), .IN2(r843_n38), .QN(r843_n276) );
  OR2X1 r843_U301 ( .IN2(P2_N5075), .IN1(r843_n38), .Q(r843_n278) );
  NAND2X0 r843_U300 ( .IN1(P2_N2236), .IN2(r843_n278), .QN(r843_n277) );
  NAND2X0 r843_U299 ( .IN1(r843_n276), .IN2(r843_n277), .QN(r843_n31) );
  NAND2X0 r843_U298 ( .IN1(P2_N5076), .IN2(r843_n31), .QN(r843_n273) );
  OR2X1 r843_U297 ( .IN2(P2_N5076), .IN1(r843_n31), .Q(r843_n275) );
  NAND2X0 r843_U296 ( .IN1(P2_N2237), .IN2(r843_n275), .QN(r843_n274) );
  NAND2X0 r843_U295 ( .IN1(r843_n273), .IN2(r843_n274), .QN(r843_n24) );
  NAND2X0 r843_U294 ( .IN1(n7162), .IN2(r843_n24), .QN(r843_n270) );
  OR2X1 r843_U293 ( .IN2(n7162), .IN1(r843_n24), .Q(r843_n272) );
  NAND2X0 r843_U292 ( .IN1(P2_N2238), .IN2(r843_n272), .QN(r843_n271) );
  NAND2X0 r843_U291 ( .IN1(r843_n270), .IN2(r843_n271), .QN(r843_n17) );
  NAND2X0 r843_U290 ( .IN1(P2_N5078), .IN2(r843_n17), .QN(r843_n267) );
  OR2X1 r843_U289 ( .IN2(P2_N5078), .IN1(r843_n17), .Q(r843_n269) );
  NAND2X0 r843_U288 ( .IN1(P2_N2239), .IN2(r843_n269), .QN(r843_n268) );
  NAND2X0 r843_U287 ( .IN1(r843_n267), .IN2(r843_n268), .QN(r843_n10) );
  NAND2X0 r843_U286 ( .IN1(n7154), .IN2(r843_n10), .QN(r843_n264) );
  OR2X1 r843_U285 ( .IN2(n7154), .IN1(r843_n10), .Q(r843_n266) );
  NAND2X0 r843_U284 ( .IN1(P2_N2240), .IN2(r843_n266), .QN(r843_n265) );
  NAND2X0 r843_U283 ( .IN1(r843_n264), .IN2(r843_n265), .QN(r843_n3) );
  NAND2X0 r843_U282 ( .IN1(n7151), .IN2(r843_n3), .QN(r843_n261) );
  OR2X1 r843_U281 ( .IN2(n7151), .IN1(r843_n3), .Q(r843_n263) );
  NAND2X0 r843_U280 ( .IN1(P2_N2241), .IN2(r843_n263), .QN(r843_n262) );
  NAND2X0 r843_U279 ( .IN1(r843_n261), .IN2(r843_n262), .QN(r843_n254) );
  OR2X1 r843_U277 ( .IN2(P2_N2242), .IN1(n7219), .Q(r843_n258) );
  NAND2X0 r843_U276 ( .IN1(P2_N2242), .IN2(n7219), .QN(r843_n259) );
  NAND2X0 r843_U275 ( .IN1(r843_n258), .IN2(r843_n259), .QN(r843_n257) );
  NOR2X0 r843_U274 ( .QN(r843_n255), .IN1(r843_n254), .IN2(r843_n257) );
  AND2X1 r843_U273 ( .IN1(r843_n254), .IN2(r843_n257), .Q(r843_n256) );
  NOR2X0 r843_U272 ( .QN(P2_N2394), .IN1(r843_n255), .IN2(r843_n256) );
  NAND2X0 r843_U271 ( .IN1(P2_N5081), .IN2(r843_n254), .QN(r843_n251) );
  OR2X1 r843_U270 ( .IN2(P2_N5081), .IN1(r843_n254), .Q(r843_n253) );
  NAND2X0 r843_U269 ( .IN1(P2_N2242), .IN2(r843_n253), .QN(r843_n252) );
  NAND2X0 r843_U268 ( .IN1(r843_n251), .IN2(r843_n252), .QN(r843_n244) );
  OR2X1 r843_U266 ( .IN2(P2_N2243), .IN1(n7214), .Q(r843_n248) );
  OR2X1 r800_U5 ( .IN2(n7070), .IN1(r800_n7), .Q(r800_n6) );
  NAND2X0 r800_U4 ( .IN1(r800_n5), .IN2(r800_n6), .QN(r800_n3) );
  NAND2X0 r800_U3 ( .IN1(r800_n3), .IN2(r800_n4), .QN(r800_n1) );
  OR2X1 r800_U2 ( .IN2(r800_n4), .IN1(r800_n3), .Q(r800_n2) );
  NAND2X0 r800_U1 ( .IN1(r800_n1), .IN2(r800_n2), .QN(P1_N2519) );
  OR2X1 r800_U98 ( .IN2(n7138), .IN1(r800_n106), .Q(r800_n104) );
  NAND2X0 r800_U97 ( .IN1(r800_n104), .IN2(r800_n105), .QN(r800_n103) );
  NAND2X0 r800_U96 ( .IN1(r800_n102), .IN2(r800_n103), .QN(r800_n96) );
  NAND2X0 r800_U95 ( .IN1(r800_n101), .IN2(r800_n96), .QN(r800_n99) );
  OR2X1 r800_U94 ( .IN2(r800_n96), .IN1(r800_n101), .Q(r800_n100) );
  NAND2X0 r800_U93 ( .IN1(r800_n99), .IN2(r800_n100), .QN(P1_N2535) );
  INVX0 r800_U92 ( .ZN(r800_n85), .INP(P1_N2384) );
  NAND2X0 r800_U91 ( .IN1(n7124), .IN2(r800_n85), .QN(r800_n97) );
  OR2X1 r800_U90 ( .IN2(n7124), .IN1(r800_n85), .Q(r800_n98) );
  NAND2X0 r800_U89 ( .IN1(r800_n97), .IN2(r800_n98), .QN(r800_n91) );
  NAND2X0 r800_U88 ( .IN1(P1_N5174), .IN2(r800_n96), .QN(r800_n92) );
  OR2X1 r800_U87 ( .IN2(P1_N5174), .IN1(r800_n96), .Q(r800_n94) );
  NAND2X0 r800_U86 ( .IN1(r800_n94), .IN2(r800_n95), .QN(r800_n93) );
  NAND2X0 r800_U85 ( .IN1(r800_n92), .IN2(r800_n93), .QN(r800_n86) );
  NAND2X0 r800_U84 ( .IN1(r800_n91), .IN2(r800_n86), .QN(r800_n89) );
  OR2X1 r800_U83 ( .IN2(r800_n86), .IN1(r800_n91), .Q(r800_n90) );
  NAND2X0 r800_U82 ( .IN1(r800_n89), .IN2(r800_n90), .QN(P1_N2536) );
  INVX0 r800_U81 ( .ZN(r800_n75), .INP(P1_N2385) );
  NAND2X0 r800_U80 ( .IN1(P1_N5176), .IN2(r800_n75), .QN(r800_n87) );
  OR2X1 r800_U79 ( .IN2(P1_N5176), .IN1(r800_n75), .Q(r800_n88) );
  NAND2X0 r800_U78 ( .IN1(r800_n87), .IN2(r800_n88), .QN(r800_n81) );
  NAND2X0 r800_U77 ( .IN1(n7124), .IN2(r800_n86), .QN(r800_n82) );
  OR2X1 r800_U76 ( .IN2(n7124), .IN1(r800_n86), .Q(r800_n84) );
  NAND2X0 r800_U75 ( .IN1(r800_n84), .IN2(r800_n85), .QN(r800_n83) );
  NAND2X0 r800_U74 ( .IN1(r800_n82), .IN2(r800_n83), .QN(r800_n76) );
  NAND2X0 r800_U73 ( .IN1(r800_n81), .IN2(r800_n76), .QN(r800_n79) );
  OR2X1 r800_U72 ( .IN2(r800_n76), .IN1(r800_n81), .Q(r800_n80) );
  NAND2X0 r800_U71 ( .IN1(r800_n79), .IN2(r800_n80), .QN(P1_N2537) );
  INVX0 r800_U70 ( .ZN(r800_n64), .INP(P1_N2386) );
  NAND2X0 r800_U69 ( .IN1(P1_N5177), .IN2(r800_n64), .QN(r800_n77) );
  OR2X1 r800_U68 ( .IN2(P1_N5177), .IN1(r800_n64), .Q(r800_n78) );
  NAND2X0 r800_U67 ( .IN1(r800_n77), .IN2(r800_n78), .QN(r800_n71) );
  NAND2X0 r800_U66 ( .IN1(n7122), .IN2(r800_n76), .QN(r800_n72) );
  OR2X1 r800_U65 ( .IN2(P1_N5176), .IN1(r800_n76), .Q(r800_n74) );
  NAND2X0 r800_U64 ( .IN1(r800_n74), .IN2(r800_n75), .QN(r800_n73) );
  NAND2X0 r800_U63 ( .IN1(r800_n72), .IN2(r800_n73), .QN(r800_n65) );
  NAND2X0 r800_U62 ( .IN1(r800_n71), .IN2(r800_n65), .QN(r800_n69) );
  OR2X1 r800_U61 ( .IN2(r800_n65), .IN1(r800_n71), .Q(r800_n70) );
  NAND2X0 r800_U60 ( .IN1(r800_n69), .IN2(r800_n70), .QN(P1_N2538) );
  OR2X1 r800_U58 ( .IN2(P1_N2387), .IN1(n7146), .Q(r800_n66) );
  NAND2X0 r800_U57 ( .IN1(P1_N2387), .IN2(n7146), .QN(r800_n67) );
  NAND2X0 r800_U56 ( .IN1(r800_n66), .IN2(r800_n67), .QN(r800_n60) );
  NAND2X0 r800_U55 ( .IN1(P1_N5177), .IN2(r800_n65), .QN(r800_n61) );
  OR2X1 r800_U54 ( .IN2(P1_N5177), .IN1(r800_n65), .Q(r800_n63) );
  NAND2X0 r800_U53 ( .IN1(r800_n63), .IN2(r800_n64), .QN(r800_n62) );
  NAND2X0 r800_U52 ( .IN1(r800_n61), .IN2(r800_n62), .QN(r800_n59) );
  NAND2X0 r800_U51 ( .IN1(r800_n60), .IN2(r800_n59), .QN(r800_n57) );
  OR2X1 r800_U50 ( .IN2(r800_n60), .IN1(r800_n59), .Q(r800_n58) );
  NAND2X0 r800_U49 ( .IN1(r800_n57), .IN2(r800_n58), .QN(P1_N2539) );
  NAND2X0 r800_U48 ( .IN1(P1_N5151), .IN2(r800_n56), .QN(r800_n54) );
  OR2X1 r800_U47 ( .IN2(P1_N5151), .IN1(r800_n56), .Q(r800_n55) );
  NAND2X0 r800_U46 ( .IN1(r800_n54), .IN2(r800_n55), .QN(r800_n52) );
  NAND2X0 r800_U45 ( .IN1(r800_n52), .IN2(r800_n53), .QN(r800_n50) );
  OR2X1 r800_U44 ( .IN2(r800_n53), .IN1(r800_n52), .Q(r800_n51) );
  NAND2X0 r800_U43 ( .IN1(r800_n50), .IN2(r800_n51), .QN(P1_N2512) );
  NAND2X0 r800_U42 ( .IN1(P1_N5152), .IN2(r800_n49), .QN(r800_n47) );
  OR2X1 r800_U41 ( .IN2(P1_N5152), .IN1(r800_n49), .Q(r800_n48) );
  NAND2X0 r800_U40 ( .IN1(r800_n47), .IN2(r800_n48), .QN(r800_n45) );
  NAND2X0 r800_U39 ( .IN1(r800_n45), .IN2(r800_n46), .QN(r800_n43) );
  OR2X1 r800_U38 ( .IN2(r800_n46), .IN1(r800_n45), .Q(r800_n44) );
  NAND2X0 r800_U37 ( .IN1(r800_n43), .IN2(r800_n44), .QN(P1_N2513) );
  NAND2X0 r800_U36 ( .IN1(P1_N5153), .IN2(r800_n42), .QN(r800_n40) );
  OR2X1 r800_U35 ( .IN2(P1_N5153), .IN1(r800_n42), .Q(r800_n41) );
  NAND2X0 r800_U34 ( .IN1(r800_n40), .IN2(r800_n41), .QN(r800_n38) );
  NAND2X0 r800_U33 ( .IN1(r800_n38), .IN2(r800_n39), .QN(r800_n36) );
  OR2X1 r800_U32 ( .IN2(r800_n39), .IN1(r800_n38), .Q(r800_n37) );
  NAND2X0 r800_U31 ( .IN1(r800_n36), .IN2(r800_n37), .QN(P1_N2514) );
  NAND2X0 r800_U30 ( .IN1(P1_N5154), .IN2(r800_n35), .QN(r800_n33) );
  OR2X1 r800_U29 ( .IN2(P1_N5154), .IN1(r800_n35), .Q(r800_n34) );
  NAND2X0 r800_U28 ( .IN1(r800_n33), .IN2(r800_n34), .QN(r800_n31) );
  NAND2X0 r800_U27 ( .IN1(r800_n31), .IN2(r800_n32), .QN(r800_n29) );
  OR2X1 r800_U26 ( .IN2(r800_n32), .IN1(r800_n31), .Q(r800_n30) );
  NAND2X0 r800_U25 ( .IN1(r800_n29), .IN2(r800_n30), .QN(P1_N2515) );
  NAND2X0 r800_U24 ( .IN1(n7080), .IN2(r800_n28), .QN(r800_n26) );
  OR2X1 r800_U23 ( .IN2(n7080), .IN1(r800_n28), .Q(r800_n27) );
  NAND2X0 r800_U22 ( .IN1(r800_n26), .IN2(r800_n27), .QN(r800_n24) );
  NAND2X0 r800_U21 ( .IN1(r800_n24), .IN2(r800_n25), .QN(r800_n22) );
  OR2X1 r800_U20 ( .IN2(r800_n25), .IN1(r800_n24), .Q(r800_n23) );
  NAND2X0 r800_U19 ( .IN1(r800_n22), .IN2(r800_n23), .QN(P1_N2516) );
  NAND2X0 r800_U18 ( .IN1(n7075), .IN2(r800_n21), .QN(r800_n19) );
  OR2X1 r800_U17 ( .IN2(n7075), .IN1(r800_n21), .Q(r800_n20) );
  NAND2X0 r800_U16 ( .IN1(r800_n19), .IN2(r800_n20), .QN(r800_n17) );
  NAND2X0 r800_U15 ( .IN1(r800_n17), .IN2(r800_n18), .QN(r800_n15) );
  OR2X1 r800_U14 ( .IN2(r800_n18), .IN1(r800_n17), .Q(r800_n16) );
  NAND2X0 r800_U13 ( .IN1(r800_n15), .IN2(r800_n16), .QN(P1_N2517) );
  NAND2X0 r800_U12 ( .IN1(n7072), .IN2(r800_n14), .QN(r800_n12) );
  OR2X1 r800_U11 ( .IN2(n7072), .IN1(r800_n14), .Q(r800_n13) );
  NAND2X0 r800_U10 ( .IN1(r800_n12), .IN2(r800_n13), .QN(r800_n10) );
  NAND2X0 r800_U9 ( .IN1(r800_n10), .IN2(r800_n11), .QN(r800_n8) );
  OR2X1 r800_U8 ( .IN2(r800_n11), .IN1(r800_n10), .Q(r800_n9) );
  NAND2X0 r800_U7 ( .IN1(r800_n8), .IN2(r800_n9), .QN(P1_N2518) );
  NAND2X0 r800_U6 ( .IN1(n7070), .IN2(r800_n7), .QN(r800_n5) );
  NAND2X0 r800_U191 ( .IN1(r800_n192), .IN2(r800_n193), .QN(r800_n191) );
  NAND2X0 r800_U190 ( .IN1(r800_n190), .IN2(r800_n191), .QN(r800_n184) );
  NAND2X0 r800_U189 ( .IN1(r800_n189), .IN2(r800_n184), .QN(r800_n187) );
  OR2X1 r800_U188 ( .IN2(r800_n184), .IN1(r800_n189), .Q(r800_n188) );
  NAND2X0 r800_U187 ( .IN1(r800_n187), .IN2(r800_n188), .QN(P1_N2527) );
  INVX0 r800_U186 ( .ZN(r800_n173), .INP(P1_N2376) );
  NAND2X0 r800_U185 ( .IN1(P1_N5167), .IN2(r800_n173), .QN(r800_n185) );
  OR2X1 r800_U184 ( .IN2(P1_N5167), .IN1(r800_n173), .Q(r800_n186) );
  NAND2X0 r800_U183 ( .IN1(r800_n185), .IN2(r800_n186), .QN(r800_n179) );
  NAND2X0 r800_U182 ( .IN1(n7106), .IN2(r800_n184), .QN(r800_n180) );
  OR2X1 r800_U181 ( .IN2(n7106), .IN1(r800_n184), .Q(r800_n182) );
  NAND2X0 r800_U180 ( .IN1(r800_n182), .IN2(r800_n183), .QN(r800_n181) );
  NAND2X0 r800_U179 ( .IN1(r800_n180), .IN2(r800_n181), .QN(r800_n174) );
  NAND2X0 r800_U178 ( .IN1(r800_n179), .IN2(r800_n174), .QN(r800_n177) );
  OR2X1 r800_U177 ( .IN2(r800_n174), .IN1(r800_n179), .Q(r800_n178) );
  NAND2X0 r800_U176 ( .IN1(r800_n177), .IN2(r800_n178), .QN(P1_N2528) );
  INVX0 r800_U175 ( .ZN(r800_n155), .INP(P1_N2377) );
  NAND2X0 r800_U174 ( .IN1(n7099), .IN2(r800_n155), .QN(r800_n175) );
  OR2X1 r800_U173 ( .IN2(n7099), .IN1(r800_n155), .Q(r800_n176) );
  NAND2X0 r800_U172 ( .IN1(r800_n175), .IN2(r800_n176), .QN(r800_n169) );
  NAND2X0 r800_U171 ( .IN1(P1_N5167), .IN2(r800_n174), .QN(r800_n170) );
  OR2X1 r800_U170 ( .IN2(P1_N5167), .IN1(r800_n174), .Q(r800_n172) );
  NAND2X0 r800_U169 ( .IN1(r800_n172), .IN2(r800_n173), .QN(r800_n171) );
  NAND2X0 r800_U168 ( .IN1(r800_n170), .IN2(r800_n171), .QN(r800_n156) );
  NAND2X0 r800_U167 ( .IN1(r800_n169), .IN2(r800_n156), .QN(r800_n167) );
  OR2X1 r800_U166 ( .IN2(r800_n156), .IN1(r800_n169), .Q(r800_n168) );
  NAND2X0 r800_U165 ( .IN1(r800_n167), .IN2(r800_n168), .QN(P1_N2529) );
  NAND2X0 r800_U164 ( .IN1(P1_N5150), .IN2(r800_n166), .QN(r800_n163) );
  NAND2X0 r800_U163 ( .IN1(P1_N2359), .IN2(n7048), .QN(r800_n164) );
  NAND2X0 r800_U162 ( .IN1(r800_n163), .IN2(r800_n164), .QN(r800_n161) );
  NAND2X0 r800_U161 ( .IN1(r800_n161), .IN2(r800_n162), .QN(r800_n159) );
  OR2X1 r800_U160 ( .IN2(r800_n162), .IN1(r800_n161), .Q(r800_n160) );
  NAND2X0 r800_U159 ( .IN1(r800_n159), .IN2(r800_n160), .QN(P1_N2511) );
  INVX0 r800_U158 ( .ZN(r800_n145), .INP(P1_N2378) );
  NAND2X0 r800_U157 ( .IN1(P1_N5169), .IN2(r800_n145), .QN(r800_n157) );
  OR2X1 r800_U156 ( .IN2(P1_N5169), .IN1(r800_n145), .Q(r800_n158) );
  NAND2X0 r800_U155 ( .IN1(r800_n157), .IN2(r800_n158), .QN(r800_n151) );
  NAND2X0 r800_U154 ( .IN1(n7099), .IN2(r800_n156), .QN(r800_n152) );
  OR2X1 r800_U153 ( .IN2(n7099), .IN1(r800_n156), .Q(r800_n154) );
  NAND2X0 r800_U152 ( .IN1(r800_n154), .IN2(r800_n155), .QN(r800_n153) );
  NAND2X0 r800_U151 ( .IN1(r800_n152), .IN2(r800_n153), .QN(r800_n146) );
  NAND2X0 r800_U150 ( .IN1(r800_n151), .IN2(r800_n146), .QN(r800_n149) );
  OR2X1 r800_U149 ( .IN2(r800_n146), .IN1(r800_n151), .Q(r800_n150) );
  NAND2X0 r800_U148 ( .IN1(r800_n149), .IN2(r800_n150), .QN(P1_N2530) );
  INVX0 r800_U147 ( .ZN(r800_n135), .INP(P1_N2379) );
  NAND2X0 r800_U146 ( .IN1(P1_N5170), .IN2(r800_n135), .QN(r800_n147) );
  OR2X1 r800_U145 ( .IN2(P1_N5170), .IN1(r800_n135), .Q(r800_n148) );
  NAND2X0 r800_U144 ( .IN1(r800_n147), .IN2(r800_n148), .QN(r800_n141) );
  NAND2X0 r800_U143 ( .IN1(P1_N5169), .IN2(r800_n146), .QN(r800_n142) );
  OR2X1 r800_U142 ( .IN2(P1_N5169), .IN1(r800_n146), .Q(r800_n144) );
  NAND2X0 r800_U141 ( .IN1(r800_n144), .IN2(r800_n145), .QN(r800_n143) );
  NAND2X0 r800_U140 ( .IN1(r800_n142), .IN2(r800_n143), .QN(r800_n136) );
  NAND2X0 r800_U139 ( .IN1(r800_n141), .IN2(r800_n136), .QN(r800_n139) );
  OR2X1 r800_U138 ( .IN2(r800_n136), .IN1(r800_n141), .Q(r800_n140) );
  NAND2X0 r800_U137 ( .IN1(r800_n139), .IN2(r800_n140), .QN(P1_N2531) );
  INVX0 r800_U136 ( .ZN(r800_n125), .INP(P1_N2380) );
  NAND2X0 r800_U135 ( .IN1(P1_N5171), .IN2(r800_n125), .QN(r800_n137) );
  OR2X1 r800_U134 ( .IN2(P1_N5171), .IN1(r800_n125), .Q(r800_n138) );
  NAND2X0 r800_U133 ( .IN1(r800_n137), .IN2(r800_n138), .QN(r800_n131) );
  NAND2X0 r800_U132 ( .IN1(P1_N5170), .IN2(r800_n136), .QN(r800_n132) );
  OR2X1 r800_U131 ( .IN2(P1_N5170), .IN1(r800_n136), .Q(r800_n134) );
  NAND2X0 r800_U130 ( .IN1(r800_n134), .IN2(r800_n135), .QN(r800_n133) );
  NAND2X0 r800_U129 ( .IN1(r800_n132), .IN2(r800_n133), .QN(r800_n126) );
  NAND2X0 r800_U128 ( .IN1(r800_n131), .IN2(r800_n126), .QN(r800_n129) );
  OR2X1 r800_U127 ( .IN2(r800_n126), .IN1(r800_n131), .Q(r800_n130) );
  NAND2X0 r800_U126 ( .IN1(r800_n129), .IN2(r800_n130), .QN(P1_N2532) );
  INVX0 r800_U125 ( .ZN(r800_n115), .INP(P1_N2381) );
  NAND2X0 r800_U124 ( .IN1(n7141), .IN2(r800_n115), .QN(r800_n127) );
  OR2X1 r800_U123 ( .IN2(n7141), .IN1(r800_n115), .Q(r800_n128) );
  NAND2X0 r800_U122 ( .IN1(r800_n127), .IN2(r800_n128), .QN(r800_n121) );
  NAND2X0 r800_U121 ( .IN1(P1_N5171), .IN2(r800_n126), .QN(r800_n122) );
  OR2X1 r800_U120 ( .IN2(P1_N5171), .IN1(r800_n126), .Q(r800_n124) );
  NAND2X0 r800_U119 ( .IN1(r800_n124), .IN2(r800_n125), .QN(r800_n123) );
  NAND2X0 r800_U118 ( .IN1(r800_n122), .IN2(r800_n123), .QN(r800_n116) );
  NAND2X0 r800_U117 ( .IN1(r800_n121), .IN2(r800_n116), .QN(r800_n119) );
  OR2X1 r800_U116 ( .IN2(r800_n116), .IN1(r800_n121), .Q(r800_n120) );
  NAND2X0 r800_U115 ( .IN1(r800_n119), .IN2(r800_n120), .QN(P1_N2533) );
  INVX0 r800_U114 ( .ZN(r800_n105), .INP(P1_N2382) );
  NAND2X0 r800_U113 ( .IN1(n7138), .IN2(r800_n105), .QN(r800_n117) );
  OR2X1 r800_U112 ( .IN2(n7138), .IN1(r800_n105), .Q(r800_n118) );
  NAND2X0 r800_U111 ( .IN1(r800_n117), .IN2(r800_n118), .QN(r800_n111) );
  NAND2X0 r800_U110 ( .IN1(n7141), .IN2(r800_n116), .QN(r800_n112) );
  OR2X1 r800_U109 ( .IN2(n7141), .IN1(r800_n116), .Q(r800_n114) );
  NAND2X0 r800_U108 ( .IN1(r800_n114), .IN2(r800_n115), .QN(r800_n113) );
  NAND2X0 r800_U107 ( .IN1(r800_n112), .IN2(r800_n113), .QN(r800_n106) );
  NAND2X0 r800_U106 ( .IN1(r800_n111), .IN2(r800_n106), .QN(r800_n109) );
  OR2X1 r800_U105 ( .IN2(r800_n106), .IN1(r800_n111), .Q(r800_n110) );
  NAND2X0 r800_U104 ( .IN1(r800_n109), .IN2(r800_n110), .QN(P1_N2534) );
  INVX0 r800_U103 ( .ZN(r800_n95), .INP(P1_N2383) );
  NAND2X0 r800_U102 ( .IN1(P1_N5174), .IN2(r800_n95), .QN(r800_n107) );
  OR2X1 r800_U101 ( .IN2(P1_N5174), .IN1(r800_n95), .Q(r800_n108) );
  NAND2X0 r800_U100 ( .IN1(r800_n107), .IN2(r800_n108), .QN(r800_n101) );
  NAND2X0 r800_U99 ( .IN1(n7138), .IN2(r800_n106), .QN(r800_n102) );
  INVX0 r800_U284 ( .ZN(r800_n28), .INP(P1_N2364) );
  NAND2X0 r800_U283 ( .IN1(r800_n271), .IN2(r800_n28), .QN(r800_n270) );
  NAND2X0 r800_U282 ( .IN1(r800_n269), .IN2(r800_n270), .QN(r800_n18) );
  NAND2X0 r800_U281 ( .IN1(n7075), .IN2(r800_n18), .QN(r800_n266) );
  OR2X1 r800_U280 ( .IN2(n7075), .IN1(r800_n18), .Q(r800_n268) );
  INVX0 r800_U279 ( .ZN(r800_n21), .INP(P1_N2365) );
  NAND2X0 r800_U278 ( .IN1(r800_n268), .IN2(r800_n21), .QN(r800_n267) );
  NAND2X0 r800_U277 ( .IN1(r800_n266), .IN2(r800_n267), .QN(r800_n11) );
  NAND2X0 r800_U276 ( .IN1(n7072), .IN2(r800_n11), .QN(r800_n263) );
  OR2X1 r800_U275 ( .IN2(n7072), .IN1(r800_n11), .Q(r800_n265) );
  INVX0 r800_U274 ( .ZN(r800_n14), .INP(P1_N2366) );
  NAND2X0 r800_U273 ( .IN1(r800_n265), .IN2(r800_n14), .QN(r800_n264) );
  NAND2X0 r800_U272 ( .IN1(r800_n263), .IN2(r800_n264), .QN(r800_n4) );
  NAND2X0 r800_U271 ( .IN1(n7070), .IN2(r800_n4), .QN(r800_n260) );
  OR2X1 r800_U270 ( .IN2(n7070), .IN1(r800_n4), .Q(r800_n262) );
  INVX0 r800_U269 ( .ZN(r800_n7), .INP(P1_N2367) );
  NAND2X0 r800_U268 ( .IN1(r800_n262), .IN2(r800_n7), .QN(r800_n261) );
  NAND2X0 r800_U267 ( .IN1(r800_n260), .IN2(r800_n261), .QN(r800_n254) );
  NAND2X0 r800_U266 ( .IN1(r800_n259), .IN2(r800_n254), .QN(r800_n257) );
  OR2X1 r800_U265 ( .IN2(r800_n254), .IN1(r800_n259), .Q(r800_n258) );
  NAND2X0 r800_U264 ( .IN1(r800_n257), .IN2(r800_n258), .QN(P1_N2520) );
  INVX0 r800_U263 ( .ZN(r800_n243), .INP(P1_N2369) );
  NAND2X0 r800_U262 ( .IN1(P1_N5160), .IN2(r800_n243), .QN(r800_n255) );
  OR2X1 r800_U261 ( .IN2(P1_N5160), .IN1(r800_n243), .Q(r800_n256) );
  NAND2X0 r800_U260 ( .IN1(r800_n255), .IN2(r800_n256), .QN(r800_n249) );
  NAND2X0 r800_U259 ( .IN1(n7066), .IN2(r800_n254), .QN(r800_n250) );
  OR2X1 r800_U258 ( .IN2(n7066), .IN1(r800_n254), .Q(r800_n252) );
  NAND2X0 r800_U257 ( .IN1(r800_n252), .IN2(r800_n253), .QN(r800_n251) );
  NAND2X0 r800_U256 ( .IN1(r800_n250), .IN2(r800_n251), .QN(r800_n244) );
  NAND2X0 r800_U255 ( .IN1(r800_n249), .IN2(r800_n244), .QN(r800_n247) );
  OR2X1 r800_U254 ( .IN2(r800_n244), .IN1(r800_n249), .Q(r800_n248) );
  NAND2X0 r800_U253 ( .IN1(r800_n247), .IN2(r800_n248), .QN(P1_N2521) );
  INVX0 r800_U252 ( .ZN(r800_n233), .INP(P1_N2370) );
  NAND2X0 r800_U251 ( .IN1(n7059), .IN2(r800_n233), .QN(r800_n245) );
  OR2X1 r800_U250 ( .IN2(n7059), .IN1(r800_n233), .Q(r800_n246) );
  NAND2X0 r800_U249 ( .IN1(r800_n245), .IN2(r800_n246), .QN(r800_n239) );
  NAND2X0 r800_U248 ( .IN1(P1_N5160), .IN2(r800_n244), .QN(r800_n240) );
  OR2X1 r800_U247 ( .IN2(P1_N5160), .IN1(r800_n244), .Q(r800_n242) );
  NAND2X0 r800_U246 ( .IN1(r800_n242), .IN2(r800_n243), .QN(r800_n241) );
  NAND2X0 r800_U245 ( .IN1(r800_n240), .IN2(r800_n241), .QN(r800_n234) );
  NAND2X0 r800_U244 ( .IN1(r800_n239), .IN2(r800_n234), .QN(r800_n237) );
  OR2X1 r800_U243 ( .IN2(r800_n234), .IN1(r800_n239), .Q(r800_n238) );
  NAND2X0 r800_U242 ( .IN1(r800_n237), .IN2(r800_n238), .QN(P1_N2522) );
  INVX0 r800_U241 ( .ZN(r800_n223), .INP(P1_N2371) );
  NAND2X0 r800_U240 ( .IN1(n7055), .IN2(r800_n223), .QN(r800_n235) );
  OR2X1 r800_U239 ( .IN2(n7055), .IN1(r800_n223), .Q(r800_n236) );
  NAND2X0 r800_U238 ( .IN1(r800_n235), .IN2(r800_n236), .QN(r800_n229) );
  NAND2X0 r800_U237 ( .IN1(n7059), .IN2(r800_n234), .QN(r800_n230) );
  OR2X1 r800_U236 ( .IN2(n7059), .IN1(r800_n234), .Q(r800_n232) );
  NAND2X0 r800_U235 ( .IN1(r800_n232), .IN2(r800_n233), .QN(r800_n231) );
  NAND2X0 r800_U234 ( .IN1(r800_n230), .IN2(r800_n231), .QN(r800_n224) );
  NAND2X0 r800_U233 ( .IN1(r800_n229), .IN2(r800_n224), .QN(r800_n227) );
  OR2X1 r800_U232 ( .IN2(r800_n224), .IN1(r800_n229), .Q(r800_n228) );
  NAND2X0 r800_U231 ( .IN1(r800_n227), .IN2(r800_n228), .QN(P1_N2523) );
  INVX0 r800_U230 ( .ZN(r800_n213), .INP(P1_N2372) );
  NAND2X0 r800_U229 ( .IN1(P1_N5163), .IN2(r800_n213), .QN(r800_n225) );
  OR2X1 r800_U228 ( .IN2(P1_N5163), .IN1(r800_n213), .Q(r800_n226) );
  NAND2X0 r800_U227 ( .IN1(r800_n225), .IN2(r800_n226), .QN(r800_n219) );
  NAND2X0 r800_U226 ( .IN1(n7055), .IN2(r800_n224), .QN(r800_n220) );
  OR2X1 r800_U225 ( .IN2(n7055), .IN1(r800_n224), .Q(r800_n222) );
  NAND2X0 r800_U224 ( .IN1(r800_n222), .IN2(r800_n223), .QN(r800_n221) );
  NAND2X0 r800_U223 ( .IN1(r800_n220), .IN2(r800_n221), .QN(r800_n214) );
  NAND2X0 r800_U222 ( .IN1(r800_n219), .IN2(r800_n214), .QN(r800_n217) );
  OR2X1 r800_U221 ( .IN2(r800_n214), .IN1(r800_n219), .Q(r800_n218) );
  NAND2X0 r800_U220 ( .IN1(r800_n217), .IN2(r800_n218), .QN(P1_N2524) );
  INVX0 r800_U219 ( .ZN(r800_n203), .INP(P1_N2373) );
  NAND2X0 r800_U218 ( .IN1(n7113), .IN2(r800_n203), .QN(r800_n215) );
  OR2X1 r800_U217 ( .IN2(n7113), .IN1(r800_n203), .Q(r800_n216) );
  NAND2X0 r800_U216 ( .IN1(r800_n215), .IN2(r800_n216), .QN(r800_n209) );
  NAND2X0 r800_U215 ( .IN1(P1_N5163), .IN2(r800_n214), .QN(r800_n210) );
  OR2X1 r800_U214 ( .IN2(P1_N5163), .IN1(r800_n214), .Q(r800_n212) );
  NAND2X0 r800_U213 ( .IN1(r800_n212), .IN2(r800_n213), .QN(r800_n211) );
  NAND2X0 r800_U212 ( .IN1(r800_n210), .IN2(r800_n211), .QN(r800_n204) );
  NAND2X0 r800_U211 ( .IN1(r800_n209), .IN2(r800_n204), .QN(r800_n207) );
  OR2X1 r800_U210 ( .IN2(r800_n204), .IN1(r800_n209), .Q(r800_n208) );
  NAND2X0 r800_U209 ( .IN1(r800_n207), .IN2(r800_n208), .QN(P1_N2525) );
  INVX0 r800_U208 ( .ZN(r800_n193), .INP(P1_N2374) );
  NAND2X0 r800_U207 ( .IN1(n7110), .IN2(r800_n193), .QN(r800_n205) );
  OR2X1 r800_U206 ( .IN2(n7110), .IN1(r800_n193), .Q(r800_n206) );
  NAND2X0 r800_U205 ( .IN1(r800_n205), .IN2(r800_n206), .QN(r800_n199) );
  NAND2X0 r800_U204 ( .IN1(n7113), .IN2(r800_n204), .QN(r800_n200) );
  OR2X1 r800_U203 ( .IN2(n7113), .IN1(r800_n204), .Q(r800_n202) );
  NAND2X0 r800_U202 ( .IN1(r800_n202), .IN2(r800_n203), .QN(r800_n201) );
  NAND2X0 r800_U201 ( .IN1(r800_n200), .IN2(r800_n201), .QN(r800_n194) );
  NAND2X0 r800_U200 ( .IN1(r800_n199), .IN2(r800_n194), .QN(r800_n197) );
  OR2X1 r800_U199 ( .IN2(r800_n194), .IN1(r800_n199), .Q(r800_n198) );
  NAND2X0 r800_U198 ( .IN1(r800_n197), .IN2(r800_n198), .QN(P1_N2526) );
  INVX0 r800_U197 ( .ZN(r800_n183), .INP(P1_N2375) );
  NAND2X0 r800_U196 ( .IN1(n7106), .IN2(r800_n183), .QN(r800_n195) );
  OR2X1 r800_U195 ( .IN2(n7106), .IN1(r800_n183), .Q(r800_n196) );
  NAND2X0 r800_U194 ( .IN1(r800_n195), .IN2(r800_n196), .QN(r800_n189) );
  NAND2X0 r800_U193 ( .IN1(n7110), .IN2(r800_n194), .QN(r800_n190) );
  OR2X1 r800_U192 ( .IN2(n7110), .IN1(r800_n194), .Q(r800_n192) );
  INVX0 r800_U321 ( .ZN(r800_n291), .INP(P1_N2358) );
  NOR2X0 r800_U320 ( .QN(r800_n287), .IN1(r800_n291), .IN2(n7034) );
  INVX0 r800_U319 ( .ZN(r800_n162), .INP(r800_n287) );
  NAND2X0 r800_U318 ( .IN1(n7034), .IN2(r800_n291), .QN(r800_n290) );
  NAND2X0 r800_U317 ( .IN1(r800_n162), .IN2(r800_n290), .QN(P1_N2510) );
  INVX0 r800_U316 ( .ZN(r800_n253), .INP(P1_N2368) );
  NAND2X0 r800_U315 ( .IN1(n7066), .IN2(r800_n253), .QN(r800_n288) );
  OR2X1 r800_U314 ( .IN2(n7066), .IN1(r800_n253), .Q(r800_n289) );
  NAND2X0 r800_U313 ( .IN1(r800_n288), .IN2(r800_n289), .QN(r800_n259) );
  NAND2X0 r800_U312 ( .IN1(P1_N5150), .IN2(r800_n162), .QN(r800_n284) );
  NAND2X0 r800_U310 ( .IN1(r800_n287), .IN2(n7048), .QN(r800_n286) );
  INVX0 r800_U309 ( .ZN(r800_n166), .INP(P1_N2359) );
  NAND2X0 r800_U308 ( .IN1(r800_n286), .IN2(r800_n166), .QN(r800_n285) );
  NAND2X0 r800_U307 ( .IN1(r800_n284), .IN2(r800_n285), .QN(r800_n53) );
  NAND2X0 r800_U306 ( .IN1(P1_N5151), .IN2(r800_n53), .QN(r800_n281) );
  OR2X1 r800_U305 ( .IN2(P1_N5151), .IN1(r800_n53), .Q(r800_n283) );
  INVX0 r800_U304 ( .ZN(r800_n56), .INP(P1_N2360) );
  NAND2X0 r800_U303 ( .IN1(r800_n283), .IN2(r800_n56), .QN(r800_n282) );
  NAND2X0 r800_U302 ( .IN1(r800_n281), .IN2(r800_n282), .QN(r800_n46) );
  NAND2X0 r800_U301 ( .IN1(P1_N5152), .IN2(r800_n46), .QN(r800_n278) );
  OR2X1 r800_U300 ( .IN2(P1_N5152), .IN1(r800_n46), .Q(r800_n280) );
  INVX0 r800_U299 ( .ZN(r800_n49), .INP(P1_N2361) );
  NAND2X0 r800_U298 ( .IN1(r800_n280), .IN2(r800_n49), .QN(r800_n279) );
  NAND2X0 r800_U297 ( .IN1(r800_n278), .IN2(r800_n279), .QN(r800_n39) );
  NAND2X0 r800_U296 ( .IN1(P1_N5153), .IN2(r800_n39), .QN(r800_n275) );
  OR2X1 r800_U295 ( .IN2(P1_N5153), .IN1(r800_n39), .Q(r800_n277) );
  INVX0 r800_U294 ( .ZN(r800_n42), .INP(P1_N2362) );
  NAND2X0 r800_U293 ( .IN1(r800_n277), .IN2(r800_n42), .QN(r800_n276) );
  NAND2X0 r800_U292 ( .IN1(r800_n275), .IN2(r800_n276), .QN(r800_n32) );
  NAND2X0 r800_U291 ( .IN1(P1_N5154), .IN2(r800_n32), .QN(r800_n272) );
  OR2X1 r800_U290 ( .IN2(P1_N5154), .IN1(r800_n32), .Q(r800_n274) );
  INVX0 r800_U289 ( .ZN(r800_n35), .INP(P1_N2363) );
  NAND2X0 r800_U288 ( .IN1(r800_n274), .IN2(r800_n35), .QN(r800_n273) );
  NAND2X0 r800_U287 ( .IN1(r800_n272), .IN2(r800_n273), .QN(r800_n25) );
  NAND2X0 r800_U286 ( .IN1(n7080), .IN2(r800_n25), .QN(r800_n269) );
  OR2X1 r800_U285 ( .IN2(n7080), .IN1(r800_n25), .Q(r800_n271) );
  OR2X1 r802_U47 ( .IN2(P1_N5151), .IN1(r802_n56), .Q(r802_n55) );
  NAND2X0 r802_U46 ( .IN1(r802_n54), .IN2(r802_n55), .QN(r802_n52) );
  NAND2X0 r802_U45 ( .IN1(r802_n52), .IN2(r802_n53), .QN(r802_n50) );
  OR2X1 r802_U44 ( .IN2(r802_n53), .IN1(r802_n52), .Q(r802_n51) );
  NAND2X0 r802_U43 ( .IN1(r802_n50), .IN2(r802_n51), .QN(P1_N2885) );
  NAND2X0 r802_U42 ( .IN1(n7041), .IN2(r802_n49), .QN(r802_n47) );
  OR2X1 r802_U41 ( .IN2(n7041), .IN1(r802_n49), .Q(r802_n48) );
  NAND2X0 r802_U40 ( .IN1(r802_n47), .IN2(r802_n48), .QN(r802_n45) );
  NAND2X0 r802_U39 ( .IN1(r802_n45), .IN2(r802_n46), .QN(r802_n43) );
  OR2X1 r802_U38 ( .IN2(r802_n46), .IN1(r802_n45), .Q(r802_n44) );
  NAND2X0 r802_U37 ( .IN1(r802_n43), .IN2(r802_n44), .QN(P1_N2886) );
  NAND2X0 r802_U36 ( .IN1(P1_N5153), .IN2(r802_n42), .QN(r802_n40) );
  OR2X1 r802_U35 ( .IN2(P1_N5153), .IN1(r802_n42), .Q(r802_n41) );
  NAND2X0 r802_U34 ( .IN1(r802_n40), .IN2(r802_n41), .QN(r802_n38) );
  NAND2X0 r802_U33 ( .IN1(r802_n38), .IN2(r802_n39), .QN(r802_n36) );
  OR2X1 r802_U32 ( .IN2(r802_n39), .IN1(r802_n38), .Q(r802_n37) );
  NAND2X0 r802_U31 ( .IN1(r802_n36), .IN2(r802_n37), .QN(P1_N2887) );
  NAND2X0 r802_U30 ( .IN1(n7081), .IN2(r802_n35), .QN(r802_n33) );
  OR2X1 r802_U29 ( .IN2(n7081), .IN1(r802_n35), .Q(r802_n34) );
  NAND2X0 r802_U28 ( .IN1(r802_n33), .IN2(r802_n34), .QN(r802_n31) );
  NAND2X0 r802_U27 ( .IN1(r802_n31), .IN2(r802_n32), .QN(r802_n29) );
  OR2X1 r802_U26 ( .IN2(r802_n32), .IN1(r802_n31), .Q(r802_n30) );
  NAND2X0 r802_U25 ( .IN1(r802_n29), .IN2(r802_n30), .QN(P1_N2888) );
  NAND2X0 r802_U24 ( .IN1(P1_N5155), .IN2(r802_n28), .QN(r802_n26) );
  OR2X1 r802_U23 ( .IN2(P1_N5155), .IN1(r802_n28), .Q(r802_n27) );
  NAND2X0 r802_U22 ( .IN1(r802_n26), .IN2(r802_n27), .QN(r802_n24) );
  NAND2X0 r802_U21 ( .IN1(r802_n24), .IN2(r802_n25), .QN(r802_n22) );
  OR2X1 r802_U20 ( .IN2(r802_n25), .IN1(r802_n24), .Q(r802_n23) );
  NAND2X0 r802_U19 ( .IN1(r802_n22), .IN2(r802_n23), .QN(P1_N2889) );
  NAND2X0 r802_U18 ( .IN1(n7075), .IN2(r802_n21), .QN(r802_n19) );
  OR2X1 r802_U17 ( .IN2(n7075), .IN1(r802_n21), .Q(r802_n20) );
  NAND2X0 r802_U16 ( .IN1(r802_n19), .IN2(r802_n20), .QN(r802_n17) );
  NAND2X0 r802_U15 ( .IN1(r802_n17), .IN2(r802_n18), .QN(r802_n15) );
  OR2X1 r802_U14 ( .IN2(r802_n18), .IN1(r802_n17), .Q(r802_n16) );
  NAND2X0 r802_U13 ( .IN1(r802_n15), .IN2(r802_n16), .QN(P1_N2890) );
  NAND2X0 r802_U12 ( .IN1(n7072), .IN2(r802_n14), .QN(r802_n12) );
  OR2X1 r802_U11 ( .IN2(n7072), .IN1(r802_n14), .Q(r802_n13) );
  NAND2X0 r802_U10 ( .IN1(r802_n12), .IN2(r802_n13), .QN(r802_n10) );
  NAND2X0 r802_U9 ( .IN1(r802_n10), .IN2(r802_n11), .QN(r802_n8) );
  OR2X1 r802_U8 ( .IN2(r802_n11), .IN1(r802_n10), .Q(r802_n9) );
  NAND2X0 r802_U7 ( .IN1(r802_n8), .IN2(r802_n9), .QN(P1_N2891) );
  NAND2X0 r802_U6 ( .IN1(P1_N5158), .IN2(r802_n7), .QN(r802_n5) );
  OR2X1 r802_U5 ( .IN2(P1_N5158), .IN1(r802_n7), .Q(r802_n6) );
  NAND2X0 r802_U4 ( .IN1(r802_n5), .IN2(r802_n6), .QN(r802_n3) );
  NAND2X0 r802_U3 ( .IN1(r802_n3), .IN2(r802_n4), .QN(r802_n1) );
  OR2X1 r802_U2 ( .IN2(r802_n4), .IN1(r802_n3), .Q(r802_n2) );
  NAND2X0 r802_U1 ( .IN1(r802_n1), .IN2(r802_n2), .QN(P1_N2892) );
  NAND2X0 r802_U140 ( .IN1(r802_n142), .IN2(r802_n143), .QN(r802_n136) );
  NAND2X0 r802_U139 ( .IN1(r802_n141), .IN2(r802_n136), .QN(r802_n139) );
  OR2X1 r802_U138 ( .IN2(r802_n136), .IN1(r802_n141), .Q(r802_n140) );
  NAND2X0 r802_U137 ( .IN1(r802_n139), .IN2(r802_n140), .QN(P1_N2904) );
  INVX0 r802_U136 ( .ZN(r802_n125), .INP(P1_N2753) );
  NAND2X0 r802_U135 ( .IN1(n7089), .IN2(r802_n125), .QN(r802_n137) );
  OR2X1 r802_U134 ( .IN2(n7089), .IN1(r802_n125), .Q(r802_n138) );
  NAND2X0 r802_U133 ( .IN1(r802_n137), .IN2(r802_n138), .QN(r802_n131) );
  NAND2X0 r802_U132 ( .IN1(n7093), .IN2(r802_n136), .QN(r802_n132) );
  OR2X1 r802_U131 ( .IN2(n7093), .IN1(r802_n136), .Q(r802_n134) );
  NAND2X0 r802_U130 ( .IN1(r802_n134), .IN2(r802_n135), .QN(r802_n133) );
  NAND2X0 r802_U129 ( .IN1(r802_n132), .IN2(r802_n133), .QN(r802_n126) );
  NAND2X0 r802_U128 ( .IN1(r802_n131), .IN2(r802_n126), .QN(r802_n129) );
  OR2X1 r802_U127 ( .IN2(r802_n126), .IN1(r802_n131), .Q(r802_n130) );
  NAND2X0 r802_U126 ( .IN1(r802_n129), .IN2(r802_n130), .QN(P1_N2905) );
  INVX0 r802_U125 ( .ZN(r802_n115), .INP(P1_N2754) );
  NAND2X0 r802_U124 ( .IN1(P1_N5172), .IN2(r802_n115), .QN(r802_n127) );
  OR2X1 r802_U123 ( .IN2(P1_N5172), .IN1(r802_n115), .Q(r802_n128) );
  NAND2X0 r802_U122 ( .IN1(r802_n127), .IN2(r802_n128), .QN(r802_n121) );
  NAND2X0 r802_U121 ( .IN1(n7089), .IN2(r802_n126), .QN(r802_n122) );
  OR2X1 r802_U120 ( .IN2(n7089), .IN1(r802_n126), .Q(r802_n124) );
  NAND2X0 r802_U119 ( .IN1(r802_n124), .IN2(r802_n125), .QN(r802_n123) );
  NAND2X0 r802_U118 ( .IN1(r802_n122), .IN2(r802_n123), .QN(r802_n116) );
  NAND2X0 r802_U117 ( .IN1(r802_n121), .IN2(r802_n116), .QN(r802_n119) );
  OR2X1 r802_U116 ( .IN2(r802_n116), .IN1(r802_n121), .Q(r802_n120) );
  NAND2X0 r802_U115 ( .IN1(r802_n119), .IN2(r802_n120), .QN(P1_N2906) );
  INVX0 r802_U114 ( .ZN(r802_n105), .INP(P1_N2755) );
  NAND2X0 r802_U113 ( .IN1(n7138), .IN2(r802_n105), .QN(r802_n117) );
  OR2X1 r802_U112 ( .IN2(n7138), .IN1(r802_n105), .Q(r802_n118) );
  NAND2X0 r802_U111 ( .IN1(r802_n117), .IN2(r802_n118), .QN(r802_n111) );
  NAND2X0 r802_U110 ( .IN1(P1_N5172), .IN2(r802_n116), .QN(r802_n112) );
  OR2X1 r802_U109 ( .IN2(P1_N5172), .IN1(r802_n116), .Q(r802_n114) );
  NAND2X0 r802_U108 ( .IN1(r802_n114), .IN2(r802_n115), .QN(r802_n113) );
  NAND2X0 r802_U107 ( .IN1(r802_n112), .IN2(r802_n113), .QN(r802_n106) );
  NAND2X0 r802_U106 ( .IN1(r802_n111), .IN2(r802_n106), .QN(r802_n109) );
  OR2X1 r802_U105 ( .IN2(r802_n106), .IN1(r802_n111), .Q(r802_n110) );
  NAND2X0 r802_U104 ( .IN1(r802_n109), .IN2(r802_n110), .QN(P1_N2907) );
  INVX0 r802_U103 ( .ZN(r802_n95), .INP(P1_N2756) );
  NAND2X0 r802_U102 ( .IN1(P1_N5174), .IN2(r802_n95), .QN(r802_n107) );
  OR2X1 r802_U101 ( .IN2(P1_N5174), .IN1(r802_n95), .Q(r802_n108) );
  NAND2X0 r802_U100 ( .IN1(r802_n107), .IN2(r802_n108), .QN(r802_n101) );
  NAND2X0 r802_U99 ( .IN1(n7138), .IN2(r802_n106), .QN(r802_n102) );
  OR2X1 r802_U98 ( .IN2(n7138), .IN1(r802_n106), .Q(r802_n104) );
  NAND2X0 r802_U97 ( .IN1(r802_n104), .IN2(r802_n105), .QN(r802_n103) );
  NAND2X0 r802_U96 ( .IN1(r802_n102), .IN2(r802_n103), .QN(r802_n96) );
  NAND2X0 r802_U95 ( .IN1(r802_n101), .IN2(r802_n96), .QN(r802_n99) );
  OR2X1 r802_U94 ( .IN2(r802_n96), .IN1(r802_n101), .Q(r802_n100) );
  NAND2X0 r802_U93 ( .IN1(r802_n99), .IN2(r802_n100), .QN(P1_N2908) );
  INVX0 r802_U92 ( .ZN(r802_n85), .INP(P1_N2757) );
  NAND2X0 r802_U91 ( .IN1(n7124), .IN2(r802_n85), .QN(r802_n97) );
  OR2X1 r802_U90 ( .IN2(n7124), .IN1(r802_n85), .Q(r802_n98) );
  NAND2X0 r802_U89 ( .IN1(r802_n97), .IN2(r802_n98), .QN(r802_n91) );
  NAND2X0 r802_U88 ( .IN1(P1_N5174), .IN2(r802_n96), .QN(r802_n92) );
  OR2X1 r802_U87 ( .IN2(P1_N5174), .IN1(r802_n96), .Q(r802_n94) );
  NAND2X0 r802_U86 ( .IN1(r802_n94), .IN2(r802_n95), .QN(r802_n93) );
  NAND2X0 r802_U85 ( .IN1(r802_n92), .IN2(r802_n93), .QN(r802_n86) );
  NAND2X0 r802_U84 ( .IN1(r802_n91), .IN2(r802_n86), .QN(r802_n89) );
  OR2X1 r802_U83 ( .IN2(r802_n86), .IN1(r802_n91), .Q(r802_n90) );
  NAND2X0 r802_U82 ( .IN1(r802_n89), .IN2(r802_n90), .QN(P1_N2909) );
  INVX0 r802_U81 ( .ZN(r802_n75), .INP(P1_N2758) );
  NAND2X0 r802_U80 ( .IN1(n7122), .IN2(r802_n75), .QN(r802_n87) );
  OR2X1 r802_U79 ( .IN2(n7122), .IN1(r802_n75), .Q(r802_n88) );
  NAND2X0 r802_U78 ( .IN1(r802_n87), .IN2(r802_n88), .QN(r802_n81) );
  NAND2X0 r802_U77 ( .IN1(n7124), .IN2(r802_n86), .QN(r802_n82) );
  OR2X1 r802_U76 ( .IN2(n7124), .IN1(r802_n86), .Q(r802_n84) );
  NAND2X0 r802_U75 ( .IN1(r802_n84), .IN2(r802_n85), .QN(r802_n83) );
  NAND2X0 r802_U74 ( .IN1(r802_n82), .IN2(r802_n83), .QN(r802_n76) );
  NAND2X0 r802_U73 ( .IN1(r802_n81), .IN2(r802_n76), .QN(r802_n79) );
  OR2X1 r802_U72 ( .IN2(r802_n76), .IN1(r802_n81), .Q(r802_n80) );
  NAND2X0 r802_U71 ( .IN1(r802_n79), .IN2(r802_n80), .QN(P1_N2910) );
  INVX0 r802_U70 ( .ZN(r802_n64), .INP(P1_N2759) );
  NAND2X0 r802_U69 ( .IN1(P1_N5177), .IN2(r802_n64), .QN(r802_n77) );
  OR2X1 r802_U68 ( .IN2(P1_N5177), .IN1(r802_n64), .Q(r802_n78) );
  NAND2X0 r802_U67 ( .IN1(r802_n77), .IN2(r802_n78), .QN(r802_n71) );
  NAND2X0 r802_U66 ( .IN1(n7122), .IN2(r802_n76), .QN(r802_n72) );
  OR2X1 r802_U65 ( .IN2(n7122), .IN1(r802_n76), .Q(r802_n74) );
  NAND2X0 r802_U64 ( .IN1(r802_n74), .IN2(r802_n75), .QN(r802_n73) );
  NAND2X0 r802_U63 ( .IN1(r802_n72), .IN2(r802_n73), .QN(r802_n65) );
  NAND2X0 r802_U62 ( .IN1(r802_n71), .IN2(r802_n65), .QN(r802_n69) );
  OR2X1 r802_U61 ( .IN2(r802_n65), .IN1(r802_n71), .Q(r802_n70) );
  NAND2X0 r802_U60 ( .IN1(r802_n69), .IN2(r802_n70), .QN(P1_N2911) );
  OR2X1 r802_U58 ( .IN2(P1_N2760), .IN1(n7146), .Q(r802_n66) );
  NAND2X0 r802_U57 ( .IN1(P1_N2760), .IN2(n7146), .QN(r802_n67) );
  NAND2X0 r802_U56 ( .IN1(r802_n66), .IN2(r802_n67), .QN(r802_n60) );
  NAND2X0 r802_U55 ( .IN1(P1_N5177), .IN2(r802_n65), .QN(r802_n61) );
  OR2X1 r802_U54 ( .IN2(P1_N5177), .IN1(r802_n65), .Q(r802_n63) );
  NAND2X0 r802_U53 ( .IN1(r802_n63), .IN2(r802_n64), .QN(r802_n62) );
  NAND2X0 r802_U52 ( .IN1(r802_n61), .IN2(r802_n62), .QN(r802_n59) );
  NAND2X0 r802_U51 ( .IN1(r802_n60), .IN2(r802_n59), .QN(r802_n57) );
  OR2X1 r802_U50 ( .IN2(r802_n60), .IN1(r802_n59), .Q(r802_n58) );
  NAND2X0 r802_U49 ( .IN1(r802_n57), .IN2(r802_n58), .QN(P1_N2912) );
  NAND2X0 r802_U48 ( .IN1(P1_N5151), .IN2(r802_n56), .QN(r802_n54) );
  NAND2X0 r802_U233 ( .IN1(r802_n229), .IN2(r802_n224), .QN(r802_n227) );
  OR2X1 r802_U232 ( .IN2(r802_n224), .IN1(r802_n229), .Q(r802_n228) );
  NAND2X0 r802_U231 ( .IN1(r802_n227), .IN2(r802_n228), .QN(P1_N2896) );
  INVX0 r802_U230 ( .ZN(r802_n213), .INP(P1_N2745) );
  NAND2X0 r802_U229 ( .IN1(P1_N5163), .IN2(r802_n213), .QN(r802_n225) );
  OR2X1 r802_U228 ( .IN2(P1_N5163), .IN1(r802_n213), .Q(r802_n226) );
  NAND2X0 r802_U227 ( .IN1(r802_n225), .IN2(r802_n226), .QN(r802_n219) );
  NAND2X0 r802_U226 ( .IN1(P1_N5162), .IN2(r802_n224), .QN(r802_n220) );
  OR2X1 r802_U225 ( .IN2(P1_N5162), .IN1(r802_n224), .Q(r802_n222) );
  NAND2X0 r802_U224 ( .IN1(r802_n222), .IN2(r802_n223), .QN(r802_n221) );
  NAND2X0 r802_U223 ( .IN1(r802_n220), .IN2(r802_n221), .QN(r802_n214) );
  NAND2X0 r802_U222 ( .IN1(r802_n219), .IN2(r802_n214), .QN(r802_n217) );
  OR2X1 r802_U221 ( .IN2(r802_n214), .IN1(r802_n219), .Q(r802_n218) );
  NAND2X0 r802_U220 ( .IN1(r802_n217), .IN2(r802_n218), .QN(P1_N2897) );
  INVX0 r802_U219 ( .ZN(r802_n203), .INP(P1_N2746) );
  NAND2X0 r802_U218 ( .IN1(P1_N5164), .IN2(r802_n203), .QN(r802_n215) );
  OR2X1 r802_U217 ( .IN2(P1_N5164), .IN1(r802_n203), .Q(r802_n216) );
  NAND2X0 r802_U216 ( .IN1(r802_n215), .IN2(r802_n216), .QN(r802_n209) );
  NAND2X0 r802_U215 ( .IN1(P1_N5163), .IN2(r802_n214), .QN(r802_n210) );
  OR2X1 r802_U214 ( .IN2(P1_N5163), .IN1(r802_n214), .Q(r802_n212) );
  NAND2X0 r802_U213 ( .IN1(r802_n212), .IN2(r802_n213), .QN(r802_n211) );
  NAND2X0 r802_U212 ( .IN1(r802_n210), .IN2(r802_n211), .QN(r802_n204) );
  NAND2X0 r802_U211 ( .IN1(r802_n209), .IN2(r802_n204), .QN(r802_n207) );
  OR2X1 r802_U210 ( .IN2(r802_n204), .IN1(r802_n209), .Q(r802_n208) );
  NAND2X0 r802_U209 ( .IN1(r802_n207), .IN2(r802_n208), .QN(P1_N2898) );
  INVX0 r802_U208 ( .ZN(r802_n193), .INP(P1_N2747) );
  NAND2X0 r802_U207 ( .IN1(P1_N5165), .IN2(r802_n193), .QN(r802_n205) );
  OR2X1 r802_U206 ( .IN2(P1_N5165), .IN1(r802_n193), .Q(r802_n206) );
  NAND2X0 r802_U205 ( .IN1(r802_n205), .IN2(r802_n206), .QN(r802_n199) );
  NAND2X0 r802_U204 ( .IN1(P1_N5164), .IN2(r802_n204), .QN(r802_n200) );
  OR2X1 r802_U203 ( .IN2(P1_N5164), .IN1(r802_n204), .Q(r802_n202) );
  NAND2X0 r802_U202 ( .IN1(r802_n202), .IN2(r802_n203), .QN(r802_n201) );
  NAND2X0 r802_U201 ( .IN1(r802_n200), .IN2(r802_n201), .QN(r802_n194) );
  NAND2X0 r802_U200 ( .IN1(r802_n199), .IN2(r802_n194), .QN(r802_n197) );
  OR2X1 r802_U199 ( .IN2(r802_n194), .IN1(r802_n199), .Q(r802_n198) );
  NAND2X0 r802_U198 ( .IN1(r802_n197), .IN2(r802_n198), .QN(P1_N2899) );
  INVX0 r802_U197 ( .ZN(r802_n183), .INP(P1_N2748) );
  NAND2X0 r802_U196 ( .IN1(n7106), .IN2(r802_n183), .QN(r802_n195) );
  OR2X1 r802_U195 ( .IN2(n7106), .IN1(r802_n183), .Q(r802_n196) );
  NAND2X0 r802_U194 ( .IN1(r802_n195), .IN2(r802_n196), .QN(r802_n189) );
  NAND2X0 r802_U193 ( .IN1(P1_N5165), .IN2(r802_n194), .QN(r802_n190) );
  OR2X1 r802_U192 ( .IN2(P1_N5165), .IN1(r802_n194), .Q(r802_n192) );
  NAND2X0 r802_U191 ( .IN1(r802_n192), .IN2(r802_n193), .QN(r802_n191) );
  NAND2X0 r802_U190 ( .IN1(r802_n190), .IN2(r802_n191), .QN(r802_n184) );
  NAND2X0 r802_U189 ( .IN1(r802_n189), .IN2(r802_n184), .QN(r802_n187) );
  OR2X1 r802_U188 ( .IN2(r802_n184), .IN1(r802_n189), .Q(r802_n188) );
  NAND2X0 r802_U187 ( .IN1(r802_n187), .IN2(r802_n188), .QN(P1_N2900) );
  INVX0 r802_U186 ( .ZN(r802_n173), .INP(P1_N2749) );
  NAND2X0 r802_U185 ( .IN1(P1_N5167), .IN2(r802_n173), .QN(r802_n185) );
  OR2X1 r802_U184 ( .IN2(P1_N5167), .IN1(r802_n173), .Q(r802_n186) );
  NAND2X0 r802_U183 ( .IN1(r802_n185), .IN2(r802_n186), .QN(r802_n179) );
  NAND2X0 r802_U182 ( .IN1(n7106), .IN2(r802_n184), .QN(r802_n180) );
  OR2X1 r802_U181 ( .IN2(n7106), .IN1(r802_n184), .Q(r802_n182) );
  NAND2X0 r802_U180 ( .IN1(r802_n182), .IN2(r802_n183), .QN(r802_n181) );
  NAND2X0 r802_U179 ( .IN1(r802_n180), .IN2(r802_n181), .QN(r802_n174) );
  NAND2X0 r802_U178 ( .IN1(r802_n179), .IN2(r802_n174), .QN(r802_n177) );
  OR2X1 r802_U177 ( .IN2(r802_n174), .IN1(r802_n179), .Q(r802_n178) );
  NAND2X0 r802_U176 ( .IN1(r802_n177), .IN2(r802_n178), .QN(P1_N2901) );
  INVX0 r802_U175 ( .ZN(r802_n155), .INP(P1_N2750) );
  NAND2X0 r802_U174 ( .IN1(n7099), .IN2(r802_n155), .QN(r802_n175) );
  OR2X1 r802_U173 ( .IN2(n7099), .IN1(r802_n155), .Q(r802_n176) );
  NAND2X0 r802_U172 ( .IN1(r802_n175), .IN2(r802_n176), .QN(r802_n169) );
  NAND2X0 r802_U171 ( .IN1(P1_N5167), .IN2(r802_n174), .QN(r802_n170) );
  OR2X1 r802_U170 ( .IN2(P1_N5167), .IN1(r802_n174), .Q(r802_n172) );
  NAND2X0 r802_U169 ( .IN1(r802_n172), .IN2(r802_n173), .QN(r802_n171) );
  NAND2X0 r802_U168 ( .IN1(r802_n170), .IN2(r802_n171), .QN(r802_n156) );
  NAND2X0 r802_U167 ( .IN1(r802_n169), .IN2(r802_n156), .QN(r802_n167) );
  OR2X1 r802_U166 ( .IN2(r802_n156), .IN1(r802_n169), .Q(r802_n168) );
  NAND2X0 r802_U165 ( .IN1(r802_n167), .IN2(r802_n168), .QN(P1_N2902) );
  NAND2X0 r802_U164 ( .IN1(P1_N5150), .IN2(r802_n166), .QN(r802_n163) );
  NAND2X0 r802_U163 ( .IN1(P1_N2732), .IN2(n7048), .QN(r802_n164) );
  NAND2X0 r802_U162 ( .IN1(r802_n163), .IN2(r802_n164), .QN(r802_n161) );
  NAND2X0 r802_U161 ( .IN1(r802_n161), .IN2(r802_n162), .QN(r802_n159) );
  OR2X1 r802_U160 ( .IN2(r802_n162), .IN1(r802_n161), .Q(r802_n160) );
  NAND2X0 r802_U159 ( .IN1(r802_n159), .IN2(r802_n160), .QN(P1_N2884) );
  INVX0 r802_U158 ( .ZN(r802_n145), .INP(P1_N2751) );
  NAND2X0 r802_U157 ( .IN1(P1_N5169), .IN2(r802_n145), .QN(r802_n157) );
  OR2X1 r802_U156 ( .IN2(P1_N5169), .IN1(r802_n145), .Q(r802_n158) );
  NAND2X0 r802_U155 ( .IN1(r802_n157), .IN2(r802_n158), .QN(r802_n151) );
  NAND2X0 r802_U154 ( .IN1(P1_N5168), .IN2(r802_n156), .QN(r802_n152) );
  OR2X1 r802_U153 ( .IN2(P1_N5168), .IN1(r802_n156), .Q(r802_n154) );
  NAND2X0 r802_U152 ( .IN1(r802_n154), .IN2(r802_n155), .QN(r802_n153) );
  NAND2X0 r802_U151 ( .IN1(r802_n152), .IN2(r802_n153), .QN(r802_n146) );
  NAND2X0 r802_U150 ( .IN1(r802_n151), .IN2(r802_n146), .QN(r802_n149) );
  OR2X1 r802_U149 ( .IN2(r802_n146), .IN1(r802_n151), .Q(r802_n150) );
  NAND2X0 r802_U148 ( .IN1(r802_n149), .IN2(r802_n150), .QN(P1_N2903) );
  INVX0 r802_U147 ( .ZN(r802_n135), .INP(P1_N2752) );
  NAND2X0 r802_U146 ( .IN1(n7093), .IN2(r802_n135), .QN(r802_n147) );
  OR2X1 r802_U145 ( .IN2(n7093), .IN1(r802_n135), .Q(r802_n148) );
  NAND2X0 r802_U144 ( .IN1(r802_n147), .IN2(r802_n148), .QN(r802_n141) );
  NAND2X0 r802_U143 ( .IN1(P1_N5169), .IN2(r802_n146), .QN(r802_n142) );
  OR2X1 r802_U142 ( .IN2(P1_N5169), .IN1(r802_n146), .Q(r802_n144) );
  NAND2X0 r802_U141 ( .IN1(r802_n144), .IN2(r802_n145), .QN(r802_n143) );
  INVX0 r802_U321 ( .ZN(r802_n291), .INP(P1_N2731) );
  NOR2X0 r802_U320 ( .QN(r802_n287), .IN1(r802_n291), .IN2(n7034) );
  INVX0 r802_U319 ( .ZN(r802_n162), .INP(r802_n287) );
  NAND2X0 r802_U318 ( .IN1(n7034), .IN2(r802_n291), .QN(r802_n290) );
  NAND2X0 r802_U317 ( .IN1(r802_n162), .IN2(r802_n290), .QN(P1_N2883) );
  INVX0 r802_U316 ( .ZN(r802_n253), .INP(P1_N2741) );
  NAND2X0 r802_U315 ( .IN1(n7066), .IN2(r802_n253), .QN(r802_n288) );
  OR2X1 r802_U314 ( .IN2(n7066), .IN1(r802_n253), .Q(r802_n289) );
  NAND2X0 r802_U313 ( .IN1(r802_n288), .IN2(r802_n289), .QN(r802_n259) );
  NAND2X0 r802_U312 ( .IN1(P1_N5150), .IN2(r802_n162), .QN(r802_n284) );
  NAND2X0 r802_U310 ( .IN1(r802_n287), .IN2(n7048), .QN(r802_n286) );
  INVX0 r802_U309 ( .ZN(r802_n166), .INP(P1_N2732) );
  NAND2X0 r802_U308 ( .IN1(r802_n286), .IN2(r802_n166), .QN(r802_n285) );
  NAND2X0 r802_U307 ( .IN1(r802_n284), .IN2(r802_n285), .QN(r802_n53) );
  NAND2X0 r802_U306 ( .IN1(P1_N5151), .IN2(r802_n53), .QN(r802_n281) );
  OR2X1 r802_U305 ( .IN2(P1_N5151), .IN1(r802_n53), .Q(r802_n283) );
  INVX0 r802_U304 ( .ZN(r802_n56), .INP(P1_N2733) );
  NAND2X0 r802_U303 ( .IN1(r802_n283), .IN2(r802_n56), .QN(r802_n282) );
  NAND2X0 r802_U302 ( .IN1(r802_n281), .IN2(r802_n282), .QN(r802_n46) );
  NAND2X0 r802_U301 ( .IN1(n7041), .IN2(r802_n46), .QN(r802_n278) );
  OR2X1 r802_U300 ( .IN2(n7041), .IN1(r802_n46), .Q(r802_n280) );
  INVX0 r802_U299 ( .ZN(r802_n49), .INP(P1_N2734) );
  NAND2X0 r802_U298 ( .IN1(r802_n280), .IN2(r802_n49), .QN(r802_n279) );
  NAND2X0 r802_U297 ( .IN1(r802_n278), .IN2(r802_n279), .QN(r802_n39) );
  NAND2X0 r802_U296 ( .IN1(P1_N5153), .IN2(r802_n39), .QN(r802_n275) );
  OR2X1 r802_U295 ( .IN2(P1_N5153), .IN1(r802_n39), .Q(r802_n277) );
  INVX0 r802_U294 ( .ZN(r802_n42), .INP(P1_N2735) );
  NAND2X0 r802_U293 ( .IN1(r802_n277), .IN2(r802_n42), .QN(r802_n276) );
  NAND2X0 r802_U292 ( .IN1(r802_n275), .IN2(r802_n276), .QN(r802_n32) );
  NAND2X0 r802_U291 ( .IN1(n7081), .IN2(r802_n32), .QN(r802_n272) );
  OR2X1 r802_U290 ( .IN2(n7081), .IN1(r802_n32), .Q(r802_n274) );
  INVX0 r802_U289 ( .ZN(r802_n35), .INP(P1_N2736) );
  NAND2X0 r802_U288 ( .IN1(r802_n274), .IN2(r802_n35), .QN(r802_n273) );
  NAND2X0 r802_U287 ( .IN1(r802_n272), .IN2(r802_n273), .QN(r802_n25) );
  NAND2X0 r802_U286 ( .IN1(n7080), .IN2(r802_n25), .QN(r802_n269) );
  OR2X1 r802_U285 ( .IN2(P1_N5155), .IN1(r802_n25), .Q(r802_n271) );
  INVX0 r802_U284 ( .ZN(r802_n28), .INP(P1_N2737) );
  NAND2X0 r802_U283 ( .IN1(r802_n271), .IN2(r802_n28), .QN(r802_n270) );
  NAND2X0 r802_U282 ( .IN1(r802_n269), .IN2(r802_n270), .QN(r802_n18) );
  NAND2X0 r802_U281 ( .IN1(n7075), .IN2(r802_n18), .QN(r802_n266) );
  OR2X1 r802_U280 ( .IN2(n7075), .IN1(r802_n18), .Q(r802_n268) );
  INVX0 r802_U279 ( .ZN(r802_n21), .INP(P1_N2738) );
  NAND2X0 r802_U278 ( .IN1(r802_n268), .IN2(r802_n21), .QN(r802_n267) );
  NAND2X0 r802_U277 ( .IN1(r802_n266), .IN2(r802_n267), .QN(r802_n11) );
  NAND2X0 r802_U276 ( .IN1(n7072), .IN2(r802_n11), .QN(r802_n263) );
  OR2X1 r802_U275 ( .IN2(n7072), .IN1(r802_n11), .Q(r802_n265) );
  INVX0 r802_U274 ( .ZN(r802_n14), .INP(P1_N2739) );
  NAND2X0 r802_U273 ( .IN1(r802_n265), .IN2(r802_n14), .QN(r802_n264) );
  NAND2X0 r802_U272 ( .IN1(r802_n263), .IN2(r802_n264), .QN(r802_n4) );
  NAND2X0 r802_U271 ( .IN1(P1_N5158), .IN2(r802_n4), .QN(r802_n260) );
  OR2X1 r802_U270 ( .IN2(P1_N5158), .IN1(r802_n4), .Q(r802_n262) );
  INVX0 r802_U269 ( .ZN(r802_n7), .INP(P1_N2740) );
  NAND2X0 r802_U268 ( .IN1(r802_n262), .IN2(r802_n7), .QN(r802_n261) );
  NAND2X0 r802_U267 ( .IN1(r802_n260), .IN2(r802_n261), .QN(r802_n254) );
  NAND2X0 r802_U266 ( .IN1(r802_n259), .IN2(r802_n254), .QN(r802_n257) );
  OR2X1 r802_U265 ( .IN2(r802_n254), .IN1(r802_n259), .Q(r802_n258) );
  NAND2X0 r802_U264 ( .IN1(r802_n257), .IN2(r802_n258), .QN(P1_N2893) );
  INVX0 r802_U263 ( .ZN(r802_n243), .INP(P1_N2742) );
  NAND2X0 r802_U262 ( .IN1(P1_N5160), .IN2(r802_n243), .QN(r802_n255) );
  OR2X1 r802_U261 ( .IN2(P1_N5160), .IN1(r802_n243), .Q(r802_n256) );
  NAND2X0 r802_U260 ( .IN1(r802_n255), .IN2(r802_n256), .QN(r802_n249) );
  NAND2X0 r802_U259 ( .IN1(n7066), .IN2(r802_n254), .QN(r802_n250) );
  OR2X1 r802_U258 ( .IN2(n7066), .IN1(r802_n254), .Q(r802_n252) );
  NAND2X0 r802_U257 ( .IN1(r802_n252), .IN2(r802_n253), .QN(r802_n251) );
  NAND2X0 r802_U256 ( .IN1(r802_n250), .IN2(r802_n251), .QN(r802_n244) );
  NAND2X0 r802_U255 ( .IN1(r802_n249), .IN2(r802_n244), .QN(r802_n247) );
  OR2X1 r802_U254 ( .IN2(r802_n244), .IN1(r802_n249), .Q(r802_n248) );
  NAND2X0 r802_U253 ( .IN1(r802_n247), .IN2(r802_n248), .QN(P1_N2894) );
  INVX0 r802_U252 ( .ZN(r802_n233), .INP(P1_N2743) );
  NAND2X0 r802_U251 ( .IN1(P1_N5161), .IN2(r802_n233), .QN(r802_n245) );
  OR2X1 r802_U250 ( .IN2(P1_N5161), .IN1(r802_n233), .Q(r802_n246) );
  NAND2X0 r802_U249 ( .IN1(r802_n245), .IN2(r802_n246), .QN(r802_n239) );
  NAND2X0 r802_U248 ( .IN1(P1_N5160), .IN2(r802_n244), .QN(r802_n240) );
  OR2X1 r802_U247 ( .IN2(P1_N5160), .IN1(r802_n244), .Q(r802_n242) );
  NAND2X0 r802_U246 ( .IN1(r802_n242), .IN2(r802_n243), .QN(r802_n241) );
  NAND2X0 r802_U245 ( .IN1(r802_n240), .IN2(r802_n241), .QN(r802_n234) );
  NAND2X0 r802_U244 ( .IN1(r802_n239), .IN2(r802_n234), .QN(r802_n237) );
  OR2X1 r802_U243 ( .IN2(r802_n234), .IN1(r802_n239), .Q(r802_n238) );
  NAND2X0 r802_U242 ( .IN1(r802_n237), .IN2(r802_n238), .QN(P1_N2895) );
  INVX0 r802_U241 ( .ZN(r802_n223), .INP(P1_N2744) );
  NAND2X0 r802_U240 ( .IN1(P1_N5162), .IN2(r802_n223), .QN(r802_n235) );
  OR2X1 r802_U239 ( .IN2(P1_N5162), .IN1(r802_n223), .Q(r802_n236) );
  NAND2X0 r802_U238 ( .IN1(r802_n235), .IN2(r802_n236), .QN(r802_n229) );
  NAND2X0 r802_U237 ( .IN1(P1_N5161), .IN2(r802_n234), .QN(r802_n230) );
  OR2X1 r802_U236 ( .IN2(P1_N5161), .IN1(r802_n234), .Q(r802_n232) );
  NAND2X0 r802_U235 ( .IN1(r802_n232), .IN2(r802_n233), .QN(r802_n231) );
  NAND2X0 r802_U234 ( .IN1(r802_n230), .IN2(r802_n231), .QN(r802_n224) );
  OR2X1 r804_U88 ( .IN2(P1_N5175), .IN1(r804_n87), .Q(r804_n86) );
  NAND2X0 r804_U87 ( .IN1(P1_N3130), .IN2(r804_n86), .QN(r804_n85) );
  NAND2X0 r804_U86 ( .IN1(r804_n84), .IN2(r804_n85), .QN(r804_n77) );
  OR2X1 r804_U84 ( .IN2(P1_N3131), .IN1(n7119), .Q(r804_n81) );
  NAND2X0 r804_U83 ( .IN1(P1_N3131), .IN2(n7119), .QN(r804_n82) );
  NAND2X0 r804_U82 ( .IN1(r804_n81), .IN2(r804_n82), .QN(r804_n80) );
  NOR2X0 r804_U81 ( .QN(r804_n78), .IN1(r804_n77), .IN2(r804_n80) );
  AND2X1 r804_U80 ( .IN1(r804_n77), .IN2(r804_n80), .Q(r804_n79) );
  NOR2X0 r804_U79 ( .QN(P1_N3283), .IN1(r804_n78), .IN2(r804_n79) );
  NAND2X0 r804_U78 ( .IN1(n7122), .IN2(r804_n77), .QN(r804_n74) );
  OR2X1 r804_U77 ( .IN2(n7122), .IN1(r804_n77), .Q(r804_n76) );
  NAND2X0 r804_U76 ( .IN1(P1_N3131), .IN2(r804_n76), .QN(r804_n75) );
  NAND2X0 r804_U75 ( .IN1(r804_n74), .IN2(r804_n75), .QN(r804_n64) );
  OR2X1 r804_U73 ( .IN2(P1_N3132), .IN1(n7117), .Q(r804_n71) );
  NAND2X0 r804_U72 ( .IN1(P1_N3132), .IN2(n7117), .QN(r804_n72) );
  NAND2X0 r804_U71 ( .IN1(r804_n71), .IN2(r804_n72), .QN(r804_n70) );
  NOR2X0 r804_U70 ( .QN(r804_n68), .IN1(r804_n64), .IN2(r804_n70) );
  AND2X1 r804_U69 ( .IN1(r804_n64), .IN2(r804_n70), .Q(r804_n69) );
  NOR2X0 r804_U68 ( .QN(P1_N3284), .IN1(r804_n68), .IN2(r804_n69) );
  OR2X1 r804_U66 ( .IN2(P1_N3133), .IN1(n7146), .Q(r804_n65) );
  NAND2X0 r804_U65 ( .IN1(P1_N3133), .IN2(n7146), .QN(r804_n66) );
  NAND2X0 r804_U64 ( .IN1(r804_n65), .IN2(r804_n66), .QN(r804_n60) );
  NAND2X0 r804_U63 ( .IN1(P1_N5177), .IN2(r804_n64), .QN(r804_n61) );
  OR2X1 r804_U62 ( .IN2(P1_N5177), .IN1(r804_n64), .Q(r804_n63) );
  NAND2X0 r804_U61 ( .IN1(P1_N3132), .IN2(r804_n63), .QN(r804_n62) );
  NAND2X0 r804_U60 ( .IN1(r804_n61), .IN2(r804_n62), .QN(r804_n59) );
  NOR2X0 r804_U59 ( .QN(r804_n57), .IN1(r804_n60), .IN2(r804_n59) );
  AND2X1 r804_U58 ( .IN1(r804_n59), .IN2(r804_n60), .Q(r804_n58) );
  NOR2X0 r804_U57 ( .QN(P1_N3285), .IN1(r804_n57), .IN2(r804_n58) );
  OR2X1 r804_U55 ( .IN2(P1_N3106), .IN1(n7045), .Q(r804_n54) );
  NAND2X0 r804_U54 ( .IN1(P1_N3106), .IN2(n7045), .QN(r804_n55) );
  NAND2X0 r804_U53 ( .IN1(r804_n54), .IN2(r804_n55), .QN(r804_n53) );
  NOR2X0 r804_U52 ( .QN(r804_n50), .IN1(r804_n52), .IN2(r804_n53) );
  AND2X1 r804_U51 ( .IN1(r804_n52), .IN2(r804_n53), .Q(r804_n51) );
  NOR2X0 r804_U50 ( .QN(P1_N3258), .IN1(r804_n50), .IN2(r804_n51) );
  OR2X1 r804_U48 ( .IN2(P1_N3107), .IN1(n7043), .Q(r804_n47) );
  NAND2X0 r804_U47 ( .IN1(P1_N3107), .IN2(n7043), .QN(r804_n48) );
  NAND2X0 r804_U46 ( .IN1(r804_n47), .IN2(r804_n48), .QN(r804_n46) );
  NOR2X0 r804_U45 ( .QN(r804_n43), .IN1(r804_n45), .IN2(r804_n46) );
  AND2X1 r804_U44 ( .IN1(r804_n45), .IN2(r804_n46), .Q(r804_n44) );
  NOR2X0 r804_U43 ( .QN(P1_N3259), .IN1(r804_n43), .IN2(r804_n44) );
  OR2X1 r804_U41 ( .IN2(P1_N3108), .IN1(n7037), .Q(r804_n40) );
  NAND2X0 r804_U40 ( .IN1(P1_N3108), .IN2(n7037), .QN(r804_n41) );
  NAND2X0 r804_U39 ( .IN1(r804_n40), .IN2(r804_n41), .QN(r804_n39) );
  NOR2X0 r804_U38 ( .QN(r804_n36), .IN1(r804_n38), .IN2(r804_n39) );
  AND2X1 r804_U37 ( .IN1(r804_n38), .IN2(r804_n39), .Q(r804_n37) );
  NOR2X0 r804_U36 ( .QN(P1_N3260), .IN1(r804_n36), .IN2(r804_n37) );
  OR2X1 r804_U34 ( .IN2(P1_N3109), .IN1(n7082), .Q(r804_n33) );
  NAND2X0 r804_U33 ( .IN1(P1_N3109), .IN2(n7082), .QN(r804_n34) );
  NAND2X0 r804_U32 ( .IN1(r804_n33), .IN2(r804_n34), .QN(r804_n32) );
  NOR2X0 r804_U31 ( .QN(r804_n29), .IN1(r804_n31), .IN2(r804_n32) );
  AND2X1 r804_U30 ( .IN1(r804_n31), .IN2(r804_n32), .Q(r804_n30) );
  NOR2X0 r804_U29 ( .QN(P1_N3261), .IN1(r804_n29), .IN2(r804_n30) );
  OR2X1 r804_U27 ( .IN2(P1_N3110), .IN1(n7079), .Q(r804_n26) );
  NAND2X0 r804_U26 ( .IN1(P1_N3110), .IN2(n7079), .QN(r804_n27) );
  NAND2X0 r804_U25 ( .IN1(r804_n26), .IN2(r804_n27), .QN(r804_n25) );
  NOR2X0 r804_U24 ( .QN(r804_n22), .IN1(r804_n24), .IN2(r804_n25) );
  AND2X1 r804_U23 ( .IN1(r804_n24), .IN2(r804_n25), .Q(r804_n23) );
  NOR2X0 r804_U22 ( .QN(P1_N3262), .IN1(r804_n22), .IN2(r804_n23) );
  OR2X1 r804_U20 ( .IN2(P1_N3111), .IN1(n7076), .Q(r804_n19) );
  NAND2X0 r804_U19 ( .IN1(P1_N3111), .IN2(n7076), .QN(r804_n20) );
  NAND2X0 r804_U18 ( .IN1(r804_n19), .IN2(r804_n20), .QN(r804_n18) );
  NOR2X0 r804_U17 ( .QN(r804_n15), .IN1(r804_n17), .IN2(r804_n18) );
  AND2X1 r804_U16 ( .IN1(r804_n17), .IN2(r804_n18), .Q(r804_n16) );
  NOR2X0 r804_U15 ( .QN(P1_N3263), .IN1(r804_n15), .IN2(r804_n16) );
  OR2X1 r804_U13 ( .IN2(P1_N3112), .IN1(n7073), .Q(r804_n12) );
  NAND2X0 r804_U12 ( .IN1(P1_N3112), .IN2(n7073), .QN(r804_n13) );
  NAND2X0 r804_U11 ( .IN1(r804_n12), .IN2(r804_n13), .QN(r804_n11) );
  NOR2X0 r804_U10 ( .QN(r804_n8), .IN1(r804_n10), .IN2(r804_n11) );
  AND2X1 r804_U9 ( .IN1(r804_n10), .IN2(r804_n11), .Q(r804_n9) );
  NOR2X0 r804_U8 ( .QN(P1_N3264), .IN1(r804_n8), .IN2(r804_n9) );
  OR2X1 r804_U6 ( .IN2(P1_N3113), .IN1(n7071), .Q(r804_n5) );
  NAND2X0 r804_U5 ( .IN1(P1_N3113), .IN2(n7071), .QN(r804_n6) );
  NAND2X0 r804_U4 ( .IN1(r804_n5), .IN2(r804_n6), .QN(r804_n4) );
  NOR2X0 r804_U3 ( .QN(r804_n1), .IN1(r804_n3), .IN2(r804_n4) );
  AND2X1 r804_U2 ( .IN1(r804_n3), .IN2(r804_n4), .Q(r804_n2) );
  NOR2X0 r804_U1 ( .QN(P1_N3265), .IN1(r804_n1), .IN2(r804_n2) );
  NAND2X0 r804_U181 ( .IN1(P1_N3122), .IN2(r804_n173), .QN(r804_n172) );
  NAND2X0 r804_U180 ( .IN1(r804_n171), .IN2(r804_n172), .QN(r804_n157) );
  OR2X1 r804_U178 ( .IN2(P1_N3123), .IN1(n7098), .Q(r804_n168) );
  NAND2X0 r804_U177 ( .IN1(P1_N3123), .IN2(n7098), .QN(r804_n169) );
  NAND2X0 r804_U176 ( .IN1(r804_n168), .IN2(r804_n169), .QN(r804_n167) );
  NOR2X0 r804_U175 ( .QN(r804_n165), .IN1(r804_n157), .IN2(r804_n167) );
  AND2X1 r804_U174 ( .IN1(r804_n157), .IN2(r804_n167), .Q(r804_n166) );
  NOR2X0 r804_U173 ( .QN(P1_N3275), .IN1(r804_n165), .IN2(r804_n166) );
  OR2X1 r804_U172 ( .IN2(P1_N3105), .IN1(n7051), .Q(r804_n162) );
  NAND2X0 r804_U171 ( .IN1(P1_N3105), .IN2(n7051), .QN(r804_n163) );
  NAND2X0 r804_U170 ( .IN1(r804_n162), .IN2(r804_n163), .QN(r804_n160) );
  NAND2X0 r804_U169 ( .IN1(r804_n160), .IN2(r804_n161), .QN(r804_n158) );
  OR2X1 r804_U168 ( .IN2(r804_n161), .IN1(r804_n160), .Q(r804_n159) );
  NAND2X0 r804_U167 ( .IN1(r804_n158), .IN2(r804_n159), .QN(P1_N3257) );
  NAND2X0 r804_U166 ( .IN1(n7099), .IN2(r804_n157), .QN(r804_n154) );
  OR2X1 r804_U165 ( .IN2(n7099), .IN1(r804_n157), .Q(r804_n156) );
  NAND2X0 r804_U164 ( .IN1(P1_N3123), .IN2(r804_n156), .QN(r804_n155) );
  NAND2X0 r804_U163 ( .IN1(r804_n154), .IN2(r804_n155), .QN(r804_n147) );
  OR2X1 r804_U161 ( .IN2(P1_N3124), .IN1(n7095), .Q(r804_n151) );
  NAND2X0 r804_U160 ( .IN1(P1_N3124), .IN2(n7095), .QN(r804_n152) );
  NAND2X0 r804_U159 ( .IN1(r804_n151), .IN2(r804_n152), .QN(r804_n150) );
  NOR2X0 r804_U158 ( .QN(r804_n148), .IN1(r804_n147), .IN2(r804_n150) );
  AND2X1 r804_U157 ( .IN1(r804_n147), .IN2(r804_n150), .Q(r804_n149) );
  NOR2X0 r804_U156 ( .QN(P1_N3276), .IN1(r804_n148), .IN2(r804_n149) );
  NAND2X0 r804_U155 ( .IN1(P1_N5169), .IN2(r804_n147), .QN(r804_n144) );
  OR2X1 r804_U154 ( .IN2(P1_N5169), .IN1(r804_n147), .Q(r804_n146) );
  NAND2X0 r804_U153 ( .IN1(P1_N3124), .IN2(r804_n146), .QN(r804_n145) );
  NAND2X0 r804_U152 ( .IN1(r804_n144), .IN2(r804_n145), .QN(r804_n137) );
  OR2X1 r804_U150 ( .IN2(P1_N3125), .IN1(n7092), .Q(r804_n141) );
  NAND2X0 r804_U149 ( .IN1(P1_N3125), .IN2(n7092), .QN(r804_n142) );
  NAND2X0 r804_U148 ( .IN1(r804_n141), .IN2(r804_n142), .QN(r804_n140) );
  NOR2X0 r804_U147 ( .QN(r804_n138), .IN1(r804_n137), .IN2(r804_n140) );
  AND2X1 r804_U146 ( .IN1(r804_n137), .IN2(r804_n140), .Q(r804_n139) );
  NOR2X0 r804_U145 ( .QN(P1_N3277), .IN1(r804_n138), .IN2(r804_n139) );
  NAND2X0 r804_U144 ( .IN1(P1_N5170), .IN2(r804_n137), .QN(r804_n134) );
  OR2X1 r804_U143 ( .IN2(P1_N5170), .IN1(r804_n137), .Q(r804_n136) );
  NAND2X0 r804_U142 ( .IN1(P1_N3125), .IN2(r804_n136), .QN(r804_n135) );
  NAND2X0 r804_U141 ( .IN1(r804_n134), .IN2(r804_n135), .QN(r804_n127) );
  OR2X1 r804_U139 ( .IN2(P1_N3126), .IN1(n7090), .Q(r804_n131) );
  NAND2X0 r804_U138 ( .IN1(P1_N3126), .IN2(n7090), .QN(r804_n132) );
  NAND2X0 r804_U137 ( .IN1(r804_n131), .IN2(r804_n132), .QN(r804_n130) );
  NOR2X0 r804_U136 ( .QN(r804_n128), .IN1(r804_n127), .IN2(r804_n130) );
  AND2X1 r804_U135 ( .IN1(r804_n127), .IN2(r804_n130), .Q(r804_n129) );
  NOR2X0 r804_U134 ( .QN(P1_N3278), .IN1(r804_n128), .IN2(r804_n129) );
  NAND2X0 r804_U133 ( .IN1(n7089), .IN2(r804_n127), .QN(r804_n124) );
  OR2X1 r804_U132 ( .IN2(n7089), .IN1(r804_n127), .Q(r804_n126) );
  NAND2X0 r804_U131 ( .IN1(P1_N3126), .IN2(r804_n126), .QN(r804_n125) );
  NAND2X0 r804_U130 ( .IN1(r804_n124), .IN2(r804_n125), .QN(r804_n117) );
  OR2X1 r804_U128 ( .IN2(P1_N3127), .IN1(n7144), .Q(r804_n121) );
  NAND2X0 r804_U127 ( .IN1(P1_N3127), .IN2(n7144), .QN(r804_n122) );
  NAND2X0 r804_U126 ( .IN1(r804_n121), .IN2(r804_n122), .QN(r804_n120) );
  NOR2X0 r804_U125 ( .QN(r804_n118), .IN1(r804_n117), .IN2(r804_n120) );
  AND2X1 r804_U124 ( .IN1(r804_n117), .IN2(r804_n120), .Q(r804_n119) );
  NOR2X0 r804_U123 ( .QN(P1_N3279), .IN1(r804_n118), .IN2(r804_n119) );
  NAND2X0 r804_U122 ( .IN1(n7141), .IN2(r804_n117), .QN(r804_n114) );
  OR2X1 r804_U121 ( .IN2(n7141), .IN1(r804_n117), .Q(r804_n116) );
  NAND2X0 r804_U120 ( .IN1(P1_N3127), .IN2(r804_n116), .QN(r804_n115) );
  NAND2X0 r804_U119 ( .IN1(r804_n114), .IN2(r804_n115), .QN(r804_n107) );
  OR2X1 r804_U117 ( .IN2(P1_N3128), .IN1(n7136), .Q(r804_n111) );
  NAND2X0 r804_U116 ( .IN1(P1_N3128), .IN2(n7136), .QN(r804_n112) );
  NAND2X0 r804_U115 ( .IN1(r804_n111), .IN2(r804_n112), .QN(r804_n110) );
  NOR2X0 r804_U114 ( .QN(r804_n108), .IN1(r804_n107), .IN2(r804_n110) );
  AND2X1 r804_U113 ( .IN1(r804_n107), .IN2(r804_n110), .Q(r804_n109) );
  NOR2X0 r804_U112 ( .QN(P1_N3280), .IN1(r804_n108), .IN2(r804_n109) );
  NAND2X0 r804_U111 ( .IN1(P1_N5173), .IN2(r804_n107), .QN(r804_n104) );
  OR2X1 r804_U110 ( .IN2(P1_N5173), .IN1(r804_n107), .Q(r804_n106) );
  NAND2X0 r804_U109 ( .IN1(P1_N3128), .IN2(r804_n106), .QN(r804_n105) );
  NAND2X0 r804_U108 ( .IN1(r804_n104), .IN2(r804_n105), .QN(r804_n97) );
  OR2X1 r804_U106 ( .IN2(P1_N3129), .IN1(n7130), .Q(r804_n101) );
  NAND2X0 r804_U105 ( .IN1(P1_N3129), .IN2(n7130), .QN(r804_n102) );
  NAND2X0 r804_U104 ( .IN1(r804_n101), .IN2(r804_n102), .QN(r804_n100) );
  NOR2X0 r804_U103 ( .QN(r804_n98), .IN1(r804_n97), .IN2(r804_n100) );
  AND2X1 r804_U102 ( .IN1(r804_n97), .IN2(r804_n100), .Q(r804_n99) );
  NOR2X0 r804_U101 ( .QN(P1_N3281), .IN1(r804_n98), .IN2(r804_n99) );
  NAND2X0 r804_U100 ( .IN1(n7129), .IN2(r804_n97), .QN(r804_n94) );
  OR2X1 r804_U99 ( .IN2(n7129), .IN1(r804_n97), .Q(r804_n96) );
  NAND2X0 r804_U98 ( .IN1(P1_N3129), .IN2(r804_n96), .QN(r804_n95) );
  NAND2X0 r804_U97 ( .IN1(r804_n94), .IN2(r804_n95), .QN(r804_n87) );
  OR2X1 r804_U95 ( .IN2(P1_N3130), .IN1(n7125), .Q(r804_n91) );
  NAND2X0 r804_U94 ( .IN1(P1_N3130), .IN2(n7125), .QN(r804_n92) );
  NAND2X0 r804_U93 ( .IN1(r804_n91), .IN2(r804_n92), .QN(r804_n90) );
  NOR2X0 r804_U92 ( .QN(r804_n88), .IN1(r804_n87), .IN2(r804_n90) );
  AND2X1 r804_U91 ( .IN1(r804_n87), .IN2(r804_n90), .Q(r804_n89) );
  NOR2X0 r804_U90 ( .QN(P1_N3282), .IN1(r804_n88), .IN2(r804_n89) );
  NAND2X0 r804_U89 ( .IN1(P1_N5175), .IN2(r804_n87), .QN(r804_n84) );
  NOR2X0 r804_U274 ( .QN(r804_n255), .IN1(r804_n254), .IN2(r804_n257) );
  AND2X1 r804_U273 ( .IN1(r804_n254), .IN2(r804_n257), .Q(r804_n256) );
  NOR2X0 r804_U272 ( .QN(P1_N3266), .IN1(r804_n255), .IN2(r804_n256) );
  NAND2X0 r804_U271 ( .IN1(P1_N5159), .IN2(r804_n254), .QN(r804_n251) );
  OR2X1 r804_U270 ( .IN2(P1_N5159), .IN1(r804_n254), .Q(r804_n253) );
  NAND2X0 r804_U269 ( .IN1(P1_N3114), .IN2(r804_n253), .QN(r804_n252) );
  NAND2X0 r804_U268 ( .IN1(r804_n251), .IN2(r804_n252), .QN(r804_n244) );
  OR2X1 r804_U266 ( .IN2(P1_N3115), .IN1(n7063), .Q(r804_n248) );
  NAND2X0 r804_U265 ( .IN1(P1_N3115), .IN2(n7063), .QN(r804_n249) );
  NAND2X0 r804_U264 ( .IN1(r804_n248), .IN2(r804_n249), .QN(r804_n247) );
  NOR2X0 r804_U263 ( .QN(r804_n245), .IN1(r804_n244), .IN2(r804_n247) );
  AND2X1 r804_U262 ( .IN1(r804_n244), .IN2(r804_n247), .Q(r804_n246) );
  NOR2X0 r804_U261 ( .QN(P1_N3267), .IN1(r804_n245), .IN2(r804_n246) );
  NAND2X0 r804_U260 ( .IN1(P1_N5160), .IN2(r804_n244), .QN(r804_n241) );
  OR2X1 r804_U259 ( .IN2(P1_N5160), .IN1(r804_n244), .Q(r804_n243) );
  NAND2X0 r804_U258 ( .IN1(P1_N3115), .IN2(r804_n243), .QN(r804_n242) );
  NAND2X0 r804_U257 ( .IN1(r804_n241), .IN2(r804_n242), .QN(r804_n234) );
  OR2X1 r804_U255 ( .IN2(P1_N3116), .IN1(n7058), .Q(r804_n238) );
  NAND2X0 r804_U254 ( .IN1(P1_N3116), .IN2(n7058), .QN(r804_n239) );
  NAND2X0 r804_U253 ( .IN1(r804_n238), .IN2(r804_n239), .QN(r804_n237) );
  NOR2X0 r804_U252 ( .QN(r804_n235), .IN1(r804_n234), .IN2(r804_n237) );
  AND2X1 r804_U251 ( .IN1(r804_n234), .IN2(r804_n237), .Q(r804_n236) );
  NOR2X0 r804_U250 ( .QN(P1_N3268), .IN1(r804_n235), .IN2(r804_n236) );
  NAND2X0 r804_U249 ( .IN1(P1_N5161), .IN2(r804_n234), .QN(r804_n231) );
  OR2X1 r804_U248 ( .IN2(P1_N5161), .IN1(r804_n234), .Q(r804_n233) );
  NAND2X0 r804_U247 ( .IN1(P1_N3116), .IN2(r804_n233), .QN(r804_n232) );
  NAND2X0 r804_U246 ( .IN1(r804_n231), .IN2(r804_n232), .QN(r804_n224) );
  OR2X1 r804_U244 ( .IN2(P1_N3117), .IN1(n7056), .Q(r804_n228) );
  NAND2X0 r804_U243 ( .IN1(P1_N3117), .IN2(n7056), .QN(r804_n229) );
  NAND2X0 r804_U242 ( .IN1(r804_n228), .IN2(r804_n229), .QN(r804_n227) );
  NOR2X0 r804_U241 ( .QN(r804_n225), .IN1(r804_n224), .IN2(r804_n227) );
  AND2X1 r804_U240 ( .IN1(r804_n224), .IN2(r804_n227), .Q(r804_n226) );
  NOR2X0 r804_U239 ( .QN(P1_N3269), .IN1(r804_n225), .IN2(r804_n226) );
  NAND2X0 r804_U238 ( .IN1(P1_N5162), .IN2(r804_n224), .QN(r804_n221) );
  OR2X1 r804_U237 ( .IN2(P1_N5162), .IN1(r804_n224), .Q(r804_n223) );
  NAND2X0 r804_U236 ( .IN1(P1_N3117), .IN2(r804_n223), .QN(r804_n222) );
  NAND2X0 r804_U235 ( .IN1(r804_n221), .IN2(r804_n222), .QN(r804_n214) );
  OR2X1 r804_U233 ( .IN2(P1_N3118), .IN1(n7115), .Q(r804_n218) );
  NAND2X0 r804_U232 ( .IN1(P1_N3118), .IN2(n7115), .QN(r804_n219) );
  NAND2X0 r804_U231 ( .IN1(r804_n218), .IN2(r804_n219), .QN(r804_n217) );
  NOR2X0 r804_U230 ( .QN(r804_n215), .IN1(r804_n214), .IN2(r804_n217) );
  AND2X1 r804_U229 ( .IN1(r804_n214), .IN2(r804_n217), .Q(r804_n216) );
  NOR2X0 r804_U228 ( .QN(P1_N3270), .IN1(r804_n215), .IN2(r804_n216) );
  NAND2X0 r804_U227 ( .IN1(P1_N5163), .IN2(r804_n214), .QN(r804_n211) );
  OR2X1 r804_U226 ( .IN2(P1_N5163), .IN1(r804_n214), .Q(r804_n213) );
  NAND2X0 r804_U225 ( .IN1(P1_N3118), .IN2(r804_n213), .QN(r804_n212) );
  NAND2X0 r804_U224 ( .IN1(r804_n211), .IN2(r804_n212), .QN(r804_n204) );
  OR2X1 r804_U222 ( .IN2(P1_N3119), .IN1(n7112), .Q(r804_n208) );
  NAND2X0 r804_U221 ( .IN1(P1_N3119), .IN2(n7112), .QN(r804_n209) );
  NAND2X0 r804_U220 ( .IN1(r804_n208), .IN2(r804_n209), .QN(r804_n207) );
  NOR2X0 r804_U219 ( .QN(r804_n205), .IN1(r804_n204), .IN2(r804_n207) );
  AND2X1 r804_U218 ( .IN1(r804_n204), .IN2(r804_n207), .Q(r804_n206) );
  NOR2X0 r804_U217 ( .QN(P1_N3271), .IN1(r804_n205), .IN2(r804_n206) );
  NAND2X0 r804_U216 ( .IN1(P1_N5164), .IN2(r804_n204), .QN(r804_n201) );
  OR2X1 r804_U215 ( .IN2(P1_N5164), .IN1(r804_n204), .Q(r804_n203) );
  NAND2X0 r804_U214 ( .IN1(P1_N3119), .IN2(r804_n203), .QN(r804_n202) );
  NAND2X0 r804_U213 ( .IN1(r804_n201), .IN2(r804_n202), .QN(r804_n194) );
  OR2X1 r804_U211 ( .IN2(P1_N3120), .IN1(n7109), .Q(r804_n198) );
  NAND2X0 r804_U210 ( .IN1(P1_N3120), .IN2(n7109), .QN(r804_n199) );
  NAND2X0 r804_U209 ( .IN1(r804_n198), .IN2(r804_n199), .QN(r804_n197) );
  NOR2X0 r804_U208 ( .QN(r804_n195), .IN1(r804_n194), .IN2(r804_n197) );
  AND2X1 r804_U207 ( .IN1(r804_n194), .IN2(r804_n197), .Q(r804_n196) );
  NOR2X0 r804_U206 ( .QN(P1_N3272), .IN1(r804_n195), .IN2(r804_n196) );
  NAND2X0 r804_U205 ( .IN1(P1_N5165), .IN2(r804_n194), .QN(r804_n191) );
  OR2X1 r804_U204 ( .IN2(P1_N5165), .IN1(r804_n194), .Q(r804_n193) );
  NAND2X0 r804_U203 ( .IN1(P1_N3120), .IN2(r804_n193), .QN(r804_n192) );
  NAND2X0 r804_U202 ( .IN1(r804_n191), .IN2(r804_n192), .QN(r804_n184) );
  OR2X1 r804_U200 ( .IN2(P1_N3121), .IN1(n7105), .Q(r804_n188) );
  NAND2X0 r804_U199 ( .IN1(P1_N3121), .IN2(n7105), .QN(r804_n189) );
  NAND2X0 r804_U198 ( .IN1(r804_n188), .IN2(r804_n189), .QN(r804_n187) );
  NOR2X0 r804_U197 ( .QN(r804_n185), .IN1(r804_n184), .IN2(r804_n187) );
  AND2X1 r804_U196 ( .IN1(r804_n184), .IN2(r804_n187), .Q(r804_n186) );
  NOR2X0 r804_U195 ( .QN(P1_N3273), .IN1(r804_n185), .IN2(r804_n186) );
  NAND2X0 r804_U194 ( .IN1(n7106), .IN2(r804_n184), .QN(r804_n181) );
  OR2X1 r804_U193 ( .IN2(n7106), .IN1(r804_n184), .Q(r804_n183) );
  NAND2X0 r804_U192 ( .IN1(P1_N3121), .IN2(r804_n183), .QN(r804_n182) );
  NAND2X0 r804_U191 ( .IN1(r804_n181), .IN2(r804_n182), .QN(r804_n174) );
  OR2X1 r804_U189 ( .IN2(P1_N3122), .IN1(n7102), .Q(r804_n178) );
  NAND2X0 r804_U188 ( .IN1(P1_N3122), .IN2(n7102), .QN(r804_n179) );
  NAND2X0 r804_U187 ( .IN1(r804_n178), .IN2(r804_n179), .QN(r804_n177) );
  NOR2X0 r804_U186 ( .QN(r804_n175), .IN1(r804_n174), .IN2(r804_n177) );
  AND2X1 r804_U185 ( .IN1(r804_n174), .IN2(r804_n177), .Q(r804_n176) );
  NOR2X0 r804_U184 ( .QN(P1_N3274), .IN1(r804_n175), .IN2(r804_n176) );
  NAND2X0 r804_U183 ( .IN1(P1_N5167), .IN2(r804_n174), .QN(r804_n171) );
  OR2X1 r804_U182 ( .IN2(P1_N5167), .IN1(r804_n174), .Q(r804_n173) );
  OR2X1 r804_U319 ( .IN2(P1_N3104), .IN1(n4803), .Q(r804_n288) );
  NAND2X0 r804_U318 ( .IN1(P1_N3104), .IN2(n4803), .QN(r804_n289) );
  NAND2X0 r804_U317 ( .IN1(r804_n288), .IN2(r804_n289), .QN(P1_N3256) );
  NAND2X0 r804_U315 ( .IN1(P1_N3104), .IN2(n7034), .QN(r804_n161) );
  OR2X1 r804_U314 ( .IN2(r804_n161), .IN1(n7051), .Q(r804_n285) );
  NAND2X0 r804_U313 ( .IN1(n7051), .IN2(r804_n161), .QN(r804_n287) );
  NAND2X0 r804_U312 ( .IN1(P1_N3105), .IN2(r804_n287), .QN(r804_n286) );
  NAND2X0 r804_U311 ( .IN1(r804_n285), .IN2(r804_n286), .QN(r804_n52) );
  NAND2X0 r804_U310 ( .IN1(P1_N5151), .IN2(r804_n52), .QN(r804_n282) );
  OR2X1 r804_U309 ( .IN2(P1_N5151), .IN1(r804_n52), .Q(r804_n284) );
  NAND2X0 r804_U308 ( .IN1(P1_N3106), .IN2(r804_n284), .QN(r804_n283) );
  NAND2X0 r804_U307 ( .IN1(r804_n282), .IN2(r804_n283), .QN(r804_n45) );
  NAND2X0 r804_U306 ( .IN1(n7041), .IN2(r804_n45), .QN(r804_n279) );
  OR2X1 r804_U305 ( .IN2(n7041), .IN1(r804_n45), .Q(r804_n281) );
  NAND2X0 r804_U304 ( .IN1(P1_N3107), .IN2(r804_n281), .QN(r804_n280) );
  NAND2X0 r804_U303 ( .IN1(r804_n279), .IN2(r804_n280), .QN(r804_n38) );
  NAND2X0 r804_U302 ( .IN1(n7036), .IN2(r804_n38), .QN(r804_n276) );
  OR2X1 r804_U301 ( .IN2(n7036), .IN1(r804_n38), .Q(r804_n278) );
  NAND2X0 r804_U300 ( .IN1(P1_N3108), .IN2(r804_n278), .QN(r804_n277) );
  NAND2X0 r804_U299 ( .IN1(r804_n276), .IN2(r804_n277), .QN(r804_n31) );
  NAND2X0 r804_U298 ( .IN1(P1_N5154), .IN2(r804_n31), .QN(r804_n273) );
  OR2X1 r804_U297 ( .IN2(P1_N5154), .IN1(r804_n31), .Q(r804_n275) );
  NAND2X0 r804_U296 ( .IN1(P1_N3109), .IN2(r804_n275), .QN(r804_n274) );
  NAND2X0 r804_U295 ( .IN1(r804_n273), .IN2(r804_n274), .QN(r804_n24) );
  NAND2X0 r804_U294 ( .IN1(P1_N5155), .IN2(r804_n24), .QN(r804_n270) );
  OR2X1 r804_U293 ( .IN2(P1_N5155), .IN1(r804_n24), .Q(r804_n272) );
  NAND2X0 r804_U292 ( .IN1(P1_N3110), .IN2(r804_n272), .QN(r804_n271) );
  NAND2X0 r804_U291 ( .IN1(r804_n270), .IN2(r804_n271), .QN(r804_n17) );
  NAND2X0 r804_U290 ( .IN1(n7075), .IN2(r804_n17), .QN(r804_n267) );
  OR2X1 r804_U289 ( .IN2(n7075), .IN1(r804_n17), .Q(r804_n269) );
  NAND2X0 r804_U288 ( .IN1(P1_N3111), .IN2(r804_n269), .QN(r804_n268) );
  NAND2X0 r804_U287 ( .IN1(r804_n267), .IN2(r804_n268), .QN(r804_n10) );
  NAND2X0 r804_U286 ( .IN1(n7072), .IN2(r804_n10), .QN(r804_n264) );
  OR2X1 r804_U285 ( .IN2(n7072), .IN1(r804_n10), .Q(r804_n266) );
  NAND2X0 r804_U284 ( .IN1(P1_N3112), .IN2(r804_n266), .QN(r804_n265) );
  NAND2X0 r804_U283 ( .IN1(r804_n264), .IN2(r804_n265), .QN(r804_n3) );
  NAND2X0 r804_U282 ( .IN1(P1_N5158), .IN2(r804_n3), .QN(r804_n261) );
  OR2X1 r804_U281 ( .IN2(P1_N5158), .IN1(r804_n3), .Q(r804_n263) );
  NAND2X0 r804_U280 ( .IN1(P1_N3113), .IN2(r804_n263), .QN(r804_n262) );
  NAND2X0 r804_U279 ( .IN1(r804_n261), .IN2(r804_n262), .QN(r804_n254) );
  OR2X1 r804_U277 ( .IN2(P1_N3114), .IN1(n7067), .Q(r804_n258) );
  NAND2X0 r804_U276 ( .IN1(P1_N3114), .IN2(n7067), .QN(r804_n259) );
  NAND2X0 r804_U275 ( .IN1(r804_n258), .IN2(r804_n259), .QN(r804_n257) );
  NAND2X0 r806_U37 ( .IN1(r806_n43), .IN2(r806_n44), .QN(P1_N3632) );
  NAND2X0 r806_U36 ( .IN1(P1_N5153), .IN2(r806_n42), .QN(r806_n40) );
  OR2X1 r806_U35 ( .IN2(P1_N5153), .IN1(r806_n42), .Q(r806_n41) );
  NAND2X0 r806_U34 ( .IN1(r806_n40), .IN2(r806_n41), .QN(r806_n38) );
  NAND2X0 r806_U33 ( .IN1(r806_n38), .IN2(r806_n39), .QN(r806_n36) );
  OR2X1 r806_U32 ( .IN2(r806_n39), .IN1(r806_n38), .Q(r806_n37) );
  NAND2X0 r806_U31 ( .IN1(r806_n36), .IN2(r806_n37), .QN(P1_N3633) );
  NAND2X0 r806_U30 ( .IN1(P1_N5154), .IN2(r806_n35), .QN(r806_n33) );
  OR2X1 r806_U29 ( .IN2(P1_N5154), .IN1(r806_n35), .Q(r806_n34) );
  NAND2X0 r806_U28 ( .IN1(r806_n33), .IN2(r806_n34), .QN(r806_n31) );
  NAND2X0 r806_U27 ( .IN1(r806_n31), .IN2(r806_n32), .QN(r806_n29) );
  OR2X1 r806_U26 ( .IN2(r806_n32), .IN1(r806_n31), .Q(r806_n30) );
  NAND2X0 r806_U25 ( .IN1(r806_n29), .IN2(r806_n30), .QN(P1_N3634) );
  NAND2X0 r806_U24 ( .IN1(P1_N5155), .IN2(r806_n28), .QN(r806_n26) );
  OR2X1 r806_U23 ( .IN2(P1_N5155), .IN1(r806_n28), .Q(r806_n27) );
  NAND2X0 r806_U22 ( .IN1(r806_n26), .IN2(r806_n27), .QN(r806_n24) );
  NAND2X0 r806_U21 ( .IN1(r806_n24), .IN2(r806_n25), .QN(r806_n22) );
  OR2X1 r806_U20 ( .IN2(r806_n25), .IN1(r806_n24), .Q(r806_n23) );
  NAND2X0 r806_U19 ( .IN1(r806_n22), .IN2(r806_n23), .QN(P1_N3635) );
  NAND2X0 r806_U18 ( .IN1(n7075), .IN2(r806_n21), .QN(r806_n19) );
  OR2X1 r806_U17 ( .IN2(n7075), .IN1(r806_n21), .Q(r806_n20) );
  NAND2X0 r806_U16 ( .IN1(r806_n19), .IN2(r806_n20), .QN(r806_n17) );
  NAND2X0 r806_U15 ( .IN1(r806_n17), .IN2(r806_n18), .QN(r806_n15) );
  OR2X1 r806_U14 ( .IN2(r806_n18), .IN1(r806_n17), .Q(r806_n16) );
  NAND2X0 r806_U13 ( .IN1(r806_n15), .IN2(r806_n16), .QN(P1_N3636) );
  NAND2X0 r806_U12 ( .IN1(n7072), .IN2(r806_n14), .QN(r806_n12) );
  OR2X1 r806_U11 ( .IN2(n7072), .IN1(r806_n14), .Q(r806_n13) );
  NAND2X0 r806_U10 ( .IN1(r806_n12), .IN2(r806_n13), .QN(r806_n10) );
  NAND2X0 r806_U9 ( .IN1(r806_n10), .IN2(r806_n11), .QN(r806_n8) );
  OR2X1 r806_U8 ( .IN2(r806_n11), .IN1(r806_n10), .Q(r806_n9) );
  NAND2X0 r806_U7 ( .IN1(r806_n8), .IN2(r806_n9), .QN(P1_N3637) );
  NAND2X0 r806_U6 ( .IN1(P1_N5158), .IN2(r806_n7), .QN(r806_n5) );
  OR2X1 r806_U5 ( .IN2(P1_N5158), .IN1(r806_n7), .Q(r806_n6) );
  NAND2X0 r806_U4 ( .IN1(r806_n5), .IN2(r806_n6), .QN(r806_n3) );
  NAND2X0 r806_U3 ( .IN1(r806_n3), .IN2(r806_n4), .QN(r806_n1) );
  OR2X1 r806_U2 ( .IN2(r806_n4), .IN1(r806_n3), .Q(r806_n2) );
  NAND2X0 r806_U1 ( .IN1(r806_n1), .IN2(r806_n2), .QN(P1_N3638) );
  NAND2X0 r806_U130 ( .IN1(r806_n134), .IN2(r806_n135), .QN(r806_n133) );
  NAND2X0 r806_U129 ( .IN1(r806_n132), .IN2(r806_n133), .QN(r806_n126) );
  NAND2X0 r806_U128 ( .IN1(r806_n131), .IN2(r806_n126), .QN(r806_n129) );
  OR2X1 r806_U127 ( .IN2(r806_n126), .IN1(r806_n131), .Q(r806_n130) );
  NAND2X0 r806_U126 ( .IN1(r806_n129), .IN2(r806_n130), .QN(P1_N3651) );
  INVX0 r806_U125 ( .ZN(r806_n115), .INP(P1_N3500) );
  NAND2X0 r806_U124 ( .IN1(P1_N5172), .IN2(r806_n115), .QN(r806_n127) );
  OR2X1 r806_U123 ( .IN2(P1_N5172), .IN1(r806_n115), .Q(r806_n128) );
  NAND2X0 r806_U122 ( .IN1(r806_n127), .IN2(r806_n128), .QN(r806_n121) );
  NAND2X0 r806_U121 ( .IN1(n7089), .IN2(r806_n126), .QN(r806_n122) );
  OR2X1 r806_U120 ( .IN2(n7089), .IN1(r806_n126), .Q(r806_n124) );
  NAND2X0 r806_U119 ( .IN1(r806_n124), .IN2(r806_n125), .QN(r806_n123) );
  NAND2X0 r806_U118 ( .IN1(r806_n122), .IN2(r806_n123), .QN(r806_n116) );
  NAND2X0 r806_U117 ( .IN1(r806_n121), .IN2(r806_n116), .QN(r806_n119) );
  OR2X1 r806_U116 ( .IN2(r806_n116), .IN1(r806_n121), .Q(r806_n120) );
  NAND2X0 r806_U115 ( .IN1(r806_n119), .IN2(r806_n120), .QN(P1_N3652) );
  INVX0 r806_U114 ( .ZN(r806_n105), .INP(P1_N3501) );
  NAND2X0 r806_U113 ( .IN1(n7138), .IN2(r806_n105), .QN(r806_n117) );
  OR2X1 r806_U112 ( .IN2(n7138), .IN1(r806_n105), .Q(r806_n118) );
  NAND2X0 r806_U111 ( .IN1(r806_n117), .IN2(r806_n118), .QN(r806_n111) );
  NAND2X0 r806_U110 ( .IN1(P1_N5172), .IN2(r806_n116), .QN(r806_n112) );
  OR2X1 r806_U109 ( .IN2(P1_N5172), .IN1(r806_n116), .Q(r806_n114) );
  NAND2X0 r806_U108 ( .IN1(r806_n114), .IN2(r806_n115), .QN(r806_n113) );
  NAND2X0 r806_U107 ( .IN1(r806_n112), .IN2(r806_n113), .QN(r806_n106) );
  NAND2X0 r806_U106 ( .IN1(r806_n111), .IN2(r806_n106), .QN(r806_n109) );
  OR2X1 r806_U105 ( .IN2(r806_n106), .IN1(r806_n111), .Q(r806_n110) );
  NAND2X0 r806_U104 ( .IN1(r806_n109), .IN2(r806_n110), .QN(P1_N3653) );
  INVX0 r806_U103 ( .ZN(r806_n95), .INP(P1_N3502) );
  NAND2X0 r806_U102 ( .IN1(n7129), .IN2(r806_n95), .QN(r806_n107) );
  OR2X1 r806_U101 ( .IN2(n7129), .IN1(r806_n95), .Q(r806_n108) );
  NAND2X0 r806_U100 ( .IN1(r806_n107), .IN2(r806_n108), .QN(r806_n101) );
  NAND2X0 r806_U99 ( .IN1(n7138), .IN2(r806_n106), .QN(r806_n102) );
  OR2X1 r806_U98 ( .IN2(n7138), .IN1(r806_n106), .Q(r806_n104) );
  NAND2X0 r806_U97 ( .IN1(r806_n104), .IN2(r806_n105), .QN(r806_n103) );
  NAND2X0 r806_U96 ( .IN1(r806_n102), .IN2(r806_n103), .QN(r806_n96) );
  NAND2X0 r806_U95 ( .IN1(r806_n101), .IN2(r806_n96), .QN(r806_n99) );
  OR2X1 r806_U94 ( .IN2(r806_n96), .IN1(r806_n101), .Q(r806_n100) );
  NAND2X0 r806_U93 ( .IN1(r806_n99), .IN2(r806_n100), .QN(P1_N3654) );
  INVX0 r806_U92 ( .ZN(r806_n85), .INP(P1_N3503) );
  NAND2X0 r806_U91 ( .IN1(n7124), .IN2(r806_n85), .QN(r806_n97) );
  OR2X1 r806_U90 ( .IN2(n7124), .IN1(r806_n85), .Q(r806_n98) );
  NAND2X0 r806_U89 ( .IN1(r806_n97), .IN2(r806_n98), .QN(r806_n91) );
  NAND2X0 r806_U88 ( .IN1(n7129), .IN2(r806_n96), .QN(r806_n92) );
  OR2X1 r806_U87 ( .IN2(n7129), .IN1(r806_n96), .Q(r806_n94) );
  NAND2X0 r806_U86 ( .IN1(r806_n94), .IN2(r806_n95), .QN(r806_n93) );
  NAND2X0 r806_U85 ( .IN1(r806_n92), .IN2(r806_n93), .QN(r806_n86) );
  NAND2X0 r806_U84 ( .IN1(r806_n91), .IN2(r806_n86), .QN(r806_n89) );
  OR2X1 r806_U83 ( .IN2(r806_n86), .IN1(r806_n91), .Q(r806_n90) );
  NAND2X0 r806_U82 ( .IN1(r806_n89), .IN2(r806_n90), .QN(P1_N3655) );
  INVX0 r806_U81 ( .ZN(r806_n75), .INP(P1_N3504) );
  NAND2X0 r806_U80 ( .IN1(n7122), .IN2(r806_n75), .QN(r806_n87) );
  OR2X1 r806_U79 ( .IN2(n7122), .IN1(r806_n75), .Q(r806_n88) );
  NAND2X0 r806_U78 ( .IN1(r806_n87), .IN2(r806_n88), .QN(r806_n81) );
  NAND2X0 r806_U77 ( .IN1(n7124), .IN2(r806_n86), .QN(r806_n82) );
  OR2X1 r806_U76 ( .IN2(n7124), .IN1(r806_n86), .Q(r806_n84) );
  NAND2X0 r806_U75 ( .IN1(r806_n84), .IN2(r806_n85), .QN(r806_n83) );
  NAND2X0 r806_U74 ( .IN1(r806_n82), .IN2(r806_n83), .QN(r806_n76) );
  NAND2X0 r806_U73 ( .IN1(r806_n81), .IN2(r806_n76), .QN(r806_n79) );
  OR2X1 r806_U72 ( .IN2(r806_n76), .IN1(r806_n81), .Q(r806_n80) );
  NAND2X0 r806_U71 ( .IN1(r806_n79), .IN2(r806_n80), .QN(P1_N3656) );
  INVX0 r806_U70 ( .ZN(r806_n64), .INP(P1_N3505) );
  NAND2X0 r806_U69 ( .IN1(P1_N5177), .IN2(r806_n64), .QN(r806_n77) );
  OR2X1 r806_U68 ( .IN2(P1_N5177), .IN1(r806_n64), .Q(r806_n78) );
  NAND2X0 r806_U67 ( .IN1(r806_n77), .IN2(r806_n78), .QN(r806_n71) );
  NAND2X0 r806_U66 ( .IN1(n7122), .IN2(r806_n76), .QN(r806_n72) );
  OR2X1 r806_U65 ( .IN2(n7122), .IN1(r806_n76), .Q(r806_n74) );
  NAND2X0 r806_U64 ( .IN1(r806_n74), .IN2(r806_n75), .QN(r806_n73) );
  NAND2X0 r806_U63 ( .IN1(r806_n72), .IN2(r806_n73), .QN(r806_n65) );
  NAND2X0 r806_U62 ( .IN1(r806_n71), .IN2(r806_n65), .QN(r806_n69) );
  OR2X1 r806_U61 ( .IN2(r806_n65), .IN1(r806_n71), .Q(r806_n70) );
  NAND2X0 r806_U60 ( .IN1(r806_n69), .IN2(r806_n70), .QN(P1_N3657) );
  OR2X1 r806_U58 ( .IN2(P1_N3506), .IN1(n7146), .Q(r806_n66) );
  NAND2X0 r806_U57 ( .IN1(P1_N3506), .IN2(n7146), .QN(r806_n67) );
  NAND2X0 r806_U56 ( .IN1(r806_n66), .IN2(r806_n67), .QN(r806_n60) );
  NAND2X0 r806_U55 ( .IN1(P1_N5177), .IN2(r806_n65), .QN(r806_n61) );
  OR2X1 r806_U54 ( .IN2(P1_N5177), .IN1(r806_n65), .Q(r806_n63) );
  NAND2X0 r806_U53 ( .IN1(r806_n63), .IN2(r806_n64), .QN(r806_n62) );
  NAND2X0 r806_U52 ( .IN1(r806_n61), .IN2(r806_n62), .QN(r806_n59) );
  NAND2X0 r806_U51 ( .IN1(r806_n60), .IN2(r806_n59), .QN(r806_n57) );
  OR2X1 r806_U50 ( .IN2(r806_n60), .IN1(r806_n59), .Q(r806_n58) );
  NAND2X0 r806_U49 ( .IN1(r806_n57), .IN2(r806_n58), .QN(P1_N3658) );
  NAND2X0 r806_U48 ( .IN1(n7046), .IN2(r806_n56), .QN(r806_n54) );
  OR2X1 r806_U47 ( .IN2(n7046), .IN1(r806_n56), .Q(r806_n55) );
  NAND2X0 r806_U46 ( .IN1(r806_n54), .IN2(r806_n55), .QN(r806_n52) );
  NAND2X0 r806_U45 ( .IN1(r806_n52), .IN2(r806_n53), .QN(r806_n50) );
  OR2X1 r806_U44 ( .IN2(r806_n53), .IN1(r806_n52), .Q(r806_n51) );
  NAND2X0 r806_U43 ( .IN1(r806_n50), .IN2(r806_n51), .QN(P1_N3631) );
  NAND2X0 r806_U42 ( .IN1(P1_N5152), .IN2(r806_n49), .QN(r806_n47) );
  OR2X1 r806_U41 ( .IN2(P1_N5152), .IN1(r806_n49), .Q(r806_n48) );
  NAND2X0 r806_U40 ( .IN1(r806_n47), .IN2(r806_n48), .QN(r806_n45) );
  NAND2X0 r806_U39 ( .IN1(r806_n45), .IN2(r806_n46), .QN(r806_n43) );
  OR2X1 r806_U38 ( .IN2(r806_n46), .IN1(r806_n45), .Q(r806_n44) );
  NAND2X0 r806_U223 ( .IN1(r806_n220), .IN2(r806_n221), .QN(r806_n214) );
  NAND2X0 r806_U222 ( .IN1(r806_n219), .IN2(r806_n214), .QN(r806_n217) );
  OR2X1 r806_U221 ( .IN2(r806_n214), .IN1(r806_n219), .Q(r806_n218) );
  NAND2X0 r806_U220 ( .IN1(r806_n217), .IN2(r806_n218), .QN(P1_N3643) );
  INVX0 r806_U219 ( .ZN(r806_n203), .INP(P1_N3492) );
  NAND2X0 r806_U218 ( .IN1(n7113), .IN2(r806_n203), .QN(r806_n215) );
  OR2X1 r806_U217 ( .IN2(n7113), .IN1(r806_n203), .Q(r806_n216) );
  NAND2X0 r806_U216 ( .IN1(r806_n215), .IN2(r806_n216), .QN(r806_n209) );
  NAND2X0 r806_U215 ( .IN1(n7116), .IN2(r806_n214), .QN(r806_n210) );
  OR2X1 r806_U214 ( .IN2(n7116), .IN1(r806_n214), .Q(r806_n212) );
  NAND2X0 r806_U213 ( .IN1(r806_n212), .IN2(r806_n213), .QN(r806_n211) );
  NAND2X0 r806_U212 ( .IN1(r806_n210), .IN2(r806_n211), .QN(r806_n204) );
  NAND2X0 r806_U211 ( .IN1(r806_n209), .IN2(r806_n204), .QN(r806_n207) );
  OR2X1 r806_U210 ( .IN2(r806_n204), .IN1(r806_n209), .Q(r806_n208) );
  NAND2X0 r806_U209 ( .IN1(r806_n207), .IN2(r806_n208), .QN(P1_N3644) );
  INVX0 r806_U208 ( .ZN(r806_n193), .INP(P1_N3493) );
  NAND2X0 r806_U207 ( .IN1(n7110), .IN2(r806_n193), .QN(r806_n205) );
  OR2X1 r806_U206 ( .IN2(n7110), .IN1(r806_n193), .Q(r806_n206) );
  NAND2X0 r806_U205 ( .IN1(r806_n205), .IN2(r806_n206), .QN(r806_n199) );
  NAND2X0 r806_U204 ( .IN1(n7113), .IN2(r806_n204), .QN(r806_n200) );
  OR2X1 r806_U203 ( .IN2(n7113), .IN1(r806_n204), .Q(r806_n202) );
  NAND2X0 r806_U202 ( .IN1(r806_n202), .IN2(r806_n203), .QN(r806_n201) );
  NAND2X0 r806_U201 ( .IN1(r806_n200), .IN2(r806_n201), .QN(r806_n194) );
  NAND2X0 r806_U200 ( .IN1(r806_n199), .IN2(r806_n194), .QN(r806_n197) );
  OR2X1 r806_U199 ( .IN2(r806_n194), .IN1(r806_n199), .Q(r806_n198) );
  NAND2X0 r806_U198 ( .IN1(r806_n197), .IN2(r806_n198), .QN(P1_N3645) );
  INVX0 r806_U197 ( .ZN(r806_n183), .INP(P1_N3494) );
  NAND2X0 r806_U196 ( .IN1(P1_N5166), .IN2(r806_n183), .QN(r806_n195) );
  OR2X1 r806_U195 ( .IN2(P1_N5166), .IN1(r806_n183), .Q(r806_n196) );
  NAND2X0 r806_U194 ( .IN1(r806_n195), .IN2(r806_n196), .QN(r806_n189) );
  NAND2X0 r806_U193 ( .IN1(n7110), .IN2(r806_n194), .QN(r806_n190) );
  OR2X1 r806_U192 ( .IN2(n7110), .IN1(r806_n194), .Q(r806_n192) );
  NAND2X0 r806_U191 ( .IN1(r806_n192), .IN2(r806_n193), .QN(r806_n191) );
  NAND2X0 r806_U190 ( .IN1(r806_n190), .IN2(r806_n191), .QN(r806_n184) );
  NAND2X0 r806_U189 ( .IN1(r806_n189), .IN2(r806_n184), .QN(r806_n187) );
  OR2X1 r806_U188 ( .IN2(r806_n184), .IN1(r806_n189), .Q(r806_n188) );
  NAND2X0 r806_U187 ( .IN1(r806_n187), .IN2(r806_n188), .QN(P1_N3646) );
  INVX0 r806_U186 ( .ZN(r806_n173), .INP(P1_N3495) );
  NAND2X0 r806_U185 ( .IN1(n7103), .IN2(r806_n173), .QN(r806_n185) );
  OR2X1 r806_U184 ( .IN2(n7103), .IN1(r806_n173), .Q(r806_n186) );
  NAND2X0 r806_U183 ( .IN1(r806_n185), .IN2(r806_n186), .QN(r806_n179) );
  NAND2X0 r806_U182 ( .IN1(P1_N5166), .IN2(r806_n184), .QN(r806_n180) );
  OR2X1 r806_U181 ( .IN2(P1_N5166), .IN1(r806_n184), .Q(r806_n182) );
  NAND2X0 r806_U180 ( .IN1(r806_n182), .IN2(r806_n183), .QN(r806_n181) );
  NAND2X0 r806_U179 ( .IN1(r806_n180), .IN2(r806_n181), .QN(r806_n174) );
  NAND2X0 r806_U178 ( .IN1(r806_n179), .IN2(r806_n174), .QN(r806_n177) );
  OR2X1 r806_U177 ( .IN2(r806_n174), .IN1(r806_n179), .Q(r806_n178) );
  NAND2X0 r806_U176 ( .IN1(r806_n177), .IN2(r806_n178), .QN(P1_N3647) );
  INVX0 r806_U175 ( .ZN(r806_n155), .INP(P1_N3496) );
  NAND2X0 r806_U174 ( .IN1(n7099), .IN2(r806_n155), .QN(r806_n175) );
  OR2X1 r806_U173 ( .IN2(n7099), .IN1(r806_n155), .Q(r806_n176) );
  NAND2X0 r806_U172 ( .IN1(r806_n175), .IN2(r806_n176), .QN(r806_n169) );
  NAND2X0 r806_U171 ( .IN1(n7103), .IN2(r806_n174), .QN(r806_n170) );
  OR2X1 r806_U170 ( .IN2(n7103), .IN1(r806_n174), .Q(r806_n172) );
  NAND2X0 r806_U169 ( .IN1(r806_n172), .IN2(r806_n173), .QN(r806_n171) );
  NAND2X0 r806_U168 ( .IN1(r806_n170), .IN2(r806_n171), .QN(r806_n156) );
  NAND2X0 r806_U167 ( .IN1(r806_n169), .IN2(r806_n156), .QN(r806_n167) );
  OR2X1 r806_U166 ( .IN2(r806_n156), .IN1(r806_n169), .Q(r806_n168) );
  NAND2X0 r806_U165 ( .IN1(r806_n167), .IN2(r806_n168), .QN(P1_N3648) );
  NAND2X0 r806_U164 ( .IN1(P1_N5150), .IN2(r806_n166), .QN(r806_n163) );
  NAND2X0 r806_U163 ( .IN1(P1_N3478), .IN2(n7051), .QN(r806_n164) );
  NAND2X0 r806_U162 ( .IN1(r806_n163), .IN2(r806_n164), .QN(r806_n161) );
  NAND2X0 r806_U161 ( .IN1(r806_n161), .IN2(r806_n162), .QN(r806_n159) );
  OR2X1 r806_U160 ( .IN2(r806_n162), .IN1(r806_n161), .Q(r806_n160) );
  NAND2X0 r806_U159 ( .IN1(r806_n159), .IN2(r806_n160), .QN(P1_N3630) );
  INVX0 r806_U158 ( .ZN(r806_n145), .INP(P1_N3497) );
  NAND2X0 r806_U157 ( .IN1(n7096), .IN2(r806_n145), .QN(r806_n157) );
  OR2X1 r806_U156 ( .IN2(P1_N5169), .IN1(r806_n145), .Q(r806_n158) );
  NAND2X0 r806_U155 ( .IN1(r806_n157), .IN2(r806_n158), .QN(r806_n151) );
  NAND2X0 r806_U154 ( .IN1(n7099), .IN2(r806_n156), .QN(r806_n152) );
  OR2X1 r806_U153 ( .IN2(n7099), .IN1(r806_n156), .Q(r806_n154) );
  NAND2X0 r806_U152 ( .IN1(r806_n154), .IN2(r806_n155), .QN(r806_n153) );
  NAND2X0 r806_U151 ( .IN1(r806_n152), .IN2(r806_n153), .QN(r806_n146) );
  NAND2X0 r806_U150 ( .IN1(r806_n151), .IN2(r806_n146), .QN(r806_n149) );
  OR2X1 r806_U149 ( .IN2(r806_n146), .IN1(r806_n151), .Q(r806_n150) );
  NAND2X0 r806_U148 ( .IN1(r806_n149), .IN2(r806_n150), .QN(P1_N3649) );
  INVX0 r806_U147 ( .ZN(r806_n135), .INP(P1_N3498) );
  NAND2X0 r806_U146 ( .IN1(n7093), .IN2(r806_n135), .QN(r806_n147) );
  OR2X1 r806_U145 ( .IN2(n7093), .IN1(r806_n135), .Q(r806_n148) );
  NAND2X0 r806_U144 ( .IN1(r806_n147), .IN2(r806_n148), .QN(r806_n141) );
  NAND2X0 r806_U143 ( .IN1(n7096), .IN2(r806_n146), .QN(r806_n142) );
  OR2X1 r806_U142 ( .IN2(n7096), .IN1(r806_n146), .Q(r806_n144) );
  NAND2X0 r806_U141 ( .IN1(r806_n144), .IN2(r806_n145), .QN(r806_n143) );
  NAND2X0 r806_U140 ( .IN1(r806_n142), .IN2(r806_n143), .QN(r806_n136) );
  NAND2X0 r806_U139 ( .IN1(r806_n141), .IN2(r806_n136), .QN(r806_n139) );
  OR2X1 r806_U138 ( .IN2(r806_n136), .IN1(r806_n141), .Q(r806_n140) );
  NAND2X0 r806_U137 ( .IN1(r806_n139), .IN2(r806_n140), .QN(P1_N3650) );
  INVX0 r806_U136 ( .ZN(r806_n125), .INP(P1_N3499) );
  NAND2X0 r806_U135 ( .IN1(n7089), .IN2(r806_n125), .QN(r806_n137) );
  OR2X1 r806_U134 ( .IN2(n7089), .IN1(r806_n125), .Q(r806_n138) );
  NAND2X0 r806_U133 ( .IN1(r806_n137), .IN2(r806_n138), .QN(r806_n131) );
  NAND2X0 r806_U132 ( .IN1(P1_N5170), .IN2(r806_n136), .QN(r806_n132) );
  OR2X1 r806_U131 ( .IN2(P1_N5170), .IN1(r806_n136), .Q(r806_n134) );
  INVX0 r806_U316 ( .ZN(r806_n253), .INP(P1_N3487) );
  NAND2X0 r806_U315 ( .IN1(P1_N5159), .IN2(r806_n253), .QN(r806_n288) );
  OR2X1 r806_U314 ( .IN2(P1_N5159), .IN1(r806_n253), .Q(r806_n289) );
  NAND2X0 r806_U313 ( .IN1(r806_n288), .IN2(r806_n289), .QN(r806_n259) );
  NAND2X0 r806_U312 ( .IN1(P1_N5150), .IN2(r806_n162), .QN(r806_n284) );
  NAND2X0 r806_U310 ( .IN1(r806_n287), .IN2(n7048), .QN(r806_n286) );
  INVX0 r806_U309 ( .ZN(r806_n166), .INP(P1_N3478) );
  NAND2X0 r806_U308 ( .IN1(r806_n286), .IN2(r806_n166), .QN(r806_n285) );
  NAND2X0 r806_U307 ( .IN1(r806_n284), .IN2(r806_n285), .QN(r806_n53) );
  NAND2X0 r806_U306 ( .IN1(n7046), .IN2(r806_n53), .QN(r806_n281) );
  OR2X1 r806_U305 ( .IN2(n7046), .IN1(r806_n53), .Q(r806_n283) );
  INVX0 r806_U304 ( .ZN(r806_n56), .INP(P1_N3479) );
  NAND2X0 r806_U303 ( .IN1(r806_n283), .IN2(r806_n56), .QN(r806_n282) );
  NAND2X0 r806_U302 ( .IN1(r806_n281), .IN2(r806_n282), .QN(r806_n46) );
  NAND2X0 r806_U301 ( .IN1(P1_N5152), .IN2(r806_n46), .QN(r806_n278) );
  OR2X1 r806_U300 ( .IN2(P1_N5152), .IN1(r806_n46), .Q(r806_n280) );
  INVX0 r806_U299 ( .ZN(r806_n49), .INP(P1_N3480) );
  NAND2X0 r806_U298 ( .IN1(r806_n280), .IN2(r806_n49), .QN(r806_n279) );
  NAND2X0 r806_U297 ( .IN1(r806_n278), .IN2(r806_n279), .QN(r806_n39) );
  NAND2X0 r806_U296 ( .IN1(P1_N5153), .IN2(r806_n39), .QN(r806_n275) );
  OR2X1 r806_U295 ( .IN2(P1_N5153), .IN1(r806_n39), .Q(r806_n277) );
  INVX0 r806_U294 ( .ZN(r806_n42), .INP(P1_N3481) );
  NAND2X0 r806_U293 ( .IN1(r806_n277), .IN2(r806_n42), .QN(r806_n276) );
  NAND2X0 r806_U292 ( .IN1(r806_n275), .IN2(r806_n276), .QN(r806_n32) );
  NAND2X0 r806_U291 ( .IN1(P1_N5154), .IN2(r806_n32), .QN(r806_n272) );
  OR2X1 r806_U290 ( .IN2(P1_N5154), .IN1(r806_n32), .Q(r806_n274) );
  INVX0 r806_U289 ( .ZN(r806_n35), .INP(P1_N3482) );
  NAND2X0 r806_U288 ( .IN1(r806_n274), .IN2(r806_n35), .QN(r806_n273) );
  NAND2X0 r806_U287 ( .IN1(r806_n272), .IN2(r806_n273), .QN(r806_n25) );
  NAND2X0 r806_U286 ( .IN1(P1_N5155), .IN2(r806_n25), .QN(r806_n269) );
  OR2X1 r806_U285 ( .IN2(P1_N5155), .IN1(r806_n25), .Q(r806_n271) );
  INVX0 r806_U284 ( .ZN(r806_n28), .INP(P1_N3483) );
  NAND2X0 r806_U283 ( .IN1(r806_n271), .IN2(r806_n28), .QN(r806_n270) );
  NAND2X0 r806_U282 ( .IN1(r806_n269), .IN2(r806_n270), .QN(r806_n18) );
  NAND2X0 r806_U281 ( .IN1(n7075), .IN2(r806_n18), .QN(r806_n266) );
  OR2X1 r806_U280 ( .IN2(n7075), .IN1(r806_n18), .Q(r806_n268) );
  INVX0 r806_U279 ( .ZN(r806_n21), .INP(P1_N3484) );
  NAND2X0 r806_U278 ( .IN1(r806_n268), .IN2(r806_n21), .QN(r806_n267) );
  NAND2X0 r806_U277 ( .IN1(r806_n266), .IN2(r806_n267), .QN(r806_n11) );
  NAND2X0 r806_U276 ( .IN1(n7072), .IN2(r806_n11), .QN(r806_n263) );
  OR2X1 r806_U275 ( .IN2(n7072), .IN1(r806_n11), .Q(r806_n265) );
  INVX0 r806_U274 ( .ZN(r806_n14), .INP(P1_N3485) );
  NAND2X0 r806_U273 ( .IN1(r806_n265), .IN2(r806_n14), .QN(r806_n264) );
  NAND2X0 r806_U272 ( .IN1(r806_n263), .IN2(r806_n264), .QN(r806_n4) );
  NAND2X0 r806_U271 ( .IN1(P1_N5158), .IN2(r806_n4), .QN(r806_n260) );
  OR2X1 r806_U270 ( .IN2(P1_N5158), .IN1(r806_n4), .Q(r806_n262) );
  INVX0 r806_U269 ( .ZN(r806_n7), .INP(P1_N3486) );
  NAND2X0 r806_U268 ( .IN1(r806_n262), .IN2(r806_n7), .QN(r806_n261) );
  NAND2X0 r806_U267 ( .IN1(r806_n260), .IN2(r806_n261), .QN(r806_n254) );
  NAND2X0 r806_U266 ( .IN1(r806_n259), .IN2(r806_n254), .QN(r806_n257) );
  OR2X1 r806_U265 ( .IN2(r806_n254), .IN1(r806_n259), .Q(r806_n258) );
  NAND2X0 r806_U264 ( .IN1(r806_n257), .IN2(r806_n258), .QN(P1_N3639) );
  INVX0 r806_U263 ( .ZN(r806_n243), .INP(P1_N3488) );
  NAND2X0 r806_U262 ( .IN1(P1_N5160), .IN2(r806_n243), .QN(r806_n255) );
  OR2X1 r806_U261 ( .IN2(P1_N5160), .IN1(r806_n243), .Q(r806_n256) );
  NAND2X0 r806_U260 ( .IN1(r806_n255), .IN2(r806_n256), .QN(r806_n249) );
  NAND2X0 r806_U259 ( .IN1(P1_N5159), .IN2(r806_n254), .QN(r806_n250) );
  OR2X1 r806_U258 ( .IN2(P1_N5159), .IN1(r806_n254), .Q(r806_n252) );
  NAND2X0 r806_U257 ( .IN1(r806_n252), .IN2(r806_n253), .QN(r806_n251) );
  NAND2X0 r806_U256 ( .IN1(r806_n250), .IN2(r806_n251), .QN(r806_n244) );
  NAND2X0 r806_U255 ( .IN1(r806_n249), .IN2(r806_n244), .QN(r806_n247) );
  OR2X1 r806_U254 ( .IN2(r806_n244), .IN1(r806_n249), .Q(r806_n248) );
  NAND2X0 r806_U253 ( .IN1(r806_n247), .IN2(r806_n248), .QN(P1_N3640) );
  INVX0 r806_U252 ( .ZN(r806_n233), .INP(P1_N3489) );
  NAND2X0 r806_U251 ( .IN1(P1_N5161), .IN2(r806_n233), .QN(r806_n245) );
  OR2X1 r806_U250 ( .IN2(P1_N5161), .IN1(r806_n233), .Q(r806_n246) );
  NAND2X0 r806_U249 ( .IN1(r806_n245), .IN2(r806_n246), .QN(r806_n239) );
  NAND2X0 r806_U248 ( .IN1(P1_N5160), .IN2(r806_n244), .QN(r806_n240) );
  OR2X1 r806_U247 ( .IN2(P1_N5160), .IN1(r806_n244), .Q(r806_n242) );
  NAND2X0 r806_U246 ( .IN1(r806_n242), .IN2(r806_n243), .QN(r806_n241) );
  NAND2X0 r806_U245 ( .IN1(r806_n240), .IN2(r806_n241), .QN(r806_n234) );
  NAND2X0 r806_U244 ( .IN1(r806_n239), .IN2(r806_n234), .QN(r806_n237) );
  OR2X1 r806_U243 ( .IN2(r806_n234), .IN1(r806_n239), .Q(r806_n238) );
  NAND2X0 r806_U242 ( .IN1(r806_n237), .IN2(r806_n238), .QN(P1_N3641) );
  INVX0 r806_U241 ( .ZN(r806_n223), .INP(P1_N3490) );
  NAND2X0 r806_U240 ( .IN1(n7055), .IN2(r806_n223), .QN(r806_n235) );
  OR2X1 r806_U239 ( .IN2(n7055), .IN1(r806_n223), .Q(r806_n236) );
  NAND2X0 r806_U238 ( .IN1(r806_n235), .IN2(r806_n236), .QN(r806_n229) );
  NAND2X0 r806_U237 ( .IN1(P1_N5161), .IN2(r806_n234), .QN(r806_n230) );
  OR2X1 r806_U236 ( .IN2(P1_N5161), .IN1(r806_n234), .Q(r806_n232) );
  NAND2X0 r806_U235 ( .IN1(r806_n232), .IN2(r806_n233), .QN(r806_n231) );
  NAND2X0 r806_U234 ( .IN1(r806_n230), .IN2(r806_n231), .QN(r806_n224) );
  NAND2X0 r806_U233 ( .IN1(r806_n229), .IN2(r806_n224), .QN(r806_n227) );
  OR2X1 r806_U232 ( .IN2(r806_n224), .IN1(r806_n229), .Q(r806_n228) );
  NAND2X0 r806_U231 ( .IN1(r806_n227), .IN2(r806_n228), .QN(P1_N3642) );
  INVX0 r806_U230 ( .ZN(r806_n213), .INP(P1_N3491) );
  NAND2X0 r806_U229 ( .IN1(n7116), .IN2(r806_n213), .QN(r806_n225) );
  OR2X1 r806_U228 ( .IN2(n7116), .IN1(r806_n213), .Q(r806_n226) );
  NAND2X0 r806_U227 ( .IN1(r806_n225), .IN2(r806_n226), .QN(r806_n219) );
  NAND2X0 r806_U226 ( .IN1(P1_N5162), .IN2(r806_n224), .QN(r806_n220) );
  OR2X1 r806_U225 ( .IN2(n7055), .IN1(r806_n224), .Q(r806_n222) );
  NAND2X0 r806_U224 ( .IN1(r806_n222), .IN2(r806_n223), .QN(r806_n221) );
  INVX0 r806_U321 ( .ZN(r806_n291), .INP(P1_N3477) );
  NOR2X0 r806_U320 ( .QN(r806_n287), .IN1(r806_n291), .IN2(n7034) );
  INVX0 r806_U319 ( .ZN(r806_n162), .INP(r806_n287) );
  NAND2X0 r806_U318 ( .IN1(n7034), .IN2(r806_n291), .QN(r806_n290) );
  NAND2X0 r806_U317 ( .IN1(r806_n162), .IN2(r806_n290), .QN(P1_N3629) );
  NAND2X0 r808_U78 ( .IN1(P1_N5176), .IN2(r808_n77), .QN(r808_n74) );
  OR2X1 r808_U77 ( .IN2(P1_N5176), .IN1(r808_n77), .Q(r808_n76) );
  NAND2X0 r808_U76 ( .IN1(P1_N3877), .IN2(r808_n76), .QN(r808_n75) );
  NAND2X0 r808_U75 ( .IN1(r808_n74), .IN2(r808_n75), .QN(r808_n64) );
  OR2X1 r808_U73 ( .IN2(P1_N3878), .IN1(n7117), .Q(r808_n71) );
  NAND2X0 r808_U72 ( .IN1(P1_N3878), .IN2(n7117), .QN(r808_n72) );
  NAND2X0 r808_U71 ( .IN1(r808_n71), .IN2(r808_n72), .QN(r808_n70) );
  NOR2X0 r808_U70 ( .QN(r808_n68), .IN1(r808_n64), .IN2(r808_n70) );
  AND2X1 r808_U69 ( .IN1(r808_n64), .IN2(r808_n70), .Q(r808_n69) );
  NOR2X0 r808_U68 ( .QN(P1_N4030), .IN1(r808_n68), .IN2(r808_n69) );
  OR2X1 r808_U66 ( .IN2(P1_N3879), .IN1(n7146), .Q(r808_n65) );
  NAND2X0 r808_U65 ( .IN1(P1_N3879), .IN2(n7146), .QN(r808_n66) );
  NAND2X0 r808_U64 ( .IN1(r808_n65), .IN2(r808_n66), .QN(r808_n60) );
  NAND2X0 r808_U63 ( .IN1(P1_N5177), .IN2(r808_n64), .QN(r808_n61) );
  OR2X1 r808_U62 ( .IN2(P1_N5177), .IN1(r808_n64), .Q(r808_n63) );
  NAND2X0 r808_U61 ( .IN1(P1_N3878), .IN2(r808_n63), .QN(r808_n62) );
  NAND2X0 r808_U60 ( .IN1(r808_n61), .IN2(r808_n62), .QN(r808_n59) );
  NOR2X0 r808_U59 ( .QN(r808_n57), .IN1(r808_n60), .IN2(r808_n59) );
  AND2X1 r808_U58 ( .IN1(r808_n59), .IN2(r808_n60), .Q(r808_n58) );
  NOR2X0 r808_U57 ( .QN(P1_N4031), .IN1(r808_n57), .IN2(r808_n58) );
  OR2X1 r808_U55 ( .IN2(P1_N3852), .IN1(n7045), .Q(r808_n54) );
  NAND2X0 r808_U54 ( .IN1(P1_N3852), .IN2(n7045), .QN(r808_n55) );
  NAND2X0 r808_U53 ( .IN1(r808_n54), .IN2(r808_n55), .QN(r808_n53) );
  NOR2X0 r808_U52 ( .QN(r808_n50), .IN1(r808_n52), .IN2(r808_n53) );
  AND2X1 r808_U51 ( .IN1(r808_n52), .IN2(r808_n53), .Q(r808_n51) );
  NOR2X0 r808_U50 ( .QN(P1_N4004), .IN1(r808_n50), .IN2(r808_n51) );
  OR2X1 r808_U48 ( .IN2(P1_N3853), .IN1(n7043), .Q(r808_n47) );
  NAND2X0 r808_U47 ( .IN1(P1_N3853), .IN2(n7043), .QN(r808_n48) );
  NAND2X0 r808_U46 ( .IN1(r808_n47), .IN2(r808_n48), .QN(r808_n46) );
  NOR2X0 r808_U45 ( .QN(r808_n43), .IN1(r808_n45), .IN2(r808_n46) );
  AND2X1 r808_U44 ( .IN1(r808_n45), .IN2(r808_n46), .Q(r808_n44) );
  NOR2X0 r808_U43 ( .QN(P1_N4005), .IN1(r808_n43), .IN2(r808_n44) );
  OR2X1 r808_U41 ( .IN2(P1_N3854), .IN1(n7037), .Q(r808_n40) );
  NAND2X0 r808_U40 ( .IN1(P1_N3854), .IN2(n7037), .QN(r808_n41) );
  NAND2X0 r808_U39 ( .IN1(r808_n40), .IN2(r808_n41), .QN(r808_n39) );
  NOR2X0 r808_U38 ( .QN(r808_n36), .IN1(r808_n38), .IN2(r808_n39) );
  AND2X1 r808_U37 ( .IN1(r808_n38), .IN2(r808_n39), .Q(r808_n37) );
  NOR2X0 r808_U36 ( .QN(P1_N4006), .IN1(r808_n36), .IN2(r808_n37) );
  OR2X1 r808_U34 ( .IN2(P1_N3855), .IN1(n7082), .Q(r808_n33) );
  NAND2X0 r808_U33 ( .IN1(P1_N3855), .IN2(n7082), .QN(r808_n34) );
  NAND2X0 r808_U32 ( .IN1(r808_n33), .IN2(r808_n34), .QN(r808_n32) );
  NOR2X0 r808_U31 ( .QN(r808_n29), .IN1(r808_n31), .IN2(r808_n32) );
  AND2X1 r808_U30 ( .IN1(r808_n31), .IN2(r808_n32), .Q(r808_n30) );
  NOR2X0 r808_U29 ( .QN(P1_N4007), .IN1(r808_n29), .IN2(r808_n30) );
  OR2X1 r808_U27 ( .IN2(P1_N3856), .IN1(n7079), .Q(r808_n26) );
  NAND2X0 r808_U26 ( .IN1(P1_N3856), .IN2(n7079), .QN(r808_n27) );
  NAND2X0 r808_U25 ( .IN1(r808_n26), .IN2(r808_n27), .QN(r808_n25) );
  NOR2X0 r808_U24 ( .QN(r808_n22), .IN1(r808_n24), .IN2(r808_n25) );
  AND2X1 r808_U23 ( .IN1(r808_n24), .IN2(r808_n25), .Q(r808_n23) );
  NOR2X0 r808_U22 ( .QN(P1_N4008), .IN1(r808_n22), .IN2(r808_n23) );
  OR2X1 r808_U20 ( .IN2(P1_N3857), .IN1(n7076), .Q(r808_n19) );
  NAND2X0 r808_U19 ( .IN1(P1_N3857), .IN2(n7076), .QN(r808_n20) );
  NAND2X0 r808_U18 ( .IN1(r808_n19), .IN2(r808_n20), .QN(r808_n18) );
  NOR2X0 r808_U17 ( .QN(r808_n15), .IN1(r808_n17), .IN2(r808_n18) );
  AND2X1 r808_U16 ( .IN1(r808_n17), .IN2(r808_n18), .Q(r808_n16) );
  NOR2X0 r808_U15 ( .QN(P1_N4009), .IN1(r808_n15), .IN2(r808_n16) );
  OR2X1 r808_U13 ( .IN2(P1_N3858), .IN1(n7073), .Q(r808_n12) );
  NAND2X0 r808_U12 ( .IN1(P1_N3858), .IN2(n7073), .QN(r808_n13) );
  NAND2X0 r808_U11 ( .IN1(r808_n12), .IN2(r808_n13), .QN(r808_n11) );
  NOR2X0 r808_U10 ( .QN(r808_n8), .IN1(r808_n10), .IN2(r808_n11) );
  AND2X1 r808_U9 ( .IN1(r808_n10), .IN2(r808_n11), .Q(r808_n9) );
  NOR2X0 r808_U8 ( .QN(P1_N4010), .IN1(r808_n8), .IN2(r808_n9) );
  OR2X1 r808_U6 ( .IN2(P1_N3859), .IN1(n7071), .Q(r808_n5) );
  NAND2X0 r808_U5 ( .IN1(P1_N3859), .IN2(n7071), .QN(r808_n6) );
  NAND2X0 r808_U4 ( .IN1(r808_n5), .IN2(r808_n6), .QN(r808_n4) );
  NOR2X0 r808_U3 ( .QN(r808_n1), .IN1(r808_n3), .IN2(r808_n4) );
  AND2X1 r808_U2 ( .IN1(r808_n3), .IN2(r808_n4), .Q(r808_n2) );
  NOR2X0 r808_U1 ( .QN(P1_N4011), .IN1(r808_n1), .IN2(r808_n2) );
  NAND2X0 r808_U171 ( .IN1(P1_N3851), .IN2(n7051), .QN(r808_n163) );
  NAND2X0 r808_U170 ( .IN1(r808_n162), .IN2(r808_n163), .QN(r808_n160) );
  NAND2X0 r808_U169 ( .IN1(r808_n160), .IN2(r808_n161), .QN(r808_n158) );
  OR2X1 r808_U168 ( .IN2(r808_n161), .IN1(r808_n160), .Q(r808_n159) );
  NAND2X0 r808_U167 ( .IN1(r808_n158), .IN2(r808_n159), .QN(P1_N4003) );
  NAND2X0 r808_U166 ( .IN1(n7099), .IN2(r808_n157), .QN(r808_n154) );
  OR2X1 r808_U165 ( .IN2(n7099), .IN1(r808_n157), .Q(r808_n156) );
  NAND2X0 r808_U164 ( .IN1(P1_N3869), .IN2(r808_n156), .QN(r808_n155) );
  NAND2X0 r808_U163 ( .IN1(r808_n154), .IN2(r808_n155), .QN(r808_n147) );
  OR2X1 r808_U161 ( .IN2(P1_N3870), .IN1(n7095), .Q(r808_n151) );
  NAND2X0 r808_U160 ( .IN1(P1_N3870), .IN2(n7095), .QN(r808_n152) );
  NAND2X0 r808_U159 ( .IN1(r808_n151), .IN2(r808_n152), .QN(r808_n150) );
  NOR2X0 r808_U158 ( .QN(r808_n148), .IN1(r808_n147), .IN2(r808_n150) );
  AND2X1 r808_U157 ( .IN1(r808_n147), .IN2(r808_n150), .Q(r808_n149) );
  NOR2X0 r808_U156 ( .QN(P1_N4022), .IN1(r808_n148), .IN2(r808_n149) );
  NAND2X0 r808_U155 ( .IN1(P1_N5169), .IN2(r808_n147), .QN(r808_n144) );
  OR2X1 r808_U154 ( .IN2(P1_N5169), .IN1(r808_n147), .Q(r808_n146) );
  NAND2X0 r808_U153 ( .IN1(P1_N3870), .IN2(r808_n146), .QN(r808_n145) );
  NAND2X0 r808_U152 ( .IN1(r808_n144), .IN2(r808_n145), .QN(r808_n137) );
  OR2X1 r808_U150 ( .IN2(P1_N3871), .IN1(n7092), .Q(r808_n141) );
  NAND2X0 r808_U149 ( .IN1(P1_N3871), .IN2(n7092), .QN(r808_n142) );
  NAND2X0 r808_U148 ( .IN1(r808_n141), .IN2(r808_n142), .QN(r808_n140) );
  NOR2X0 r808_U147 ( .QN(r808_n138), .IN1(r808_n137), .IN2(r808_n140) );
  AND2X1 r808_U146 ( .IN1(r808_n137), .IN2(r808_n140), .Q(r808_n139) );
  NOR2X0 r808_U145 ( .QN(P1_N4023), .IN1(r808_n138), .IN2(r808_n139) );
  NAND2X0 r808_U144 ( .IN1(P1_N5170), .IN2(r808_n137), .QN(r808_n134) );
  OR2X1 r808_U143 ( .IN2(P1_N5170), .IN1(r808_n137), .Q(r808_n136) );
  NAND2X0 r808_U142 ( .IN1(P1_N3871), .IN2(r808_n136), .QN(r808_n135) );
  NAND2X0 r808_U141 ( .IN1(r808_n134), .IN2(r808_n135), .QN(r808_n127) );
  OR2X1 r808_U139 ( .IN2(P1_N3872), .IN1(n7090), .Q(r808_n131) );
  NAND2X0 r808_U138 ( .IN1(P1_N3872), .IN2(n7090), .QN(r808_n132) );
  NAND2X0 r808_U137 ( .IN1(r808_n131), .IN2(r808_n132), .QN(r808_n130) );
  NOR2X0 r808_U136 ( .QN(r808_n128), .IN1(r808_n127), .IN2(r808_n130) );
  AND2X1 r808_U135 ( .IN1(r808_n127), .IN2(r808_n130), .Q(r808_n129) );
  NOR2X0 r808_U134 ( .QN(P1_N4024), .IN1(r808_n128), .IN2(r808_n129) );
  NAND2X0 r808_U133 ( .IN1(P1_N5171), .IN2(r808_n127), .QN(r808_n124) );
  OR2X1 r808_U132 ( .IN2(P1_N5171), .IN1(r808_n127), .Q(r808_n126) );
  NAND2X0 r808_U131 ( .IN1(P1_N3872), .IN2(r808_n126), .QN(r808_n125) );
  NAND2X0 r808_U130 ( .IN1(r808_n124), .IN2(r808_n125), .QN(r808_n117) );
  OR2X1 r808_U128 ( .IN2(P1_N3873), .IN1(n7144), .Q(r808_n121) );
  NAND2X0 r808_U127 ( .IN1(P1_N3873), .IN2(n7144), .QN(r808_n122) );
  NAND2X0 r808_U126 ( .IN1(r808_n121), .IN2(r808_n122), .QN(r808_n120) );
  NOR2X0 r808_U125 ( .QN(r808_n118), .IN1(r808_n117), .IN2(r808_n120) );
  AND2X1 r808_U124 ( .IN1(r808_n117), .IN2(r808_n120), .Q(r808_n119) );
  NOR2X0 r808_U123 ( .QN(P1_N4025), .IN1(r808_n118), .IN2(r808_n119) );
  NAND2X0 r808_U122 ( .IN1(n7141), .IN2(r808_n117), .QN(r808_n114) );
  OR2X1 r808_U121 ( .IN2(n7141), .IN1(r808_n117), .Q(r808_n116) );
  NAND2X0 r808_U120 ( .IN1(P1_N3873), .IN2(r808_n116), .QN(r808_n115) );
  NAND2X0 r808_U119 ( .IN1(r808_n114), .IN2(r808_n115), .QN(r808_n107) );
  OR2X1 r808_U117 ( .IN2(P1_N3874), .IN1(n7136), .Q(r808_n111) );
  NAND2X0 r808_U116 ( .IN1(P1_N3874), .IN2(n7136), .QN(r808_n112) );
  NAND2X0 r808_U115 ( .IN1(r808_n111), .IN2(r808_n112), .QN(r808_n110) );
  NOR2X0 r808_U114 ( .QN(r808_n108), .IN1(r808_n107), .IN2(r808_n110) );
  AND2X1 r808_U113 ( .IN1(r808_n107), .IN2(r808_n110), .Q(r808_n109) );
  NOR2X0 r808_U112 ( .QN(P1_N4026), .IN1(r808_n108), .IN2(r808_n109) );
  NAND2X0 r808_U111 ( .IN1(n7138), .IN2(r808_n107), .QN(r808_n104) );
  OR2X1 r808_U110 ( .IN2(n7138), .IN1(r808_n107), .Q(r808_n106) );
  NAND2X0 r808_U109 ( .IN1(P1_N3874), .IN2(r808_n106), .QN(r808_n105) );
  NAND2X0 r808_U108 ( .IN1(r808_n104), .IN2(r808_n105), .QN(r808_n97) );
  OR2X1 r808_U106 ( .IN2(P1_N3875), .IN1(n7130), .Q(r808_n101) );
  NAND2X0 r808_U105 ( .IN1(P1_N3875), .IN2(n7130), .QN(r808_n102) );
  NAND2X0 r808_U104 ( .IN1(r808_n101), .IN2(r808_n102), .QN(r808_n100) );
  NOR2X0 r808_U103 ( .QN(r808_n98), .IN1(r808_n97), .IN2(r808_n100) );
  AND2X1 r808_U102 ( .IN1(r808_n97), .IN2(r808_n100), .Q(r808_n99) );
  NOR2X0 r808_U101 ( .QN(P1_N4027), .IN1(r808_n98), .IN2(r808_n99) );
  NAND2X0 r808_U100 ( .IN1(n7129), .IN2(r808_n97), .QN(r808_n94) );
  OR2X1 r808_U99 ( .IN2(n7129), .IN1(r808_n97), .Q(r808_n96) );
  NAND2X0 r808_U98 ( .IN1(P1_N3875), .IN2(r808_n96), .QN(r808_n95) );
  NAND2X0 r808_U97 ( .IN1(r808_n94), .IN2(r808_n95), .QN(r808_n87) );
  OR2X1 r808_U95 ( .IN2(P1_N3876), .IN1(n7125), .Q(r808_n91) );
  NAND2X0 r808_U94 ( .IN1(P1_N3876), .IN2(n7125), .QN(r808_n92) );
  NAND2X0 r808_U93 ( .IN1(r808_n91), .IN2(r808_n92), .QN(r808_n90) );
  NOR2X0 r808_U92 ( .QN(r808_n88), .IN1(r808_n87), .IN2(r808_n90) );
  AND2X1 r808_U91 ( .IN1(r808_n87), .IN2(r808_n90), .Q(r808_n89) );
  NOR2X0 r808_U90 ( .QN(P1_N4028), .IN1(r808_n88), .IN2(r808_n89) );
  NAND2X0 r808_U89 ( .IN1(P1_N5175), .IN2(r808_n87), .QN(r808_n84) );
  OR2X1 r808_U88 ( .IN2(P1_N5175), .IN1(r808_n87), .Q(r808_n86) );
  NAND2X0 r808_U87 ( .IN1(P1_N3876), .IN2(r808_n86), .QN(r808_n85) );
  NAND2X0 r808_U86 ( .IN1(r808_n84), .IN2(r808_n85), .QN(r808_n77) );
  OR2X1 r808_U84 ( .IN2(P1_N3877), .IN1(n7119), .Q(r808_n81) );
  NAND2X0 r808_U83 ( .IN1(P1_N3877), .IN2(n7119), .QN(r808_n82) );
  NAND2X0 r808_U82 ( .IN1(r808_n81), .IN2(r808_n82), .QN(r808_n80) );
  NOR2X0 r808_U81 ( .QN(r808_n78), .IN1(r808_n77), .IN2(r808_n80) );
  AND2X1 r808_U80 ( .IN1(r808_n77), .IN2(r808_n80), .Q(r808_n79) );
  NOR2X0 r808_U79 ( .QN(P1_N4029), .IN1(r808_n78), .IN2(r808_n79) );
  NAND2X0 r808_U264 ( .IN1(r808_n248), .IN2(r808_n249), .QN(r808_n247) );
  NOR2X0 r808_U263 ( .QN(r808_n245), .IN1(r808_n244), .IN2(r808_n247) );
  AND2X1 r808_U262 ( .IN1(r808_n244), .IN2(r808_n247), .Q(r808_n246) );
  NOR2X0 r808_U261 ( .QN(P1_N4013), .IN1(r808_n245), .IN2(r808_n246) );
  NAND2X0 r808_U260 ( .IN1(P1_N5160), .IN2(r808_n244), .QN(r808_n241) );
  OR2X1 r808_U259 ( .IN2(P1_N5160), .IN1(r808_n244), .Q(r808_n243) );
  NAND2X0 r808_U258 ( .IN1(P1_N3861), .IN2(r808_n243), .QN(r808_n242) );
  NAND2X0 r808_U257 ( .IN1(r808_n241), .IN2(r808_n242), .QN(r808_n234) );
  OR2X1 r808_U255 ( .IN2(P1_N3862), .IN1(n7058), .Q(r808_n238) );
  NAND2X0 r808_U254 ( .IN1(P1_N3862), .IN2(n7058), .QN(r808_n239) );
  NAND2X0 r808_U253 ( .IN1(r808_n238), .IN2(r808_n239), .QN(r808_n237) );
  NOR2X0 r808_U252 ( .QN(r808_n235), .IN1(r808_n234), .IN2(r808_n237) );
  AND2X1 r808_U251 ( .IN1(r808_n234), .IN2(r808_n237), .Q(r808_n236) );
  NOR2X0 r808_U250 ( .QN(P1_N4014), .IN1(r808_n235), .IN2(r808_n236) );
  NAND2X0 r808_U249 ( .IN1(P1_N5161), .IN2(r808_n234), .QN(r808_n231) );
  OR2X1 r808_U248 ( .IN2(P1_N5161), .IN1(r808_n234), .Q(r808_n233) );
  NAND2X0 r808_U247 ( .IN1(P1_N3862), .IN2(r808_n233), .QN(r808_n232) );
  NAND2X0 r808_U246 ( .IN1(r808_n231), .IN2(r808_n232), .QN(r808_n224) );
  OR2X1 r808_U244 ( .IN2(P1_N3863), .IN1(n7056), .Q(r808_n228) );
  NAND2X0 r808_U243 ( .IN1(P1_N3863), .IN2(n7056), .QN(r808_n229) );
  NAND2X0 r808_U242 ( .IN1(r808_n228), .IN2(r808_n229), .QN(r808_n227) );
  NOR2X0 r808_U241 ( .QN(r808_n225), .IN1(r808_n224), .IN2(r808_n227) );
  AND2X1 r808_U240 ( .IN1(r808_n224), .IN2(r808_n227), .Q(r808_n226) );
  NOR2X0 r808_U239 ( .QN(P1_N4015), .IN1(r808_n225), .IN2(r808_n226) );
  NAND2X0 r808_U238 ( .IN1(P1_N5162), .IN2(r808_n224), .QN(r808_n221) );
  OR2X1 r808_U237 ( .IN2(P1_N5162), .IN1(r808_n224), .Q(r808_n223) );
  NAND2X0 r808_U236 ( .IN1(P1_N3863), .IN2(r808_n223), .QN(r808_n222) );
  NAND2X0 r808_U235 ( .IN1(r808_n221), .IN2(r808_n222), .QN(r808_n214) );
  OR2X1 r808_U233 ( .IN2(P1_N3864), .IN1(n7115), .Q(r808_n218) );
  NAND2X0 r808_U232 ( .IN1(P1_N3864), .IN2(n7115), .QN(r808_n219) );
  NAND2X0 r808_U231 ( .IN1(r808_n218), .IN2(r808_n219), .QN(r808_n217) );
  NOR2X0 r808_U230 ( .QN(r808_n215), .IN1(r808_n214), .IN2(r808_n217) );
  AND2X1 r808_U229 ( .IN1(r808_n214), .IN2(r808_n217), .Q(r808_n216) );
  NOR2X0 r808_U228 ( .QN(P1_N4016), .IN1(r808_n215), .IN2(r808_n216) );
  NAND2X0 r808_U227 ( .IN1(P1_N5163), .IN2(r808_n214), .QN(r808_n211) );
  OR2X1 r808_U226 ( .IN2(P1_N5163), .IN1(r808_n214), .Q(r808_n213) );
  NAND2X0 r808_U225 ( .IN1(P1_N3864), .IN2(r808_n213), .QN(r808_n212) );
  NAND2X0 r808_U224 ( .IN1(r808_n211), .IN2(r808_n212), .QN(r808_n204) );
  OR2X1 r808_U222 ( .IN2(P1_N3865), .IN1(n7112), .Q(r808_n208) );
  NAND2X0 r808_U221 ( .IN1(P1_N3865), .IN2(n7112), .QN(r808_n209) );
  NAND2X0 r808_U220 ( .IN1(r808_n208), .IN2(r808_n209), .QN(r808_n207) );
  NOR2X0 r808_U219 ( .QN(r808_n205), .IN1(r808_n204), .IN2(r808_n207) );
  AND2X1 r808_U218 ( .IN1(r808_n204), .IN2(r808_n207), .Q(r808_n206) );
  NOR2X0 r808_U217 ( .QN(P1_N4017), .IN1(r808_n205), .IN2(r808_n206) );
  NAND2X0 r808_U216 ( .IN1(P1_N5164), .IN2(r808_n204), .QN(r808_n201) );
  OR2X1 r808_U215 ( .IN2(P1_N5164), .IN1(r808_n204), .Q(r808_n203) );
  NAND2X0 r808_U214 ( .IN1(P1_N3865), .IN2(r808_n203), .QN(r808_n202) );
  NAND2X0 r808_U213 ( .IN1(r808_n201), .IN2(r808_n202), .QN(r808_n194) );
  OR2X1 r808_U211 ( .IN2(P1_N3866), .IN1(n7109), .Q(r808_n198) );
  NAND2X0 r808_U210 ( .IN1(P1_N3866), .IN2(n7109), .QN(r808_n199) );
  NAND2X0 r808_U209 ( .IN1(r808_n198), .IN2(r808_n199), .QN(r808_n197) );
  NOR2X0 r808_U208 ( .QN(r808_n195), .IN1(r808_n194), .IN2(r808_n197) );
  AND2X1 r808_U207 ( .IN1(r808_n194), .IN2(r808_n197), .Q(r808_n196) );
  NOR2X0 r808_U206 ( .QN(P1_N4018), .IN1(r808_n195), .IN2(r808_n196) );
  NAND2X0 r808_U205 ( .IN1(P1_N5165), .IN2(r808_n194), .QN(r808_n191) );
  OR2X1 r808_U204 ( .IN2(P1_N5165), .IN1(r808_n194), .Q(r808_n193) );
  NAND2X0 r808_U203 ( .IN1(P1_N3866), .IN2(r808_n193), .QN(r808_n192) );
  NAND2X0 r808_U202 ( .IN1(r808_n191), .IN2(r808_n192), .QN(r808_n184) );
  OR2X1 r808_U200 ( .IN2(P1_N3867), .IN1(n7105), .Q(r808_n188) );
  NAND2X0 r808_U199 ( .IN1(P1_N3867), .IN2(n7105), .QN(r808_n189) );
  NAND2X0 r808_U198 ( .IN1(r808_n188), .IN2(r808_n189), .QN(r808_n187) );
  NOR2X0 r808_U197 ( .QN(r808_n185), .IN1(r808_n184), .IN2(r808_n187) );
  AND2X1 r808_U196 ( .IN1(r808_n184), .IN2(r808_n187), .Q(r808_n186) );
  NOR2X0 r808_U195 ( .QN(P1_N4019), .IN1(r808_n185), .IN2(r808_n186) );
  NAND2X0 r808_U194 ( .IN1(n7106), .IN2(r808_n184), .QN(r808_n181) );
  OR2X1 r808_U193 ( .IN2(n7106), .IN1(r808_n184), .Q(r808_n183) );
  NAND2X0 r808_U192 ( .IN1(P1_N3867), .IN2(r808_n183), .QN(r808_n182) );
  NAND2X0 r808_U191 ( .IN1(r808_n181), .IN2(r808_n182), .QN(r808_n174) );
  OR2X1 r808_U189 ( .IN2(P1_N3868), .IN1(n7102), .Q(r808_n178) );
  NAND2X0 r808_U188 ( .IN1(P1_N3868), .IN2(n7102), .QN(r808_n179) );
  NAND2X0 r808_U187 ( .IN1(r808_n178), .IN2(r808_n179), .QN(r808_n177) );
  NOR2X0 r808_U186 ( .QN(r808_n175), .IN1(r808_n174), .IN2(r808_n177) );
  AND2X1 r808_U185 ( .IN1(r808_n174), .IN2(r808_n177), .Q(r808_n176) );
  NOR2X0 r808_U184 ( .QN(P1_N4020), .IN1(r808_n175), .IN2(r808_n176) );
  NAND2X0 r808_U183 ( .IN1(P1_N5167), .IN2(r808_n174), .QN(r808_n171) );
  OR2X1 r808_U182 ( .IN2(P1_N5167), .IN1(r808_n174), .Q(r808_n173) );
  NAND2X0 r808_U181 ( .IN1(P1_N3868), .IN2(r808_n173), .QN(r808_n172) );
  NAND2X0 r808_U180 ( .IN1(r808_n171), .IN2(r808_n172), .QN(r808_n157) );
  OR2X1 r808_U178 ( .IN2(P1_N3869), .IN1(n7098), .Q(r808_n168) );
  NAND2X0 r808_U177 ( .IN1(P1_N3869), .IN2(n7098), .QN(r808_n169) );
  NAND2X0 r808_U176 ( .IN1(r808_n168), .IN2(r808_n169), .QN(r808_n167) );
  NOR2X0 r808_U175 ( .QN(r808_n165), .IN1(r808_n157), .IN2(r808_n167) );
  AND2X1 r808_U174 ( .IN1(r808_n157), .IN2(r808_n167), .Q(r808_n166) );
  NOR2X0 r808_U173 ( .QN(P1_N4021), .IN1(r808_n165), .IN2(r808_n166) );
  OR2X1 r808_U172 ( .IN2(P1_N3851), .IN1(n7051), .Q(r808_n162) );
  OR2X1 r808_U319 ( .IN2(P1_N3850), .IN1(n4803), .Q(r808_n288) );
  NAND2X0 r808_U318 ( .IN1(P1_N3850), .IN2(n4803), .QN(r808_n289) );
  NAND2X0 r808_U317 ( .IN1(r808_n288), .IN2(r808_n289), .QN(P1_N4002) );
  NAND2X0 r808_U315 ( .IN1(P1_N3850), .IN2(n7034), .QN(r808_n161) );
  OR2X1 r808_U314 ( .IN2(r808_n161), .IN1(n7051), .Q(r808_n285) );
  NAND2X0 r808_U313 ( .IN1(n7051), .IN2(r808_n161), .QN(r808_n287) );
  NAND2X0 r808_U312 ( .IN1(P1_N3851), .IN2(r808_n287), .QN(r808_n286) );
  NAND2X0 r808_U311 ( .IN1(r808_n285), .IN2(r808_n286), .QN(r808_n52) );
  NAND2X0 r808_U310 ( .IN1(P1_N5151), .IN2(r808_n52), .QN(r808_n282) );
  OR2X1 r808_U309 ( .IN2(P1_N5151), .IN1(r808_n52), .Q(r808_n284) );
  NAND2X0 r808_U308 ( .IN1(P1_N3852), .IN2(r808_n284), .QN(r808_n283) );
  NAND2X0 r808_U307 ( .IN1(r808_n282), .IN2(r808_n283), .QN(r808_n45) );
  NAND2X0 r808_U306 ( .IN1(n7041), .IN2(r808_n45), .QN(r808_n279) );
  OR2X1 r808_U305 ( .IN2(n7041), .IN1(r808_n45), .Q(r808_n281) );
  NAND2X0 r808_U304 ( .IN1(P1_N3853), .IN2(r808_n281), .QN(r808_n280) );
  NAND2X0 r808_U303 ( .IN1(r808_n279), .IN2(r808_n280), .QN(r808_n38) );
  NAND2X0 r808_U302 ( .IN1(P1_N5153), .IN2(r808_n38), .QN(r808_n276) );
  OR2X1 r808_U301 ( .IN2(P1_N5153), .IN1(r808_n38), .Q(r808_n278) );
  NAND2X0 r808_U300 ( .IN1(P1_N3854), .IN2(r808_n278), .QN(r808_n277) );
  NAND2X0 r808_U299 ( .IN1(r808_n276), .IN2(r808_n277), .QN(r808_n31) );
  NAND2X0 r808_U298 ( .IN1(P1_N5154), .IN2(r808_n31), .QN(r808_n273) );
  OR2X1 r808_U297 ( .IN2(P1_N5154), .IN1(r808_n31), .Q(r808_n275) );
  NAND2X0 r808_U296 ( .IN1(P1_N3855), .IN2(r808_n275), .QN(r808_n274) );
  NAND2X0 r808_U295 ( .IN1(r808_n273), .IN2(r808_n274), .QN(r808_n24) );
  NAND2X0 r808_U294 ( .IN1(P1_N5155), .IN2(r808_n24), .QN(r808_n270) );
  OR2X1 r808_U293 ( .IN2(P1_N5155), .IN1(r808_n24), .Q(r808_n272) );
  NAND2X0 r808_U292 ( .IN1(P1_N3856), .IN2(r808_n272), .QN(r808_n271) );
  NAND2X0 r808_U291 ( .IN1(r808_n270), .IN2(r808_n271), .QN(r808_n17) );
  NAND2X0 r808_U290 ( .IN1(n7075), .IN2(r808_n17), .QN(r808_n267) );
  OR2X1 r808_U289 ( .IN2(n7075), .IN1(r808_n17), .Q(r808_n269) );
  NAND2X0 r808_U288 ( .IN1(P1_N3857), .IN2(r808_n269), .QN(r808_n268) );
  NAND2X0 r808_U287 ( .IN1(r808_n267), .IN2(r808_n268), .QN(r808_n10) );
  NAND2X0 r808_U286 ( .IN1(n7072), .IN2(r808_n10), .QN(r808_n264) );
  OR2X1 r808_U285 ( .IN2(n7072), .IN1(r808_n10), .Q(r808_n266) );
  NAND2X0 r808_U284 ( .IN1(P1_N3858), .IN2(r808_n266), .QN(r808_n265) );
  NAND2X0 r808_U283 ( .IN1(r808_n264), .IN2(r808_n265), .QN(r808_n3) );
  NAND2X0 r808_U282 ( .IN1(P1_N5158), .IN2(r808_n3), .QN(r808_n261) );
  OR2X1 r808_U281 ( .IN2(P1_N5158), .IN1(r808_n3), .Q(r808_n263) );
  NAND2X0 r808_U280 ( .IN1(P1_N3859), .IN2(r808_n263), .QN(r808_n262) );
  NAND2X0 r808_U279 ( .IN1(r808_n261), .IN2(r808_n262), .QN(r808_n254) );
  OR2X1 r808_U277 ( .IN2(P1_N3860), .IN1(n7067), .Q(r808_n258) );
  NAND2X0 r808_U276 ( .IN1(P1_N3860), .IN2(n7067), .QN(r808_n259) );
  NAND2X0 r808_U275 ( .IN1(r808_n258), .IN2(r808_n259), .QN(r808_n257) );
  NOR2X0 r808_U274 ( .QN(r808_n255), .IN1(r808_n254), .IN2(r808_n257) );
  AND2X1 r808_U273 ( .IN1(r808_n254), .IN2(r808_n257), .Q(r808_n256) );
  NOR2X0 r808_U272 ( .QN(P1_N4012), .IN1(r808_n255), .IN2(r808_n256) );
  NAND2X0 r808_U271 ( .IN1(P1_N5159), .IN2(r808_n254), .QN(r808_n251) );
  OR2X1 r808_U270 ( .IN2(P1_N5159), .IN1(r808_n254), .Q(r808_n253) );
  NAND2X0 r808_U269 ( .IN1(P1_N3860), .IN2(r808_n253), .QN(r808_n252) );
  NAND2X0 r808_U268 ( .IN1(r808_n251), .IN2(r808_n252), .QN(r808_n244) );
  OR2X1 r808_U266 ( .IN2(P1_N3861), .IN1(n7063), .Q(r808_n248) );
  NAND2X0 r808_U265 ( .IN1(P1_N3861), .IN2(n7063), .QN(r808_n249) );
  NAND2X0 r810_U27 ( .IN1(r810_n31), .IN2(r810_n32), .QN(r810_n29) );
  OR2X1 r810_U26 ( .IN2(r810_n32), .IN1(r810_n31), .Q(r810_n30) );
  NAND2X0 r810_U25 ( .IN1(r810_n29), .IN2(r810_n30), .QN(P1_N4380) );
  NAND2X0 r810_U24 ( .IN1(n7080), .IN2(r810_n28), .QN(r810_n26) );
  OR2X1 r810_U23 ( .IN2(n7080), .IN1(r810_n28), .Q(r810_n27) );
  NAND2X0 r810_U22 ( .IN1(r810_n26), .IN2(r810_n27), .QN(r810_n24) );
  NAND2X0 r810_U21 ( .IN1(r810_n24), .IN2(r810_n25), .QN(r810_n22) );
  OR2X1 r810_U20 ( .IN2(r810_n25), .IN1(r810_n24), .Q(r810_n23) );
  NAND2X0 r810_U19 ( .IN1(r810_n22), .IN2(r810_n23), .QN(P1_N4381) );
  NAND2X0 r810_U18 ( .IN1(P1_N5156), .IN2(r810_n21), .QN(r810_n19) );
  OR2X1 r810_U17 ( .IN2(P1_N5156), .IN1(r810_n21), .Q(r810_n20) );
  NAND2X0 r810_U16 ( .IN1(r810_n19), .IN2(r810_n20), .QN(r810_n17) );
  NAND2X0 r810_U15 ( .IN1(r810_n17), .IN2(r810_n18), .QN(r810_n15) );
  OR2X1 r810_U14 ( .IN2(r810_n18), .IN1(r810_n17), .Q(r810_n16) );
  NAND2X0 r810_U13 ( .IN1(r810_n15), .IN2(r810_n16), .QN(P1_N4382) );
  NAND2X0 r810_U12 ( .IN1(P1_N5157), .IN2(r810_n14), .QN(r810_n12) );
  OR2X1 r810_U11 ( .IN2(P1_N5157), .IN1(r810_n14), .Q(r810_n13) );
  NAND2X0 r810_U10 ( .IN1(r810_n12), .IN2(r810_n13), .QN(r810_n10) );
  NAND2X0 r810_U9 ( .IN1(r810_n10), .IN2(r810_n11), .QN(r810_n8) );
  OR2X1 r810_U8 ( .IN2(r810_n11), .IN1(r810_n10), .Q(r810_n9) );
  NAND2X0 r810_U7 ( .IN1(r810_n8), .IN2(r810_n9), .QN(P1_N4383) );
  NAND2X0 r810_U6 ( .IN1(n7070), .IN2(r810_n7), .QN(r810_n5) );
  OR2X1 r810_U5 ( .IN2(n7070), .IN1(r810_n7), .Q(r810_n6) );
  NAND2X0 r810_U4 ( .IN1(r810_n5), .IN2(r810_n6), .QN(r810_n3) );
  NAND2X0 r810_U3 ( .IN1(r810_n3), .IN2(r810_n4), .QN(r810_n1) );
  OR2X1 r810_U2 ( .IN2(r810_n4), .IN1(r810_n3), .Q(r810_n2) );
  NAND2X0 r810_U1 ( .IN1(r810_n1), .IN2(r810_n2), .QN(P1_N4384) );
  OR2X1 r810_U120 ( .IN2(n7089), .IN1(r810_n126), .Q(r810_n124) );
  NAND2X0 r810_U119 ( .IN1(r810_n124), .IN2(r810_n125), .QN(r810_n123) );
  NAND2X0 r810_U118 ( .IN1(r810_n122), .IN2(r810_n123), .QN(r810_n116) );
  NAND2X0 r810_U117 ( .IN1(r810_n121), .IN2(r810_n116), .QN(r810_n119) );
  OR2X1 r810_U116 ( .IN2(r810_n116), .IN1(r810_n121), .Q(r810_n120) );
  NAND2X0 r810_U115 ( .IN1(r810_n119), .IN2(r810_n120), .QN(P1_N4398) );
  INVX0 r810_U114 ( .ZN(r810_n105), .INP(P1_N4247) );
  NAND2X0 r810_U113 ( .IN1(n7138), .IN2(r810_n105), .QN(r810_n117) );
  OR2X1 r810_U112 ( .IN2(n7138), .IN1(r810_n105), .Q(r810_n118) );
  NAND2X0 r810_U111 ( .IN1(r810_n117), .IN2(r810_n118), .QN(r810_n111) );
  NAND2X0 r810_U110 ( .IN1(P1_N5172), .IN2(r810_n116), .QN(r810_n112) );
  OR2X1 r810_U109 ( .IN2(P1_N5172), .IN1(r810_n116), .Q(r810_n114) );
  NAND2X0 r810_U108 ( .IN1(r810_n114), .IN2(r810_n115), .QN(r810_n113) );
  NAND2X0 r810_U107 ( .IN1(r810_n112), .IN2(r810_n113), .QN(r810_n106) );
  NAND2X0 r810_U106 ( .IN1(r810_n111), .IN2(r810_n106), .QN(r810_n109) );
  OR2X1 r810_U105 ( .IN2(r810_n106), .IN1(r810_n111), .Q(r810_n110) );
  NAND2X0 r810_U104 ( .IN1(r810_n109), .IN2(r810_n110), .QN(P1_N4399) );
  INVX0 r810_U103 ( .ZN(r810_n95), .INP(P1_N4248) );
  NAND2X0 r810_U102 ( .IN1(P1_N5174), .IN2(r810_n95), .QN(r810_n107) );
  OR2X1 r810_U101 ( .IN2(P1_N5174), .IN1(r810_n95), .Q(r810_n108) );
  NAND2X0 r810_U100 ( .IN1(r810_n107), .IN2(r810_n108), .QN(r810_n101) );
  NAND2X0 r810_U99 ( .IN1(n7138), .IN2(r810_n106), .QN(r810_n102) );
  OR2X1 r810_U98 ( .IN2(n7138), .IN1(r810_n106), .Q(r810_n104) );
  NAND2X0 r810_U97 ( .IN1(r810_n104), .IN2(r810_n105), .QN(r810_n103) );
  NAND2X0 r810_U96 ( .IN1(r810_n102), .IN2(r810_n103), .QN(r810_n96) );
  NAND2X0 r810_U95 ( .IN1(r810_n101), .IN2(r810_n96), .QN(r810_n99) );
  OR2X1 r810_U94 ( .IN2(r810_n96), .IN1(r810_n101), .Q(r810_n100) );
  NAND2X0 r810_U93 ( .IN1(r810_n99), .IN2(r810_n100), .QN(P1_N4400) );
  INVX0 r810_U92 ( .ZN(r810_n85), .INP(P1_N4249) );
  NAND2X0 r810_U91 ( .IN1(n7124), .IN2(r810_n85), .QN(r810_n97) );
  OR2X1 r810_U90 ( .IN2(n7124), .IN1(r810_n85), .Q(r810_n98) );
  NAND2X0 r810_U89 ( .IN1(r810_n97), .IN2(r810_n98), .QN(r810_n91) );
  NAND2X0 r810_U88 ( .IN1(P1_N5174), .IN2(r810_n96), .QN(r810_n92) );
  OR2X1 r810_U87 ( .IN2(P1_N5174), .IN1(r810_n96), .Q(r810_n94) );
  NAND2X0 r810_U86 ( .IN1(r810_n94), .IN2(r810_n95), .QN(r810_n93) );
  NAND2X0 r810_U85 ( .IN1(r810_n92), .IN2(r810_n93), .QN(r810_n86) );
  NAND2X0 r810_U84 ( .IN1(r810_n91), .IN2(r810_n86), .QN(r810_n89) );
  OR2X1 r810_U83 ( .IN2(r810_n86), .IN1(r810_n91), .Q(r810_n90) );
  NAND2X0 r810_U82 ( .IN1(r810_n89), .IN2(r810_n90), .QN(P1_N4401) );
  INVX0 r810_U81 ( .ZN(r810_n75), .INP(P1_N4250) );
  NAND2X0 r810_U80 ( .IN1(n7122), .IN2(r810_n75), .QN(r810_n87) );
  OR2X1 r810_U79 ( .IN2(n7122), .IN1(r810_n75), .Q(r810_n88) );
  NAND2X0 r810_U78 ( .IN1(r810_n87), .IN2(r810_n88), .QN(r810_n81) );
  NAND2X0 r810_U77 ( .IN1(n7124), .IN2(r810_n86), .QN(r810_n82) );
  OR2X1 r810_U76 ( .IN2(n7124), .IN1(r810_n86), .Q(r810_n84) );
  NAND2X0 r810_U75 ( .IN1(r810_n84), .IN2(r810_n85), .QN(r810_n83) );
  NAND2X0 r810_U74 ( .IN1(r810_n82), .IN2(r810_n83), .QN(r810_n76) );
  NAND2X0 r810_U73 ( .IN1(r810_n81), .IN2(r810_n76), .QN(r810_n79) );
  OR2X1 r810_U72 ( .IN2(r810_n76), .IN1(r810_n81), .Q(r810_n80) );
  NAND2X0 r810_U71 ( .IN1(r810_n79), .IN2(r810_n80), .QN(P1_N4402) );
  INVX0 r810_U70 ( .ZN(r810_n64), .INP(P1_N4251) );
  NAND2X0 r810_U69 ( .IN1(P1_N5177), .IN2(r810_n64), .QN(r810_n77) );
  OR2X1 r810_U68 ( .IN2(P1_N5177), .IN1(r810_n64), .Q(r810_n78) );
  NAND2X0 r810_U67 ( .IN1(r810_n77), .IN2(r810_n78), .QN(r810_n71) );
  NAND2X0 r810_U66 ( .IN1(n7122), .IN2(r810_n76), .QN(r810_n72) );
  OR2X1 r810_U65 ( .IN2(n7122), .IN1(r810_n76), .Q(r810_n74) );
  NAND2X0 r810_U64 ( .IN1(r810_n74), .IN2(r810_n75), .QN(r810_n73) );
  NAND2X0 r810_U63 ( .IN1(r810_n72), .IN2(r810_n73), .QN(r810_n65) );
  NAND2X0 r810_U62 ( .IN1(r810_n71), .IN2(r810_n65), .QN(r810_n69) );
  OR2X1 r810_U61 ( .IN2(r810_n65), .IN1(r810_n71), .Q(r810_n70) );
  NAND2X0 r810_U60 ( .IN1(r810_n69), .IN2(r810_n70), .QN(P1_N4403) );
  OR2X1 r810_U58 ( .IN2(P1_N4252), .IN1(n7146), .Q(r810_n66) );
  NAND2X0 r810_U57 ( .IN1(P1_N4252), .IN2(n7146), .QN(r810_n67) );
  NAND2X0 r810_U56 ( .IN1(r810_n66), .IN2(r810_n67), .QN(r810_n60) );
  NAND2X0 r810_U55 ( .IN1(P1_N5177), .IN2(r810_n65), .QN(r810_n61) );
  OR2X1 r810_U54 ( .IN2(P1_N5177), .IN1(r810_n65), .Q(r810_n63) );
  NAND2X0 r810_U53 ( .IN1(r810_n63), .IN2(r810_n64), .QN(r810_n62) );
  NAND2X0 r810_U52 ( .IN1(r810_n61), .IN2(r810_n62), .QN(r810_n59) );
  NAND2X0 r810_U51 ( .IN1(r810_n60), .IN2(r810_n59), .QN(r810_n57) );
  OR2X1 r810_U50 ( .IN2(r810_n60), .IN1(r810_n59), .Q(r810_n58) );
  NAND2X0 r810_U49 ( .IN1(r810_n57), .IN2(r810_n58), .QN(P1_N4404) );
  NAND2X0 r810_U48 ( .IN1(n7046), .IN2(r810_n56), .QN(r810_n54) );
  OR2X1 r810_U47 ( .IN2(n7046), .IN1(r810_n56), .Q(r810_n55) );
  NAND2X0 r810_U46 ( .IN1(r810_n54), .IN2(r810_n55), .QN(r810_n52) );
  NAND2X0 r810_U45 ( .IN1(r810_n52), .IN2(r810_n53), .QN(r810_n50) );
  OR2X1 r810_U44 ( .IN2(r810_n53), .IN1(r810_n52), .Q(r810_n51) );
  NAND2X0 r810_U43 ( .IN1(r810_n50), .IN2(r810_n51), .QN(P1_N4377) );
  NAND2X0 r810_U42 ( .IN1(n7041), .IN2(r810_n49), .QN(r810_n47) );
  OR2X1 r810_U41 ( .IN2(n7041), .IN1(r810_n49), .Q(r810_n48) );
  NAND2X0 r810_U40 ( .IN1(r810_n47), .IN2(r810_n48), .QN(r810_n45) );
  NAND2X0 r810_U39 ( .IN1(r810_n45), .IN2(r810_n46), .QN(r810_n43) );
  OR2X1 r810_U38 ( .IN2(r810_n46), .IN1(r810_n45), .Q(r810_n44) );
  NAND2X0 r810_U37 ( .IN1(r810_n43), .IN2(r810_n44), .QN(P1_N4378) );
  NAND2X0 r810_U36 ( .IN1(n7036), .IN2(r810_n42), .QN(r810_n40) );
  OR2X1 r810_U35 ( .IN2(n7036), .IN1(r810_n42), .Q(r810_n41) );
  NAND2X0 r810_U34 ( .IN1(r810_n40), .IN2(r810_n41), .QN(r810_n38) );
  NAND2X0 r810_U33 ( .IN1(r810_n38), .IN2(r810_n39), .QN(r810_n36) );
  OR2X1 r810_U32 ( .IN2(r810_n39), .IN1(r810_n38), .Q(r810_n37) );
  NAND2X0 r810_U31 ( .IN1(r810_n36), .IN2(r810_n37), .QN(P1_N4379) );
  NAND2X0 r810_U30 ( .IN1(n7081), .IN2(r810_n35), .QN(r810_n33) );
  OR2X1 r810_U29 ( .IN2(n7081), .IN1(r810_n35), .Q(r810_n34) );
  NAND2X0 r810_U28 ( .IN1(r810_n33), .IN2(r810_n34), .QN(r810_n31) );
  NAND2X0 r810_U213 ( .IN1(r810_n212), .IN2(r810_n213), .QN(r810_n211) );
  NAND2X0 r810_U212 ( .IN1(r810_n210), .IN2(r810_n211), .QN(r810_n204) );
  NAND2X0 r810_U211 ( .IN1(r810_n209), .IN2(r810_n204), .QN(r810_n207) );
  OR2X1 r810_U210 ( .IN2(r810_n204), .IN1(r810_n209), .Q(r810_n208) );
  NAND2X0 r810_U209 ( .IN1(r810_n207), .IN2(r810_n208), .QN(P1_N4390) );
  INVX0 r810_U208 ( .ZN(r810_n193), .INP(P1_N4239) );
  NAND2X0 r810_U207 ( .IN1(P1_N5165), .IN2(r810_n193), .QN(r810_n205) );
  OR2X1 r810_U206 ( .IN2(P1_N5165), .IN1(r810_n193), .Q(r810_n206) );
  NAND2X0 r810_U205 ( .IN1(r810_n205), .IN2(r810_n206), .QN(r810_n199) );
  NAND2X0 r810_U204 ( .IN1(P1_N5164), .IN2(r810_n204), .QN(r810_n200) );
  OR2X1 r810_U203 ( .IN2(P1_N5164), .IN1(r810_n204), .Q(r810_n202) );
  NAND2X0 r810_U202 ( .IN1(r810_n202), .IN2(r810_n203), .QN(r810_n201) );
  NAND2X0 r810_U201 ( .IN1(r810_n200), .IN2(r810_n201), .QN(r810_n194) );
  NAND2X0 r810_U200 ( .IN1(r810_n199), .IN2(r810_n194), .QN(r810_n197) );
  OR2X1 r810_U199 ( .IN2(r810_n194), .IN1(r810_n199), .Q(r810_n198) );
  NAND2X0 r810_U198 ( .IN1(r810_n197), .IN2(r810_n198), .QN(P1_N4391) );
  INVX0 r810_U197 ( .ZN(r810_n183), .INP(P1_N4240) );
  NAND2X0 r810_U196 ( .IN1(n7106), .IN2(r810_n183), .QN(r810_n195) );
  OR2X1 r810_U195 ( .IN2(n7106), .IN1(r810_n183), .Q(r810_n196) );
  NAND2X0 r810_U194 ( .IN1(r810_n195), .IN2(r810_n196), .QN(r810_n189) );
  NAND2X0 r810_U193 ( .IN1(n7110), .IN2(r810_n194), .QN(r810_n190) );
  OR2X1 r810_U192 ( .IN2(n7110), .IN1(r810_n194), .Q(r810_n192) );
  NAND2X0 r810_U191 ( .IN1(r810_n192), .IN2(r810_n193), .QN(r810_n191) );
  NAND2X0 r810_U190 ( .IN1(r810_n190), .IN2(r810_n191), .QN(r810_n184) );
  NAND2X0 r810_U189 ( .IN1(r810_n189), .IN2(r810_n184), .QN(r810_n187) );
  OR2X1 r810_U188 ( .IN2(r810_n184), .IN1(r810_n189), .Q(r810_n188) );
  NAND2X0 r810_U187 ( .IN1(r810_n187), .IN2(r810_n188), .QN(P1_N4392) );
  INVX0 r810_U186 ( .ZN(r810_n173), .INP(P1_N4241) );
  NAND2X0 r810_U185 ( .IN1(P1_N5167), .IN2(r810_n173), .QN(r810_n185) );
  OR2X1 r810_U184 ( .IN2(P1_N5167), .IN1(r810_n173), .Q(r810_n186) );
  NAND2X0 r810_U183 ( .IN1(r810_n185), .IN2(r810_n186), .QN(r810_n179) );
  NAND2X0 r810_U182 ( .IN1(n7106), .IN2(r810_n184), .QN(r810_n180) );
  OR2X1 r810_U181 ( .IN2(n7106), .IN1(r810_n184), .Q(r810_n182) );
  NAND2X0 r810_U180 ( .IN1(r810_n182), .IN2(r810_n183), .QN(r810_n181) );
  NAND2X0 r810_U179 ( .IN1(r810_n180), .IN2(r810_n181), .QN(r810_n174) );
  NAND2X0 r810_U178 ( .IN1(r810_n179), .IN2(r810_n174), .QN(r810_n177) );
  OR2X1 r810_U177 ( .IN2(r810_n174), .IN1(r810_n179), .Q(r810_n178) );
  NAND2X0 r810_U176 ( .IN1(r810_n177), .IN2(r810_n178), .QN(P1_N4393) );
  INVX0 r810_U175 ( .ZN(r810_n155), .INP(P1_N4242) );
  NAND2X0 r810_U174 ( .IN1(n7099), .IN2(r810_n155), .QN(r810_n175) );
  OR2X1 r810_U173 ( .IN2(n7099), .IN1(r810_n155), .Q(r810_n176) );
  NAND2X0 r810_U172 ( .IN1(r810_n175), .IN2(r810_n176), .QN(r810_n169) );
  NAND2X0 r810_U171 ( .IN1(P1_N5167), .IN2(r810_n174), .QN(r810_n170) );
  OR2X1 r810_U170 ( .IN2(P1_N5167), .IN1(r810_n174), .Q(r810_n172) );
  NAND2X0 r810_U169 ( .IN1(r810_n172), .IN2(r810_n173), .QN(r810_n171) );
  NAND2X0 r810_U168 ( .IN1(r810_n170), .IN2(r810_n171), .QN(r810_n156) );
  NAND2X0 r810_U167 ( .IN1(r810_n169), .IN2(r810_n156), .QN(r810_n167) );
  OR2X1 r810_U166 ( .IN2(r810_n156), .IN1(r810_n169), .Q(r810_n168) );
  NAND2X0 r810_U165 ( .IN1(r810_n167), .IN2(r810_n168), .QN(P1_N4394) );
  NAND2X0 r810_U164 ( .IN1(P1_N5150), .IN2(r810_n166), .QN(r810_n163) );
  NAND2X0 r810_U163 ( .IN1(P1_N4224), .IN2(n7051), .QN(r810_n164) );
  NAND2X0 r810_U162 ( .IN1(r810_n163), .IN2(r810_n164), .QN(r810_n161) );
  NAND2X0 r810_U161 ( .IN1(r810_n161), .IN2(r810_n162), .QN(r810_n159) );
  OR2X1 r810_U160 ( .IN2(r810_n162), .IN1(r810_n161), .Q(r810_n160) );
  NAND2X0 r810_U159 ( .IN1(r810_n159), .IN2(r810_n160), .QN(P1_N4376) );
  INVX0 r810_U158 ( .ZN(r810_n145), .INP(P1_N4243) );
  NAND2X0 r810_U157 ( .IN1(P1_N5169), .IN2(r810_n145), .QN(r810_n157) );
  OR2X1 r810_U156 ( .IN2(P1_N5169), .IN1(r810_n145), .Q(r810_n158) );
  NAND2X0 r810_U155 ( .IN1(r810_n157), .IN2(r810_n158), .QN(r810_n151) );
  NAND2X0 r810_U154 ( .IN1(n7099), .IN2(r810_n156), .QN(r810_n152) );
  OR2X1 r810_U153 ( .IN2(n7099), .IN1(r810_n156), .Q(r810_n154) );
  NAND2X0 r810_U152 ( .IN1(r810_n154), .IN2(r810_n155), .QN(r810_n153) );
  NAND2X0 r810_U151 ( .IN1(r810_n152), .IN2(r810_n153), .QN(r810_n146) );
  NAND2X0 r810_U150 ( .IN1(r810_n151), .IN2(r810_n146), .QN(r810_n149) );
  OR2X1 r810_U149 ( .IN2(r810_n146), .IN1(r810_n151), .Q(r810_n150) );
  NAND2X0 r810_U148 ( .IN1(r810_n149), .IN2(r810_n150), .QN(P1_N4395) );
  INVX0 r810_U147 ( .ZN(r810_n135), .INP(P1_N4244) );
  NAND2X0 r810_U146 ( .IN1(P1_N5170), .IN2(r810_n135), .QN(r810_n147) );
  OR2X1 r810_U145 ( .IN2(P1_N5170), .IN1(r810_n135), .Q(r810_n148) );
  NAND2X0 r810_U144 ( .IN1(r810_n147), .IN2(r810_n148), .QN(r810_n141) );
  NAND2X0 r810_U143 ( .IN1(P1_N5169), .IN2(r810_n146), .QN(r810_n142) );
  OR2X1 r810_U142 ( .IN2(P1_N5169), .IN1(r810_n146), .Q(r810_n144) );
  NAND2X0 r810_U141 ( .IN1(r810_n144), .IN2(r810_n145), .QN(r810_n143) );
  NAND2X0 r810_U140 ( .IN1(r810_n142), .IN2(r810_n143), .QN(r810_n136) );
  NAND2X0 r810_U139 ( .IN1(r810_n141), .IN2(r810_n136), .QN(r810_n139) );
  OR2X1 r810_U138 ( .IN2(r810_n136), .IN1(r810_n141), .Q(r810_n140) );
  NAND2X0 r810_U137 ( .IN1(r810_n139), .IN2(r810_n140), .QN(P1_N4396) );
  INVX0 r810_U136 ( .ZN(r810_n125), .INP(P1_N4245) );
  NAND2X0 r810_U135 ( .IN1(n7089), .IN2(r810_n125), .QN(r810_n137) );
  OR2X1 r810_U134 ( .IN2(n7089), .IN1(r810_n125), .Q(r810_n138) );
  NAND2X0 r810_U133 ( .IN1(r810_n137), .IN2(r810_n138), .QN(r810_n131) );
  NAND2X0 r810_U132 ( .IN1(P1_N5170), .IN2(r810_n136), .QN(r810_n132) );
  OR2X1 r810_U131 ( .IN2(P1_N5170), .IN1(r810_n136), .Q(r810_n134) );
  NAND2X0 r810_U130 ( .IN1(r810_n134), .IN2(r810_n135), .QN(r810_n133) );
  NAND2X0 r810_U129 ( .IN1(r810_n132), .IN2(r810_n133), .QN(r810_n126) );
  NAND2X0 r810_U128 ( .IN1(r810_n131), .IN2(r810_n126), .QN(r810_n129) );
  OR2X1 r810_U127 ( .IN2(r810_n126), .IN1(r810_n131), .Q(r810_n130) );
  NAND2X0 r810_U126 ( .IN1(r810_n129), .IN2(r810_n130), .QN(P1_N4397) );
  INVX0 r810_U125 ( .ZN(r810_n115), .INP(P1_N4246) );
  NAND2X0 r810_U124 ( .IN1(P1_N5172), .IN2(r810_n115), .QN(r810_n127) );
  OR2X1 r810_U123 ( .IN2(P1_N5172), .IN1(r810_n115), .Q(r810_n128) );
  NAND2X0 r810_U122 ( .IN1(r810_n127), .IN2(r810_n128), .QN(r810_n121) );
  NAND2X0 r810_U121 ( .IN1(n7089), .IN2(r810_n126), .QN(r810_n122) );
  NAND2X0 r810_U306 ( .IN1(n7046), .IN2(r810_n53), .QN(r810_n281) );
  OR2X1 r810_U305 ( .IN2(n7046), .IN1(r810_n53), .Q(r810_n283) );
  INVX0 r810_U304 ( .ZN(r810_n56), .INP(P1_N4225) );
  NAND2X0 r810_U303 ( .IN1(r810_n283), .IN2(r810_n56), .QN(r810_n282) );
  NAND2X0 r810_U302 ( .IN1(r810_n281), .IN2(r810_n282), .QN(r810_n46) );
  NAND2X0 r810_U301 ( .IN1(n7041), .IN2(r810_n46), .QN(r810_n278) );
  OR2X1 r810_U300 ( .IN2(n7041), .IN1(r810_n46), .Q(r810_n280) );
  INVX0 r810_U299 ( .ZN(r810_n49), .INP(P1_N4226) );
  NAND2X0 r810_U298 ( .IN1(r810_n280), .IN2(r810_n49), .QN(r810_n279) );
  NAND2X0 r810_U297 ( .IN1(r810_n278), .IN2(r810_n279), .QN(r810_n39) );
  NAND2X0 r810_U296 ( .IN1(n7036), .IN2(r810_n39), .QN(r810_n275) );
  OR2X1 r810_U295 ( .IN2(n7036), .IN1(r810_n39), .Q(r810_n277) );
  INVX0 r810_U294 ( .ZN(r810_n42), .INP(P1_N4227) );
  NAND2X0 r810_U293 ( .IN1(r810_n277), .IN2(r810_n42), .QN(r810_n276) );
  NAND2X0 r810_U292 ( .IN1(r810_n275), .IN2(r810_n276), .QN(r810_n32) );
  NAND2X0 r810_U291 ( .IN1(n7081), .IN2(r810_n32), .QN(r810_n272) );
  OR2X1 r810_U290 ( .IN2(n7081), .IN1(r810_n32), .Q(r810_n274) );
  INVX0 r810_U289 ( .ZN(r810_n35), .INP(P1_N4228) );
  NAND2X0 r810_U288 ( .IN1(r810_n274), .IN2(r810_n35), .QN(r810_n273) );
  NAND2X0 r810_U287 ( .IN1(r810_n272), .IN2(r810_n273), .QN(r810_n25) );
  NAND2X0 r810_U286 ( .IN1(n7080), .IN2(r810_n25), .QN(r810_n269) );
  OR2X1 r810_U285 ( .IN2(n7080), .IN1(r810_n25), .Q(r810_n271) );
  INVX0 r810_U284 ( .ZN(r810_n28), .INP(P1_N4229) );
  NAND2X0 r810_U283 ( .IN1(r810_n271), .IN2(r810_n28), .QN(r810_n270) );
  NAND2X0 r810_U282 ( .IN1(r810_n269), .IN2(r810_n270), .QN(r810_n18) );
  NAND2X0 r810_U281 ( .IN1(P1_N5156), .IN2(r810_n18), .QN(r810_n266) );
  OR2X1 r810_U280 ( .IN2(P1_N5156), .IN1(r810_n18), .Q(r810_n268) );
  INVX0 r810_U279 ( .ZN(r810_n21), .INP(P1_N4230) );
  NAND2X0 r810_U278 ( .IN1(r810_n268), .IN2(r810_n21), .QN(r810_n267) );
  NAND2X0 r810_U277 ( .IN1(r810_n266), .IN2(r810_n267), .QN(r810_n11) );
  NAND2X0 r810_U276 ( .IN1(P1_N5157), .IN2(r810_n11), .QN(r810_n263) );
  OR2X1 r810_U275 ( .IN2(P1_N5157), .IN1(r810_n11), .Q(r810_n265) );
  INVX0 r810_U274 ( .ZN(r810_n14), .INP(P1_N4231) );
  NAND2X0 r810_U273 ( .IN1(r810_n265), .IN2(r810_n14), .QN(r810_n264) );
  NAND2X0 r810_U272 ( .IN1(r810_n263), .IN2(r810_n264), .QN(r810_n4) );
  NAND2X0 r810_U271 ( .IN1(n7070), .IN2(r810_n4), .QN(r810_n260) );
  OR2X1 r810_U270 ( .IN2(n7070), .IN1(r810_n4), .Q(r810_n262) );
  INVX0 r810_U269 ( .ZN(r810_n7), .INP(P1_N4232) );
  NAND2X0 r810_U268 ( .IN1(r810_n262), .IN2(r810_n7), .QN(r810_n261) );
  NAND2X0 r810_U267 ( .IN1(r810_n260), .IN2(r810_n261), .QN(r810_n254) );
  NAND2X0 r810_U266 ( .IN1(r810_n259), .IN2(r810_n254), .QN(r810_n257) );
  OR2X1 r810_U265 ( .IN2(r810_n254), .IN1(r810_n259), .Q(r810_n258) );
  NAND2X0 r810_U264 ( .IN1(r810_n257), .IN2(r810_n258), .QN(P1_N4385) );
  INVX0 r810_U263 ( .ZN(r810_n243), .INP(P1_N4234) );
  NAND2X0 r810_U262 ( .IN1(n7062), .IN2(r810_n243), .QN(r810_n255) );
  OR2X1 r810_U261 ( .IN2(n7062), .IN1(r810_n243), .Q(r810_n256) );
  NAND2X0 r810_U260 ( .IN1(r810_n255), .IN2(r810_n256), .QN(r810_n249) );
  NAND2X0 r810_U259 ( .IN1(P1_N5159), .IN2(r810_n254), .QN(r810_n250) );
  OR2X1 r810_U258 ( .IN2(P1_N5159), .IN1(r810_n254), .Q(r810_n252) );
  NAND2X0 r810_U257 ( .IN1(r810_n252), .IN2(r810_n253), .QN(r810_n251) );
  NAND2X0 r810_U256 ( .IN1(r810_n250), .IN2(r810_n251), .QN(r810_n244) );
  NAND2X0 r810_U255 ( .IN1(r810_n249), .IN2(r810_n244), .QN(r810_n247) );
  OR2X1 r810_U254 ( .IN2(r810_n244), .IN1(r810_n249), .Q(r810_n248) );
  NAND2X0 r810_U253 ( .IN1(r810_n247), .IN2(r810_n248), .QN(P1_N4386) );
  INVX0 r810_U252 ( .ZN(r810_n233), .INP(P1_N4235) );
  NAND2X0 r810_U251 ( .IN1(n7059), .IN2(r810_n233), .QN(r810_n245) );
  OR2X1 r810_U250 ( .IN2(n7059), .IN1(r810_n233), .Q(r810_n246) );
  NAND2X0 r810_U249 ( .IN1(r810_n245), .IN2(r810_n246), .QN(r810_n239) );
  NAND2X0 r810_U248 ( .IN1(n7062), .IN2(r810_n244), .QN(r810_n240) );
  OR2X1 r810_U247 ( .IN2(n7062), .IN1(r810_n244), .Q(r810_n242) );
  NAND2X0 r810_U246 ( .IN1(r810_n242), .IN2(r810_n243), .QN(r810_n241) );
  NAND2X0 r810_U245 ( .IN1(r810_n240), .IN2(r810_n241), .QN(r810_n234) );
  NAND2X0 r810_U244 ( .IN1(r810_n239), .IN2(r810_n234), .QN(r810_n237) );
  OR2X1 r810_U243 ( .IN2(r810_n234), .IN1(r810_n239), .Q(r810_n238) );
  NAND2X0 r810_U242 ( .IN1(r810_n237), .IN2(r810_n238), .QN(P1_N4387) );
  INVX0 r810_U241 ( .ZN(r810_n223), .INP(P1_N4236) );
  NAND2X0 r810_U240 ( .IN1(P1_N5162), .IN2(r810_n223), .QN(r810_n235) );
  OR2X1 r810_U239 ( .IN2(P1_N5162), .IN1(r810_n223), .Q(r810_n236) );
  NAND2X0 r810_U238 ( .IN1(r810_n235), .IN2(r810_n236), .QN(r810_n229) );
  NAND2X0 r810_U237 ( .IN1(n7059), .IN2(r810_n234), .QN(r810_n230) );
  OR2X1 r810_U236 ( .IN2(n7059), .IN1(r810_n234), .Q(r810_n232) );
  NAND2X0 r810_U235 ( .IN1(r810_n232), .IN2(r810_n233), .QN(r810_n231) );
  NAND2X0 r810_U234 ( .IN1(r810_n230), .IN2(r810_n231), .QN(r810_n224) );
  NAND2X0 r810_U233 ( .IN1(r810_n229), .IN2(r810_n224), .QN(r810_n227) );
  OR2X1 r810_U232 ( .IN2(r810_n224), .IN1(r810_n229), .Q(r810_n228) );
  NAND2X0 r810_U231 ( .IN1(r810_n227), .IN2(r810_n228), .QN(P1_N4388) );
  INVX0 r810_U230 ( .ZN(r810_n213), .INP(P1_N4237) );
  NAND2X0 r810_U229 ( .IN1(n7116), .IN2(r810_n213), .QN(r810_n225) );
  OR2X1 r810_U228 ( .IN2(P1_N5163), .IN1(r810_n213), .Q(r810_n226) );
  NAND2X0 r810_U227 ( .IN1(r810_n225), .IN2(r810_n226), .QN(r810_n219) );
  NAND2X0 r810_U226 ( .IN1(P1_N5162), .IN2(r810_n224), .QN(r810_n220) );
  OR2X1 r810_U225 ( .IN2(P1_N5162), .IN1(r810_n224), .Q(r810_n222) );
  NAND2X0 r810_U224 ( .IN1(r810_n222), .IN2(r810_n223), .QN(r810_n221) );
  NAND2X0 r810_U223 ( .IN1(r810_n220), .IN2(r810_n221), .QN(r810_n214) );
  NAND2X0 r810_U222 ( .IN1(r810_n219), .IN2(r810_n214), .QN(r810_n217) );
  OR2X1 r810_U221 ( .IN2(r810_n214), .IN1(r810_n219), .Q(r810_n218) );
  NAND2X0 r810_U220 ( .IN1(r810_n217), .IN2(r810_n218), .QN(P1_N4389) );
  INVX0 r810_U219 ( .ZN(r810_n203), .INP(P1_N4238) );
  NAND2X0 r810_U218 ( .IN1(P1_N5164), .IN2(r810_n203), .QN(r810_n215) );
  OR2X1 r810_U217 ( .IN2(P1_N5164), .IN1(r810_n203), .Q(r810_n216) );
  NAND2X0 r810_U216 ( .IN1(r810_n215), .IN2(r810_n216), .QN(r810_n209) );
  NAND2X0 r810_U215 ( .IN1(P1_N5163), .IN2(r810_n214), .QN(r810_n210) );
  OR2X1 r810_U214 ( .IN2(P1_N5163), .IN1(r810_n214), .Q(r810_n212) );
  INVX0 r810_U321 ( .ZN(r810_n291), .INP(P1_N4223) );
  NOR2X0 r810_U320 ( .QN(r810_n287), .IN1(r810_n291), .IN2(n7034) );
  INVX0 r810_U319 ( .ZN(r810_n162), .INP(r810_n287) );
  NAND2X0 r810_U318 ( .IN1(n7034), .IN2(r810_n291), .QN(r810_n290) );
  NAND2X0 r810_U317 ( .IN1(r810_n162), .IN2(r810_n290), .QN(P1_N4375) );
  INVX0 r810_U316 ( .ZN(r810_n253), .INP(P1_N4233) );
  NAND2X0 r810_U315 ( .IN1(P1_N5159), .IN2(r810_n253), .QN(r810_n288) );
  OR2X1 r810_U314 ( .IN2(P1_N5159), .IN1(r810_n253), .Q(r810_n289) );
  NAND2X0 r810_U313 ( .IN1(r810_n288), .IN2(r810_n289), .QN(r810_n259) );
  NAND2X0 r810_U312 ( .IN1(P1_N5150), .IN2(r810_n162), .QN(r810_n284) );
  NAND2X0 r810_U310 ( .IN1(r810_n287), .IN2(n7048), .QN(r810_n286) );
  INVX0 r810_U309 ( .ZN(r810_n166), .INP(P1_N4224) );
  NAND2X0 r810_U308 ( .IN1(r810_n286), .IN2(r810_n166), .QN(r810_n285) );
  NAND2X0 r810_U307 ( .IN1(r810_n284), .IN2(r810_n285), .QN(r810_n53) );
  NAND2X0 r812_U90 ( .IN1(r812_n79), .IN2(r812_n80), .QN(P1_N4576) );
  NAND2X0 r812_U89 ( .IN1(P1_N5150), .IN2(P1_N4556), .QN(r812_n78) );
  OR2X1 r812_U88 ( .IN2(n7046), .IN1(r812_n78), .Q(r812_n76) );
  NAND2X0 r812_U87 ( .IN1(n7046), .IN2(r812_n78), .QN(r812_n77) );
  NAND2X0 r812_U86 ( .IN1(r812_n76), .IN2(r812_n77), .QN(P1_N4558) );
  NOR2X0 r812_U85 ( .QN(r812_n73), .IN1(r812_n74), .IN2(r812_n135) );
  NAND2X0 r812_U84 ( .IN1(r812_n73), .IN2(n7096), .QN(r812_n66) );
  OR2X1 r812_U83 ( .IN2(n7093), .IN1(r812_n66), .Q(r812_n71) );
  NAND2X0 r812_U82 ( .IN1(n7093), .IN2(r812_n66), .QN(r812_n72) );
  NAND2X0 r812_U81 ( .IN1(r812_n71), .IN2(r812_n72), .QN(P1_N4577) );
  OR2X1 r812_U79 ( .IN2(r812_n66), .IN1(r812_n131), .Q(r812_n70) );
  OR2X1 r812_U78 ( .IN2(P1_N5171), .IN1(r812_n70), .Q(r812_n68) );
  NAND2X0 r812_U77 ( .IN1(P1_N5171), .IN2(r812_n70), .QN(r812_n69) );
  NAND2X0 r812_U76 ( .IN1(r812_n68), .IN2(r812_n69), .QN(P1_N4578) );
  NOR2X0 r812_U75 ( .QN(r812_n65), .IN1(r812_n66), .IN2(r812_n131) );
  NAND2X0 r812_U74 ( .IN1(r812_n65), .IN2(P1_N5171), .QN(r812_n58) );
  OR2X1 r812_U73 ( .IN2(n7141), .IN1(r812_n58), .Q(r812_n63) );
  NAND2X0 r812_U72 ( .IN1(n7141), .IN2(r812_n58), .QN(r812_n64) );
  NAND2X0 r812_U71 ( .IN1(r812_n63), .IN2(r812_n64), .QN(P1_N4579) );
  OR2X1 r812_U69 ( .IN2(r812_n58), .IN1(n7144), .Q(r812_n62) );
  OR2X1 r812_U68 ( .IN2(P1_N5173), .IN1(r812_n62), .Q(r812_n60) );
  NAND2X0 r812_U67 ( .IN1(P1_N5173), .IN2(r812_n62), .QN(r812_n61) );
  NAND2X0 r812_U66 ( .IN1(r812_n60), .IN2(r812_n61), .QN(P1_N4580) );
  NOR2X0 r812_U65 ( .QN(r812_n57), .IN1(r812_n58), .IN2(n7144) );
  NAND2X0 r812_U64 ( .IN1(r812_n57), .IN2(P1_N5173), .QN(r812_n50) );
  OR2X1 r812_U63 ( .IN2(n7129), .IN1(r812_n50), .Q(r812_n55) );
  NAND2X0 r812_U62 ( .IN1(n7129), .IN2(r812_n50), .QN(r812_n56) );
  NAND2X0 r812_U61 ( .IN1(r812_n55), .IN2(r812_n56), .QN(P1_N4581) );
  OR2X1 r812_U59 ( .IN2(r812_n50), .IN1(n7130), .Q(r812_n54) );
  OR2X1 r812_U58 ( .IN2(P1_N5175), .IN1(r812_n54), .Q(r812_n52) );
  NAND2X0 r812_U57 ( .IN1(P1_N5175), .IN2(r812_n54), .QN(r812_n53) );
  NAND2X0 r812_U56 ( .IN1(r812_n52), .IN2(r812_n53), .QN(P1_N4582) );
  NOR2X0 r812_U55 ( .QN(r812_n49), .IN1(r812_n50), .IN2(n7130) );
  NAND2X0 r812_U54 ( .IN1(r812_n49), .IN2(P1_N5175), .QN(r812_n42) );
  OR2X1 r812_U53 ( .IN2(n7122), .IN1(r812_n42), .Q(r812_n47) );
  NAND2X0 r812_U52 ( .IN1(n7122), .IN2(r812_n42), .QN(r812_n48) );
  NAND2X0 r812_U51 ( .IN1(r812_n47), .IN2(r812_n48), .QN(P1_N4583) );
  OR2X1 r812_U49 ( .IN2(r812_n42), .IN1(n7119), .Q(r812_n46) );
  OR2X1 r812_U48 ( .IN2(P1_N5177), .IN1(r812_n46), .Q(r812_n44) );
  NAND2X0 r812_U47 ( .IN1(P1_N5177), .IN2(r812_n46), .QN(r812_n45) );
  NAND2X0 r812_U46 ( .IN1(r812_n44), .IN2(r812_n45), .QN(P1_N4584) );
  NOR2X0 r812_U45 ( .QN(r812_n41), .IN1(r812_n42), .IN2(n7119) );
  NAND2X0 r812_U44 ( .IN1(r812_n41), .IN2(P1_N5177), .QN(r812_n32) );
  OR2X1 r812_U43 ( .IN2(P1_N5178), .IN1(r812_n32), .Q(r812_n39) );
  NAND2X0 r812_U42 ( .IN1(P1_N5178), .IN2(r812_n32), .QN(r812_n40) );
  NAND2X0 r812_U41 ( .IN1(r812_n39), .IN2(r812_n40), .QN(P1_N4585) );
  OR2X1 r812_U39 ( .IN2(r812_n32), .IN1(n7146), .Q(r812_n38) );
  OR2X1 r812_U38 ( .IN2(P1_N497), .IN1(r812_n38), .Q(r812_n36) );
  NAND2X0 r812_U37 ( .IN1(P1_N497), .IN2(r812_n38), .QN(r812_n37) );
  NAND2X0 r812_U36 ( .IN1(r812_n36), .IN2(r812_n37), .QN(P1_N4586) );
  OR2X1 r812_U35 ( .IN2(n7041), .IN1(r812_n26), .Q(r812_n34) );
  NAND2X0 r812_U34 ( .IN1(n7041), .IN2(r812_n26), .QN(r812_n35) );
  NAND2X0 r812_U33 ( .IN1(r812_n34), .IN2(r812_n35), .QN(P1_N4559) );
  NOR2X0 r812_U31 ( .QN(r812_n31), .IN1(r812_n32), .IN2(n7146) );
  AND2X1 r812_U30 ( .IN1(r812_n31), .IN2(P1_N497), .Q(r812_n29) );
  NOR2X0 r812_U29 ( .QN(P1_N4588), .IN1(n4469), .IN2(r812_n29) );
  INVX0 r812_U28 ( .ZN(r812_n27), .INP(P1_N4588) );
  NAND2X0 r812_U27 ( .IN1(r812_n29), .IN2(n4469), .QN(r812_n28) );
  NAND2X0 r812_U26 ( .IN1(r812_n27), .IN2(r812_n28), .QN(P1_N4587) );
  OR2X1 r812_U25 ( .IN2(r812_n26), .IN1(r812_n18), .Q(r812_n24) );
  OR2X1 r812_U24 ( .IN2(P1_N5153), .IN1(r812_n24), .Q(r812_n22) );
  NAND2X0 r812_U23 ( .IN1(P1_N5153), .IN2(r812_n24), .QN(r812_n23) );
  NAND2X0 r812_U22 ( .IN1(r812_n22), .IN2(r812_n23), .QN(P1_N4560) );
  OR2X1 r812_U21 ( .IN2(n7081), .IN1(r812_n19), .Q(r812_n20) );
  NAND2X0 r812_U20 ( .IN1(n7081), .IN2(r812_n19), .QN(r812_n21) );
  NAND2X0 r812_U19 ( .IN1(r812_n20), .IN2(r812_n21), .QN(P1_N4561) );
  OR2X1 r812_U18 ( .IN2(r812_n19), .IN1(r812_n128), .Q(r812_n17) );
  OR2X1 r812_U17 ( .IN2(n7080), .IN1(r812_n17), .Q(r812_n15) );
  NAND2X0 r812_U16 ( .IN1(n7080), .IN2(r812_n17), .QN(r812_n16) );
  NAND2X0 r812_U15 ( .IN1(r812_n15), .IN2(r812_n16), .QN(P1_N4562) );
  OR2X1 r812_U14 ( .IN2(P1_N5156), .IN1(r812_n12), .Q(r812_n13) );
  NAND2X0 r812_U13 ( .IN1(P1_N5156), .IN2(r812_n12), .QN(r812_n14) );
  NAND2X0 r812_U12 ( .IN1(r812_n13), .IN2(r812_n14), .QN(P1_N4563) );
  OR2X1 r812_U11 ( .IN2(r812_n12), .IN1(r812_n125), .Q(r812_n10) );
  OR2X1 r812_U10 ( .IN2(n7072), .IN1(r812_n10), .Q(r812_n8) );
  NAND2X0 r812_U9 ( .IN1(n7072), .IN2(r812_n10), .QN(r812_n9) );
  NAND2X0 r812_U8 ( .IN1(r812_n8), .IN2(r812_n9), .QN(P1_N4564) );
  OR2X1 r812_U7 ( .IN2(n7070), .IN1(r812_n5), .Q(r812_n6) );
  NAND2X0 r812_U6 ( .IN1(n7070), .IN2(r812_n5), .QN(r812_n7) );
  NAND2X0 r812_U5 ( .IN1(r812_n6), .IN2(r812_n7), .QN(P1_N4565) );
  OR2X1 r812_U4 ( .IN2(r812_n5), .IN1(n7071), .Q(r812_n3) );
  OR2X1 r812_U3 ( .IN2(n7066), .IN1(r812_n3), .Q(r812_n1) );
  NAND2X0 r812_U2 ( .IN1(n7066), .IN2(r812_n3), .QN(r812_n2) );
  NAND2X0 r812_U1 ( .IN1(r812_n1), .IN2(r812_n2), .QN(P1_N4566) );
  NAND2X0 r812_U155 ( .IN1(P1_N4556), .IN2(r812_n33), .QN(r812_n123) );
  INVX0 r812_U154 ( .ZN(r812_n121), .INP(P1_N4556) );
  NAND2X0 r812_U153 ( .IN1(P1_N5150), .IN2(r812_n121), .QN(r812_n124) );
  NAND2X0 r812_U152 ( .IN1(r812_n123), .IN2(r812_n124), .QN(P1_N4557) );
  NOR2X0 r812_U151 ( .QN(r812_n120), .IN1(r812_n121), .IN2(r812_n33) );
  NAND2X0 r812_U150 ( .IN1(r812_n120), .IN2(n7046), .QN(r812_n26) );
  NOR2X0 r812_U148 ( .QN(r812_n119), .IN1(r812_n26), .IN2(r812_n18) );
  NAND2X0 r812_U147 ( .IN1(r812_n119), .IN2(P1_N5153), .QN(r812_n19) );
  NOR2X0 r812_U145 ( .QN(r812_n118), .IN1(r812_n19), .IN2(r812_n128) );
  NAND2X0 r812_U144 ( .IN1(r812_n118), .IN2(n7080), .QN(r812_n12) );
  NOR2X0 r812_U142 ( .QN(r812_n117), .IN1(r812_n12), .IN2(r812_n125) );
  NAND2X0 r812_U141 ( .IN1(r812_n117), .IN2(n7072), .QN(r812_n5) );
  NOR2X0 r812_U139 ( .QN(r812_n116), .IN1(r812_n5), .IN2(n7071) );
  NAND2X0 r812_U138 ( .IN1(r812_n116), .IN2(n7066), .QN(r812_n109) );
  OR2X1 r812_U137 ( .IN2(n7062), .IN1(r812_n109), .Q(r812_n114) );
  NAND2X0 r812_U136 ( .IN1(n7062), .IN2(r812_n109), .QN(r812_n115) );
  NAND2X0 r812_U135 ( .IN1(r812_n114), .IN2(r812_n115), .QN(P1_N4567) );
  OR2X1 r812_U133 ( .IN2(r812_n109), .IN1(n7063), .Q(r812_n113) );
  OR2X1 r812_U132 ( .IN2(n7059), .IN1(r812_n113), .Q(r812_n111) );
  NAND2X0 r812_U131 ( .IN1(n7059), .IN2(r812_n113), .QN(r812_n112) );
  NAND2X0 r812_U130 ( .IN1(r812_n111), .IN2(r812_n112), .QN(P1_N4568) );
  NOR2X0 r812_U129 ( .QN(r812_n108), .IN1(r812_n109), .IN2(n7063) );
  NAND2X0 r812_U128 ( .IN1(r812_n108), .IN2(n7059), .QN(r812_n101) );
  OR2X1 r812_U127 ( .IN2(n7055), .IN1(r812_n101), .Q(r812_n106) );
  NAND2X0 r812_U126 ( .IN1(n7055), .IN2(r812_n101), .QN(r812_n107) );
  NAND2X0 r812_U125 ( .IN1(r812_n106), .IN2(r812_n107), .QN(P1_N4569) );
  OR2X1 r812_U123 ( .IN2(r812_n101), .IN1(n7056), .Q(r812_n105) );
  OR2X1 r812_U122 ( .IN2(n7116), .IN1(r812_n105), .Q(r812_n103) );
  NAND2X0 r812_U121 ( .IN1(n7116), .IN2(r812_n105), .QN(r812_n104) );
  NAND2X0 r812_U120 ( .IN1(r812_n103), .IN2(r812_n104), .QN(P1_N4570) );
  NOR2X0 r812_U119 ( .QN(r812_n100), .IN1(r812_n101), .IN2(n7056) );
  NAND2X0 r812_U118 ( .IN1(r812_n100), .IN2(n7116), .QN(r812_n93) );
  OR2X1 r812_U117 ( .IN2(n7113), .IN1(r812_n93), .Q(r812_n98) );
  NAND2X0 r812_U116 ( .IN1(n7113), .IN2(r812_n93), .QN(r812_n99) );
  NAND2X0 r812_U115 ( .IN1(r812_n98), .IN2(r812_n99), .QN(P1_N4571) );
  OR2X1 r812_U113 ( .IN2(r812_n93), .IN1(r812_n141), .Q(r812_n97) );
  OR2X1 r812_U112 ( .IN2(n7110), .IN1(r812_n97), .Q(r812_n95) );
  NAND2X0 r812_U111 ( .IN1(n7110), .IN2(r812_n97), .QN(r812_n96) );
  NAND2X0 r812_U110 ( .IN1(r812_n95), .IN2(r812_n96), .QN(P1_N4572) );
  NOR2X0 r812_U109 ( .QN(r812_n92), .IN1(r812_n93), .IN2(r812_n141) );
  NAND2X0 r812_U108 ( .IN1(r812_n92), .IN2(n7110), .QN(r812_n85) );
  OR2X1 r812_U107 ( .IN2(n7106), .IN1(r812_n85), .Q(r812_n90) );
  NAND2X0 r812_U106 ( .IN1(n7106), .IN2(r812_n85), .QN(r812_n91) );
  NAND2X0 r812_U105 ( .IN1(r812_n90), .IN2(r812_n91), .QN(P1_N4573) );
  OR2X1 r812_U103 ( .IN2(r812_n85), .IN1(r812_n138), .Q(r812_n89) );
  OR2X1 r812_U102 ( .IN2(n7103), .IN1(r812_n89), .Q(r812_n87) );
  NAND2X0 r812_U101 ( .IN1(n7103), .IN2(r812_n89), .QN(r812_n88) );
  NAND2X0 r812_U100 ( .IN1(r812_n87), .IN2(r812_n88), .QN(P1_N4574) );
  NOR2X0 r812_U99 ( .QN(r812_n84), .IN1(r812_n85), .IN2(r812_n138) );
  NAND2X0 r812_U98 ( .IN1(r812_n84), .IN2(n7103), .QN(r812_n74) );
  OR2X1 r812_U97 ( .IN2(n7099), .IN1(r812_n74), .Q(r812_n82) );
  NAND2X0 r812_U96 ( .IN1(n7099), .IN2(r812_n74), .QN(r812_n83) );
  NAND2X0 r812_U95 ( .IN1(r812_n82), .IN2(r812_n83), .QN(P1_N4575) );
  OR2X1 r812_U93 ( .IN2(r812_n74), .IN1(r812_n135), .Q(r812_n81) );
  OR2X1 r812_U92 ( .IN2(P1_N5169), .IN1(r812_n81), .Q(r812_n79) );
  NAND2X0 r812_U91 ( .IN1(P1_N5169), .IN2(r812_n81), .QN(r812_n80) );
  INVX0 r812_U32 ( .ZN(r812_n18), .INP(n7041) );
  INVX0 r812_U40 ( .ZN(r812_n33), .INP(P1_N5150) );
  INVX0 r812_U50 ( .ZN(r812_n125), .INP(P1_N5156) );
  INVX0 r812_U60 ( .ZN(r812_n128), .INP(n7081) );
  INVX0 r812_U70 ( .ZN(r812_n131), .INP(n7093) );
  INVX0 r812_U80 ( .ZN(r812_n135), .INP(n7099) );
  INVX0 r812_U94 ( .ZN(r812_n138), .INP(n7106) );
  INVX0 r812_U104 ( .ZN(r812_n141), .INP(n7113) );
  NAND2X0 r816_U79 ( .IN1(r816_n140), .IN2(r816_n8), .QN(r816_n138) );
  NAND2X0 r816_U78 ( .IN1(r816_n138), .IN2(r816_n139), .QN(r816_n136) );
  NAND2X0 r816_U77 ( .IN1(P1_N5115), .IN2(n4469), .QN(r816_n1) );
  NAND2X0 r816_U76 ( .IN1(r816_n136), .IN2(r816_n1), .QN(r816_n135) );
  NAND2X0 r816_U75 ( .IN1(r816_n4), .IN2(r816_n135), .QN(P1_N5137) );
  NOR2X0 r816_U74 ( .QN(r816_n20), .IN1(r816_n133), .IN2(r816_n134) );
  NOR2X0 r816_U73 ( .QN(r816_n35), .IN1(r816_n131), .IN2(r816_n132) );
  NOR2X0 r816_U72 ( .QN(r816_n50), .IN1(r816_n129), .IN2(r816_n130) );
  NOR2X0 r816_U71 ( .QN(r816_n65), .IN1(r816_n127), .IN2(r816_n128) );
  NOR2X0 r816_U70 ( .QN(r816_n80), .IN1(r816_n125), .IN2(r816_n126) );
  NOR2X0 r816_U69 ( .QN(r816_n95), .IN1(r816_n123), .IN2(r816_n124) );
  NOR2X0 r816_U68 ( .QN(r816_n110), .IN1(r816_n121), .IN2(r816_n122) );
  NAND2X0 r816_U67 ( .IN1(n7034), .IN2(r816_n120), .QN(r816_n117) );
  NOR2X0 r816_U66 ( .QN(r816_n118), .IN1(n7051), .IN2(r816_n117) );
  INVX0 r816_U65 ( .ZN(r816_n119), .INP(P1_N5085) );
  NOR2X0 r816_U64 ( .QN(r816_n114), .IN1(r816_n118), .IN2(r816_n119) );
  AND2X1 r816_U63 ( .IN1(n7051), .IN2(r816_n117), .Q(r816_n115) );
  NOR2X0 r816_U62 ( .QN(r816_n112), .IN1(r816_n114), .IN2(r816_n115) );
  NAND2X0 r816_U61 ( .IN1(r816_n112), .IN2(r816_n113), .QN(r816_n111) );
  NAND2X0 r816_U60 ( .IN1(r816_n110), .IN2(r816_n111), .QN(r816_n108) );
  NAND2X0 r816_U59 ( .IN1(r816_n108), .IN2(r816_n109), .QN(r816_n107) );
  NOR2X0 r816_U58 ( .QN(r816_n101), .IN1(r816_n106), .IN2(r816_n107) );
  INVX0 r816_U57 ( .ZN(r816_n103), .INP(r816_n105) );
  NAND2X0 r816_U56 ( .IN1(r816_n103), .IN2(r816_n104), .QN(r816_n102) );
  NOR2X0 r816_U55 ( .QN(r816_n100), .IN1(r816_n101), .IN2(r816_n102) );
  NOR2X0 r816_U54 ( .QN(r816_n97), .IN1(r816_n99), .IN2(r816_n100) );
  NAND2X0 r816_U53 ( .IN1(r816_n97), .IN2(r816_n98), .QN(r816_n96) );
  NAND2X0 r816_U52 ( .IN1(r816_n95), .IN2(r816_n96), .QN(r816_n93) );
  NAND2X0 r816_U51 ( .IN1(r816_n93), .IN2(r816_n94), .QN(r816_n92) );
  NOR2X0 r816_U50 ( .QN(r816_n86), .IN1(r816_n91), .IN2(r816_n92) );
  INVX0 r816_U49 ( .ZN(r816_n88), .INP(r816_n90) );
  NAND2X0 r816_U48 ( .IN1(r816_n88), .IN2(r816_n89), .QN(r816_n87) );
  NOR2X0 r816_U47 ( .QN(r816_n85), .IN1(r816_n86), .IN2(r816_n87) );
  NOR2X0 r816_U46 ( .QN(r816_n82), .IN1(r816_n84), .IN2(r816_n85) );
  NAND2X0 r816_U45 ( .IN1(r816_n82), .IN2(r816_n83), .QN(r816_n81) );
  NAND2X0 r816_U44 ( .IN1(r816_n80), .IN2(r816_n81), .QN(r816_n78) );
  NAND2X0 r816_U43 ( .IN1(r816_n78), .IN2(r816_n79), .QN(r816_n77) );
  NOR2X0 r816_U42 ( .QN(r816_n71), .IN1(r816_n76), .IN2(r816_n77) );
  INVX0 r816_U41 ( .ZN(r816_n73), .INP(r816_n75) );
  NAND2X0 r816_U40 ( .IN1(r816_n73), .IN2(r816_n74), .QN(r816_n72) );
  NOR2X0 r816_U39 ( .QN(r816_n70), .IN1(r816_n71), .IN2(r816_n72) );
  NOR2X0 r816_U38 ( .QN(r816_n67), .IN1(r816_n69), .IN2(r816_n70) );
  NAND2X0 r816_U37 ( .IN1(r816_n67), .IN2(r816_n68), .QN(r816_n66) );
  NAND2X0 r816_U36 ( .IN1(r816_n65), .IN2(r816_n66), .QN(r816_n63) );
  NAND2X0 r816_U35 ( .IN1(r816_n63), .IN2(r816_n64), .QN(r816_n62) );
  NOR2X0 r816_U34 ( .QN(r816_n56), .IN1(r816_n61), .IN2(r816_n62) );
  INVX0 r816_U33 ( .ZN(r816_n58), .INP(r816_n60) );
  NAND2X0 r816_U32 ( .IN1(r816_n58), .IN2(r816_n59), .QN(r816_n57) );
  NOR2X0 r816_U31 ( .QN(r816_n55), .IN1(r816_n56), .IN2(r816_n57) );
  NOR2X0 r816_U30 ( .QN(r816_n52), .IN1(r816_n54), .IN2(r816_n55) );
  NAND2X0 r816_U29 ( .IN1(r816_n52), .IN2(r816_n53), .QN(r816_n51) );
  NAND2X0 r816_U28 ( .IN1(r816_n50), .IN2(r816_n51), .QN(r816_n48) );
  NAND2X0 r816_U27 ( .IN1(r816_n48), .IN2(r816_n49), .QN(r816_n47) );
  NOR2X0 r816_U26 ( .QN(r816_n41), .IN1(r816_n46), .IN2(r816_n47) );
  INVX0 r816_U25 ( .ZN(r816_n43), .INP(r816_n45) );
  NAND2X0 r816_U24 ( .IN1(r816_n43), .IN2(r816_n44), .QN(r816_n42) );
  NOR2X0 r816_U23 ( .QN(r816_n40), .IN1(r816_n41), .IN2(r816_n42) );
  NOR2X0 r816_U22 ( .QN(r816_n37), .IN1(r816_n39), .IN2(r816_n40) );
  NAND2X0 r816_U21 ( .IN1(r816_n37), .IN2(r816_n38), .QN(r816_n36) );
  NAND2X0 r816_U20 ( .IN1(r816_n35), .IN2(r816_n36), .QN(r816_n33) );
  NAND2X0 r816_U19 ( .IN1(r816_n33), .IN2(r816_n34), .QN(r816_n32) );
  NOR2X0 r816_U18 ( .QN(r816_n26), .IN1(r816_n31), .IN2(r816_n32) );
  INVX0 r816_U17 ( .ZN(r816_n28), .INP(r816_n30) );
  NAND2X0 r816_U16 ( .IN1(r816_n28), .IN2(r816_n29), .QN(r816_n27) );
  NOR2X0 r816_U15 ( .QN(r816_n25), .IN1(r816_n26), .IN2(r816_n27) );
  NOR2X0 r816_U14 ( .QN(r816_n22), .IN1(r816_n24), .IN2(r816_n25) );
  NAND2X0 r816_U13 ( .IN1(r816_n22), .IN2(r816_n23), .QN(r816_n21) );
  NAND2X0 r816_U12 ( .IN1(r816_n20), .IN2(r816_n21), .QN(r816_n18) );
  NAND2X0 r816_U11 ( .IN1(r816_n18), .IN2(r816_n19), .QN(r816_n17) );
  NOR2X0 r816_U10 ( .QN(r816_n11), .IN1(r816_n16), .IN2(r816_n17) );
  INVX0 r816_U9 ( .ZN(r816_n13), .INP(r816_n15) );
  NAND2X0 r816_U8 ( .IN1(r816_n13), .IN2(r816_n14), .QN(r816_n12) );
  NOR2X0 r816_U7 ( .QN(r816_n10), .IN1(r816_n11), .IN2(r816_n12) );
  NOR2X0 r816_U6 ( .QN(r816_n7), .IN1(r816_n9), .IN2(r816_n10) );
  NAND2X0 r816_U5 ( .IN1(r816_n7), .IN2(r816_n8), .QN(r816_n5) );
  NAND2X0 r816_U4 ( .IN1(r816_n5), .IN2(r816_n6), .QN(r816_n3) );
  NAND2X0 r816_U3 ( .IN1(r816_n3), .IN2(r816_n4), .QN(r816_n2) );
  NAND2X0 r816_U2 ( .IN1(r816_n1), .IN2(r816_n2), .QN(P1_N5143) );
  NOR2X0 r816_U1 ( .QN(P1_N5140), .IN1(P1_N5137), .IN2(P1_N5143) );
  NAND2X0 r816_U172 ( .IN1(P1_N5094), .IN2(n7067), .QN(r816_n214) );
  INVX0 r816_U171 ( .ZN(r816_n216), .INP(r816_n214) );
  NOR2X0 r816_U170 ( .QN(r816_n83), .IN1(r816_n125), .IN2(r816_n216) );
  NAND2X0 r816_U169 ( .IN1(r816_n215), .IN2(r816_n83), .QN(r816_n213) );
  NAND2X0 r816_U168 ( .IN1(r816_n213), .IN2(r816_n214), .QN(r816_n212) );
  NOR2X0 r816_U167 ( .QN(r816_n210), .IN1(r816_n211), .IN2(r816_n212) );
  NOR2X0 r816_U166 ( .QN(r816_n207), .IN1(r816_n126), .IN2(r816_n210) );
  OR2X1 r816_U164 ( .IN2(P1_N5096), .IN1(n7058), .Q(r816_n74) );
  NAND2X0 r816_U163 ( .IN1(P1_N5096), .IN2(n7058), .QN(r816_n206) );
  NAND2X0 r816_U162 ( .IN1(r816_n74), .IN2(r816_n206), .QN(r816_n76) );
  INVX0 r816_U161 ( .ZN(r816_n208), .INP(r816_n76) );
  NAND2X0 r816_U160 ( .IN1(r816_n207), .IN2(r816_n208), .QN(r816_n205) );
  NAND2X0 r816_U159 ( .IN1(r816_n205), .IN2(r816_n206), .QN(r816_n204) );
  NOR2X0 r816_U158 ( .QN(r816_n203), .IN1(r816_n69), .IN2(r816_n204) );
  NOR2X0 r816_U157 ( .QN(r816_n200), .IN1(r816_n75), .IN2(r816_n203) );
  NOR2X0 r816_U155 ( .QN(r816_n127), .IN1(n7115), .IN2(P1_N5098) );
  NAND2X0 r816_U154 ( .IN1(P1_N5098), .IN2(n7115), .QN(r816_n199) );
  INVX0 r816_U153 ( .ZN(r816_n201), .INP(r816_n199) );
  NOR2X0 r816_U152 ( .QN(r816_n68), .IN1(r816_n127), .IN2(r816_n201) );
  NAND2X0 r816_U151 ( .IN1(r816_n200), .IN2(r816_n68), .QN(r816_n198) );
  NAND2X0 r816_U150 ( .IN1(r816_n198), .IN2(r816_n199), .QN(r816_n197) );
  NOR2X0 r816_U149 ( .QN(r816_n195), .IN1(r816_n196), .IN2(r816_n197) );
  NOR2X0 r816_U148 ( .QN(r816_n192), .IN1(r816_n128), .IN2(r816_n195) );
  OR2X1 r816_U146 ( .IN2(P1_N5100), .IN1(n7109), .Q(r816_n59) );
  NAND2X0 r816_U145 ( .IN1(P1_N5100), .IN2(n7109), .QN(r816_n191) );
  NAND2X0 r816_U144 ( .IN1(r816_n59), .IN2(r816_n191), .QN(r816_n61) );
  INVX0 r816_U143 ( .ZN(r816_n193), .INP(r816_n61) );
  NAND2X0 r816_U142 ( .IN1(r816_n192), .IN2(r816_n193), .QN(r816_n190) );
  NAND2X0 r816_U141 ( .IN1(r816_n190), .IN2(r816_n191), .QN(r816_n189) );
  NOR2X0 r816_U140 ( .QN(r816_n188), .IN1(r816_n54), .IN2(r816_n189) );
  NOR2X0 r816_U139 ( .QN(r816_n185), .IN1(r816_n60), .IN2(r816_n188) );
  NOR2X0 r816_U137 ( .QN(r816_n129), .IN1(n7102), .IN2(P1_N5102) );
  NAND2X0 r816_U136 ( .IN1(P1_N5102), .IN2(n7102), .QN(r816_n184) );
  INVX0 r816_U135 ( .ZN(r816_n186), .INP(r816_n184) );
  NOR2X0 r816_U134 ( .QN(r816_n53), .IN1(r816_n129), .IN2(r816_n186) );
  NAND2X0 r816_U133 ( .IN1(r816_n185), .IN2(r816_n53), .QN(r816_n183) );
  NAND2X0 r816_U132 ( .IN1(r816_n183), .IN2(r816_n184), .QN(r816_n182) );
  NOR2X0 r816_U131 ( .QN(r816_n180), .IN1(r816_n181), .IN2(r816_n182) );
  NOR2X0 r816_U130 ( .QN(r816_n177), .IN1(r816_n130), .IN2(r816_n180) );
  OR2X1 r816_U128 ( .IN2(P1_N5104), .IN1(n7095), .Q(r816_n44) );
  NAND2X0 r816_U127 ( .IN1(P1_N5104), .IN2(n7095), .QN(r816_n176) );
  NAND2X0 r816_U126 ( .IN1(r816_n44), .IN2(r816_n176), .QN(r816_n46) );
  INVX0 r816_U125 ( .ZN(r816_n178), .INP(r816_n46) );
  NAND2X0 r816_U124 ( .IN1(r816_n177), .IN2(r816_n178), .QN(r816_n175) );
  NAND2X0 r816_U123 ( .IN1(r816_n175), .IN2(r816_n176), .QN(r816_n174) );
  NOR2X0 r816_U122 ( .QN(r816_n173), .IN1(r816_n39), .IN2(r816_n174) );
  NOR2X0 r816_U121 ( .QN(r816_n170), .IN1(r816_n45), .IN2(r816_n173) );
  NOR2X0 r816_U119 ( .QN(r816_n131), .IN1(n7090), .IN2(P1_N5106) );
  NAND2X0 r816_U118 ( .IN1(P1_N5106), .IN2(n7090), .QN(r816_n169) );
  INVX0 r816_U117 ( .ZN(r816_n171), .INP(r816_n169) );
  NOR2X0 r816_U116 ( .QN(r816_n38), .IN1(r816_n131), .IN2(r816_n171) );
  NAND2X0 r816_U115 ( .IN1(r816_n170), .IN2(r816_n38), .QN(r816_n168) );
  NAND2X0 r816_U114 ( .IN1(r816_n168), .IN2(r816_n169), .QN(r816_n167) );
  NOR2X0 r816_U113 ( .QN(r816_n165), .IN1(r816_n166), .IN2(r816_n167) );
  NOR2X0 r816_U112 ( .QN(r816_n162), .IN1(r816_n132), .IN2(r816_n165) );
  OR2X1 r816_U110 ( .IN2(P1_N5108), .IN1(r816_n304), .Q(r816_n29) );
  NAND2X0 r816_U109 ( .IN1(P1_N5108), .IN2(r816_n304), .QN(r816_n161) );
  NAND2X0 r816_U108 ( .IN1(r816_n29), .IN2(r816_n161), .QN(r816_n31) );
  INVX0 r816_U107 ( .ZN(r816_n163), .INP(r816_n31) );
  NAND2X0 r816_U106 ( .IN1(r816_n162), .IN2(r816_n163), .QN(r816_n160) );
  NAND2X0 r816_U105 ( .IN1(r816_n160), .IN2(r816_n161), .QN(r816_n159) );
  NOR2X0 r816_U104 ( .QN(r816_n158), .IN1(r816_n24), .IN2(r816_n159) );
  NOR2X0 r816_U103 ( .QN(r816_n155), .IN1(r816_n30), .IN2(r816_n158) );
  NOR2X0 r816_U101 ( .QN(r816_n133), .IN1(r816_n301), .IN2(P1_N5110) );
  NAND2X0 r816_U100 ( .IN1(P1_N5110), .IN2(r816_n301), .QN(r816_n154) );
  INVX0 r816_U99 ( .ZN(r816_n156), .INP(r816_n154) );
  NOR2X0 r816_U98 ( .QN(r816_n23), .IN1(r816_n133), .IN2(r816_n156) );
  NAND2X0 r816_U97 ( .IN1(r816_n155), .IN2(r816_n23), .QN(r816_n153) );
  NAND2X0 r816_U96 ( .IN1(r816_n153), .IN2(r816_n154), .QN(r816_n152) );
  NOR2X0 r816_U95 ( .QN(r816_n150), .IN1(r816_n151), .IN2(r816_n152) );
  NOR2X0 r816_U94 ( .QN(r816_n147), .IN1(r816_n134), .IN2(r816_n150) );
  OR2X1 r816_U92 ( .IN2(P1_N5112), .IN1(n7117), .Q(r816_n14) );
  NAND2X0 r816_U91 ( .IN1(P1_N5112), .IN2(n7117), .QN(r816_n146) );
  NAND2X0 r816_U90 ( .IN1(r816_n14), .IN2(r816_n146), .QN(r816_n16) );
  INVX0 r816_U89 ( .ZN(r816_n148), .INP(r816_n16) );
  NAND2X0 r816_U88 ( .IN1(r816_n147), .IN2(r816_n148), .QN(r816_n145) );
  NAND2X0 r816_U87 ( .IN1(r816_n145), .IN2(r816_n146), .QN(r816_n144) );
  NOR2X0 r816_U86 ( .QN(r816_n143), .IN1(r816_n9), .IN2(r816_n144) );
  NOR2X0 r816_U85 ( .QN(r816_n140), .IN1(r816_n15), .IN2(r816_n143) );
  NAND2X0 r816_U83 ( .IN1(P1_N497), .IN2(r816_n308), .QN(r816_n6) );
  NAND2X0 r816_U81 ( .IN1(P1_N5114), .IN2(n7145), .QN(r816_n139) );
  AND2X1 r816_U80 ( .IN1(r816_n6), .IN2(r816_n139), .Q(r816_n8) );
  NOR2X0 r816_U265 ( .QN(r816_n15), .IN1(n7146), .IN2(P1_N5113) );
  AND2X1 r816_U264 ( .IN1(P1_N5113), .IN2(n7146), .Q(r816_n9) );
  NOR2X0 r816_U262 ( .QN(r816_n134), .IN1(n7119), .IN2(P1_N5111) );
  NAND2X0 r816_U261 ( .IN1(P1_N5111), .IN2(n7119), .QN(r816_n19) );
  INVX0 r816_U260 ( .ZN(r816_n151), .INP(r816_n19) );
  NOR2X0 r816_U258 ( .QN(r816_n30), .IN1(n7130), .IN2(P1_N5109) );
  AND2X1 r816_U257 ( .IN1(P1_N5109), .IN2(n7130), .Q(r816_n24) );
  NOR2X0 r816_U255 ( .QN(r816_n132), .IN1(n7144), .IN2(P1_N5107) );
  NAND2X0 r816_U254 ( .IN1(P1_N5107), .IN2(n7144), .QN(r816_n34) );
  INVX0 r816_U253 ( .ZN(r816_n166), .INP(r816_n34) );
  NOR2X0 r816_U251 ( .QN(r816_n45), .IN1(n7092), .IN2(P1_N5105) );
  AND2X1 r816_U250 ( .IN1(P1_N5105), .IN2(n7092), .Q(r816_n39) );
  NOR2X0 r816_U248 ( .QN(r816_n130), .IN1(n7098), .IN2(P1_N5103) );
  NAND2X0 r816_U247 ( .IN1(P1_N5103), .IN2(n7098), .QN(r816_n49) );
  INVX0 r816_U246 ( .ZN(r816_n181), .INP(r816_n49) );
  NOR2X0 r816_U244 ( .QN(r816_n60), .IN1(n7105), .IN2(P1_N5101) );
  AND2X1 r816_U243 ( .IN1(P1_N5101), .IN2(n7105), .Q(r816_n54) );
  NOR2X0 r816_U241 ( .QN(r816_n128), .IN1(n7112), .IN2(P1_N5099) );
  NAND2X0 r816_U240 ( .IN1(P1_N5099), .IN2(n7112), .QN(r816_n64) );
  INVX0 r816_U239 ( .ZN(r816_n196), .INP(r816_n64) );
  NOR2X0 r816_U237 ( .QN(r816_n75), .IN1(n7056), .IN2(P1_N5097) );
  AND2X1 r816_U236 ( .IN1(P1_N5097), .IN2(n7056), .Q(r816_n69) );
  NOR2X0 r816_U234 ( .QN(r816_n126), .IN1(n7063), .IN2(P1_N5095) );
  NAND2X0 r816_U233 ( .IN1(P1_N5095), .IN2(n7063), .QN(r816_n79) );
  INVX0 r816_U232 ( .ZN(r816_n211), .INP(r816_n79) );
  NOR2X0 r816_U230 ( .QN(r816_n90), .IN1(n7071), .IN2(P1_N5093) );
  AND2X1 r816_U229 ( .IN1(P1_N5093), .IN2(n7071), .Q(r816_n84) );
  NOR2X0 r816_U227 ( .QN(r816_n124), .IN1(n7076), .IN2(P1_N5091) );
  NAND2X0 r816_U226 ( .IN1(P1_N5091), .IN2(n7076), .QN(r816_n94) );
  INVX0 r816_U225 ( .ZN(r816_n226), .INP(r816_n94) );
  NOR2X0 r816_U223 ( .QN(r816_n105), .IN1(n7082), .IN2(P1_N5089) );
  AND2X1 r816_U222 ( .IN1(P1_N5089), .IN2(n7082), .Q(r816_n99) );
  NOR2X0 r816_U220 ( .QN(r816_n122), .IN1(n7043), .IN2(P1_N5087) );
  NAND2X0 r816_U219 ( .IN1(P1_N5087), .IN2(n7043), .QN(r816_n109) );
  INVX0 r816_U218 ( .ZN(r816_n241), .INP(r816_n109) );
  INVX0 r816_U216 ( .ZN(r816_n120), .INP(P1_N5084) );
  NOR2X0 r816_U215 ( .QN(r816_n250), .IN1(r816_n120), .IN2(n7034) );
  AND2X1 r816_U214 ( .IN1(n7051), .IN2(r816_n250), .Q(r816_n251) );
  NOR2X0 r816_U213 ( .QN(r816_n248), .IN1(P1_N5085), .IN2(r816_n251) );
  NOR2X0 r816_U212 ( .QN(r816_n249), .IN1(r816_n250), .IN2(n7051) );
  NOR2X0 r816_U211 ( .QN(r816_n245), .IN1(r816_n248), .IN2(r816_n249) );
  NOR2X0 r816_U209 ( .QN(r816_n121), .IN1(n7045), .IN2(P1_N5086) );
  NAND2X0 r816_U208 ( .IN1(P1_N5086), .IN2(n7045), .QN(r816_n244) );
  INVX0 r816_U207 ( .ZN(r816_n246), .INP(r816_n244) );
  NOR2X0 r816_U206 ( .QN(r816_n113), .IN1(r816_n121), .IN2(r816_n246) );
  NAND2X0 r816_U205 ( .IN1(r816_n245), .IN2(r816_n113), .QN(r816_n243) );
  NAND2X0 r816_U204 ( .IN1(r816_n243), .IN2(r816_n244), .QN(r816_n242) );
  NOR2X0 r816_U203 ( .QN(r816_n240), .IN1(r816_n241), .IN2(r816_n242) );
  NOR2X0 r816_U202 ( .QN(r816_n237), .IN1(r816_n122), .IN2(r816_n240) );
  OR2X1 r816_U200 ( .IN2(P1_N5088), .IN1(r816_n276), .Q(r816_n104) );
  NAND2X0 r816_U199 ( .IN1(P1_N5088), .IN2(r816_n276), .QN(r816_n236) );
  NAND2X0 r816_U198 ( .IN1(r816_n104), .IN2(r816_n236), .QN(r816_n106) );
  INVX0 r816_U197 ( .ZN(r816_n238), .INP(r816_n106) );
  NAND2X0 r816_U196 ( .IN1(r816_n237), .IN2(r816_n238), .QN(r816_n235) );
  NAND2X0 r816_U195 ( .IN1(r816_n235), .IN2(r816_n236), .QN(r816_n234) );
  NOR2X0 r816_U194 ( .QN(r816_n233), .IN1(r816_n99), .IN2(r816_n234) );
  NOR2X0 r816_U193 ( .QN(r816_n230), .IN1(r816_n105), .IN2(r816_n233) );
  NOR2X0 r816_U191 ( .QN(r816_n123), .IN1(n7079), .IN2(P1_N5090) );
  NAND2X0 r816_U190 ( .IN1(P1_N5090), .IN2(n7079), .QN(r816_n229) );
  INVX0 r816_U189 ( .ZN(r816_n231), .INP(r816_n229) );
  NOR2X0 r816_U188 ( .QN(r816_n98), .IN1(r816_n123), .IN2(r816_n231) );
  NAND2X0 r816_U187 ( .IN1(r816_n230), .IN2(r816_n98), .QN(r816_n228) );
  NAND2X0 r816_U186 ( .IN1(r816_n228), .IN2(r816_n229), .QN(r816_n227) );
  NOR2X0 r816_U185 ( .QN(r816_n225), .IN1(r816_n226), .IN2(r816_n227) );
  NOR2X0 r816_U184 ( .QN(r816_n222), .IN1(r816_n124), .IN2(r816_n225) );
  OR2X1 r816_U182 ( .IN2(P1_N5092), .IN1(n7073), .Q(r816_n89) );
  NAND2X0 r816_U181 ( .IN1(P1_N5092), .IN2(n7073), .QN(r816_n221) );
  NAND2X0 r816_U180 ( .IN1(r816_n89), .IN2(r816_n221), .QN(r816_n91) );
  INVX0 r816_U179 ( .ZN(r816_n223), .INP(r816_n91) );
  NAND2X0 r816_U178 ( .IN1(r816_n222), .IN2(r816_n223), .QN(r816_n220) );
  NAND2X0 r816_U177 ( .IN1(r816_n220), .IN2(r816_n221), .QN(r816_n219) );
  NOR2X0 r816_U176 ( .QN(r816_n218), .IN1(r816_n84), .IN2(r816_n219) );
  NOR2X0 r816_U175 ( .QN(r816_n215), .IN1(r816_n90), .IN2(r816_n218) );
  NOR2X0 r816_U173 ( .QN(r816_n125), .IN1(n7067), .IN2(P1_N5094) );
  OR2X1 r816_U267 ( .IN2(P1_N5115), .IN1(n4469), .Q(r816_n4) );
  INVX0 r816_U82 ( .ZN(r816_n276), .INP(n7036) );
  INVX0 r816_U84 ( .ZN(r816_n301), .INP(P1_N5175) );
  INVX0 r816_U93 ( .ZN(r816_n304), .INP(n7138) );
  INVX0 r816_U102 ( .ZN(r816_n308), .INP(P1_N5114) );
  NOR2X0 P1_sub_111_U53 ( .QN(P1_sub_111_n44), .IN1(n10187), .IN2(n10381) );
  NAND2X0 P1_sub_111_U52 ( .IN1(P1_sub_111_n44), .IN2(P1_sub_111_n45), 
        .QN(P1_sub_111_n38) );
  AND2X1 P1_sub_111_U51 ( .IN1(P1_sub_111_n38), .IN2(n10373), 
        .Q(P1_sub_111_n42) );
  NOR2X0 P1_sub_111_U50 ( .QN(P1_sub_111_n43), .IN1(n10373), 
        .IN2(P1_sub_111_n38) );
  NOR2X0 P1_sub_111_U49 ( .QN(P1_N129), .IN1(P1_sub_111_n42), 
        .IN2(P1_sub_111_n43) );
  OR2X1 P1_sub_111_U48 ( .IN2(n10373), .IN1(P1_sub_111_n38), 
        .Q(P1_sub_111_n41) );
  AND2X1 P1_sub_111_U47 ( .IN1(P1_sub_111_n41), .IN2(n10145), 
        .Q(P1_sub_111_n39) );
  NOR2X0 P1_sub_111_U46 ( .QN(P1_sub_111_n40), .IN1(n10145), 
        .IN2(P1_sub_111_n41) );
  NOR2X0 P1_sub_111_U45 ( .QN(P1_N130), .IN1(P1_sub_111_n39), 
        .IN2(P1_sub_111_n40) );
  NOR2X0 P1_sub_111_U44 ( .QN(P1_sub_111_n36), .IN1(n10145), .IN2(n10373) );
  INVX0 P1_sub_111_U43 ( .ZN(P1_sub_111_n37), .INP(P1_sub_111_n38) );
  NAND2X0 P1_sub_111_U42 ( .IN1(P1_sub_111_n36), .IN2(P1_sub_111_n37), 
        .QN(P1_sub_111_n30) );
  AND2X1 P1_sub_111_U41 ( .IN1(P1_sub_111_n30), .IN2(n10125), 
        .Q(P1_sub_111_n34) );
  NOR2X0 P1_sub_111_U40 ( .QN(P1_sub_111_n35), .IN1(n10125), 
        .IN2(P1_sub_111_n30) );
  NOR2X0 P1_sub_111_U39 ( .QN(P1_N131), .IN1(P1_sub_111_n34), 
        .IN2(P1_sub_111_n35) );
  OR2X1 P1_sub_111_U38 ( .IN2(n6624), .IN1(n6625), .Q(P1_sub_111_n33) );
  AND2X1 P1_sub_111_U37 ( .IN1(P1_sub_111_n33), .IN2(n6626), 
        .Q(P1_sub_111_n31) );
  NOR2X0 P1_sub_111_U36 ( .QN(P1_sub_111_n32), .IN1(n6626), 
        .IN2(P1_sub_111_n33) );
  NOR2X0 P1_sub_111_U35 ( .QN(P1_N104), .IN1(P1_sub_111_n31), 
        .IN2(P1_sub_111_n32) );
  OR2X1 P1_sub_111_U34 ( .IN2(n10125), .IN1(P1_sub_111_n30), 
        .Q(P1_sub_111_n27) );
  AND2X1 P1_sub_111_U33 ( .IN1(P1_sub_111_n27), .IN2(n10129), 
        .Q(P1_sub_111_n28) );
  NOR2X0 P1_sub_111_U32 ( .QN(P1_sub_111_n29), .IN1(n10129), 
        .IN2(P1_sub_111_n27) );
  NOR2X0 P1_sub_111_U31 ( .QN(P1_N132), .IN1(P1_sub_111_n28), 
        .IN2(P1_sub_111_n29) );
  OR2X1 P1_sub_111_U30 ( .IN2(n10129), .IN1(P1_sub_111_n27), 
        .Q(P1_sub_111_n26) );
  AND2X1 P1_sub_111_U29 ( .IN1(P1_sub_111_n26), .IN2(n6708), 
        .Q(P1_sub_111_n24) );
  NOR2X0 P1_sub_111_U28 ( .QN(P1_sub_111_n25), .IN1(n6708), 
        .IN2(P1_sub_111_n26) );
  NOR2X0 P1_sub_111_U27 ( .QN(P1_N133), .IN1(P1_sub_111_n24), 
        .IN2(P1_sub_111_n25) );
  AND2X1 P1_sub_111_U26 ( .IN1(P1_sub_111_n21), .IN2(n6627), 
        .Q(P1_sub_111_n22) );
  NOR2X0 P1_sub_111_U25 ( .QN(P1_sub_111_n23), .IN1(n6627), 
        .IN2(P1_sub_111_n21) );
  NOR2X0 P1_sub_111_U24 ( .QN(P1_N105), .IN1(P1_sub_111_n22), 
        .IN2(P1_sub_111_n23) );
  OR2X1 P1_sub_111_U23 ( .IN2(n6627), .IN1(P1_sub_111_n21), .Q(P1_sub_111_n20)
         );
  AND2X1 P1_sub_111_U22 ( .IN1(P1_sub_111_n20), .IN2(n6628), 
        .Q(P1_sub_111_n18) );
  NOR2X0 P1_sub_111_U21 ( .QN(P1_sub_111_n19), .IN1(n6628), 
        .IN2(P1_sub_111_n20) );
  NOR2X0 P1_sub_111_U20 ( .QN(P1_N106), .IN1(P1_sub_111_n18), 
        .IN2(P1_sub_111_n19) );
  INVX0 P1_sub_111_U19 ( .ZN(P1_sub_111_n14), .INP(P1_sub_111_n17) );
  AND2X1 P1_sub_111_U18 ( .IN1(P1_sub_111_n14), .IN2(n6629), 
        .Q(P1_sub_111_n15) );
  NOR2X0 P1_sub_111_U17 ( .QN(P1_sub_111_n16), .IN1(n6629), 
        .IN2(P1_sub_111_n14) );
  NOR2X0 P1_sub_111_U16 ( .QN(P1_N107), .IN1(P1_sub_111_n15), 
        .IN2(P1_sub_111_n16) );
  OR2X1 P1_sub_111_U15 ( .IN2(n6629), .IN1(P1_sub_111_n14), .Q(P1_sub_111_n13)
         );
  AND2X1 P1_sub_111_U14 ( .IN1(P1_sub_111_n13), .IN2(n6630), 
        .Q(P1_sub_111_n11) );
  NOR2X0 P1_sub_111_U13 ( .QN(P1_sub_111_n12), .IN1(n6630), 
        .IN2(P1_sub_111_n13) );
  NOR2X0 P1_sub_111_U12 ( .QN(P1_N108), .IN1(P1_sub_111_n11), 
        .IN2(P1_sub_111_n12) );
  AND2X1 P1_sub_111_U11 ( .IN1(P1_sub_111_n8), .IN2(n6631), .Q(P1_sub_111_n9)
         );
  NOR2X0 P1_sub_111_U10 ( .QN(P1_sub_111_n10), .IN1(n6631), 
        .IN2(P1_sub_111_n8) );
  NOR2X0 P1_sub_111_U9 ( .QN(P1_N109), .IN1(P1_sub_111_n9), 
        .IN2(P1_sub_111_n10) );
  OR2X1 P1_sub_111_U8 ( .IN2(n6631), .IN1(P1_sub_111_n8), .Q(P1_sub_111_n7) );
  AND2X1 P1_sub_111_U7 ( .IN1(P1_sub_111_n7), .IN2(n6632), .Q(P1_sub_111_n5)
         );
  NOR2X0 P1_sub_111_U6 ( .QN(P1_sub_111_n6), .IN1(n6632), .IN2(P1_sub_111_n7)
         );
  NOR2X0 P1_sub_111_U5 ( .QN(P1_N110), .IN1(P1_sub_111_n5), 
        .IN2(P1_sub_111_n6) );
  AND2X1 P1_sub_111_U4 ( .IN1(P1_sub_111_n4), .IN2(n6633), .Q(P1_sub_111_n2)
         );
  NOR2X0 P1_sub_111_U3 ( .QN(P1_sub_111_n3), .IN1(n6633), .IN2(P1_sub_111_n4)
         );
  NOR2X0 P1_sub_111_U2 ( .QN(P1_N111), .IN1(P1_sub_111_n2), 
        .IN2(P1_sub_111_n3) );
  OR2X1 P1_sub_111_U146 ( .IN2(n6631), .IN1(n6632), .Q(P1_sub_111_n112) );
  NOR2X0 P1_sub_111_U145 ( .QN(P1_sub_111_n113), .IN1(n6630), .IN2(n6629) );
  OR2X1 P1_sub_111_U144 ( .IN2(n6627), .IN1(n6628), .Q(P1_sub_111_n114) );
  NOR2X0 P1_sub_111_U143 ( .QN(P1_sub_111_n115), .IN1(n6626), .IN2(n6625) );
  NAND2X0 P1_sub_111_U141 ( .IN1(P1_sub_111_n115), .IN2(n18695), 
        .QN(P1_sub_111_n21) );
  NOR2X0 P1_sub_111_U140 ( .QN(P1_sub_111_n17), .IN1(P1_sub_111_n114), 
        .IN2(P1_sub_111_n21) );
  NAND2X0 P1_sub_111_U139 ( .IN1(P1_sub_111_n113), .IN2(P1_sub_111_n17), 
        .QN(P1_sub_111_n8) );
  NOR2X0 P1_sub_111_U138 ( .QN(P1_sub_111_n108), .IN1(P1_sub_111_n112), 
        .IN2(P1_sub_111_n8) );
  INVX0 P1_sub_111_U137 ( .ZN(P1_sub_111_n4), .INP(P1_sub_111_n108) );
  OR2X1 P1_sub_111_U136 ( .IN2(n6633), .IN1(P1_sub_111_n4), 
        .Q(P1_sub_111_n111) );
  AND2X1 P1_sub_111_U135 ( .IN1(P1_sub_111_n111), .IN2(n6634), 
        .Q(P1_sub_111_n109) );
  NOR2X0 P1_sub_111_U134 ( .QN(P1_sub_111_n110), .IN1(n6634), 
        .IN2(P1_sub_111_n111) );
  NOR2X0 P1_sub_111_U133 ( .QN(P1_N112), .IN1(P1_sub_111_n109), 
        .IN2(P1_sub_111_n110) );
  NOR2X0 P1_sub_111_U132 ( .QN(P1_sub_111_n107), .IN1(n6633), .IN2(n6634) );
  NAND2X0 P1_sub_111_U131 ( .IN1(P1_sub_111_n107), .IN2(P1_sub_111_n108), 
        .QN(P1_sub_111_n101) );
  AND2X1 P1_sub_111_U130 ( .IN1(P1_sub_111_n101), .IN2(n6635), 
        .Q(P1_sub_111_n105) );
  NOR2X0 P1_sub_111_U129 ( .QN(P1_sub_111_n106), .IN1(n6635), 
        .IN2(P1_sub_111_n101) );
  NOR2X0 P1_sub_111_U128 ( .QN(P1_N113), .IN1(P1_sub_111_n105), 
        .IN2(P1_sub_111_n106) );
  OR2X1 P1_sub_111_U127 ( .IN2(n6635), .IN1(P1_sub_111_n101), 
        .Q(P1_sub_111_n104) );
  AND2X1 P1_sub_111_U126 ( .IN1(P1_sub_111_n104), .IN2(n6636), 
        .Q(P1_sub_111_n102) );
  NOR2X0 P1_sub_111_U125 ( .QN(P1_sub_111_n103), .IN1(n6636), 
        .IN2(P1_sub_111_n104) );
  NOR2X0 P1_sub_111_U124 ( .QN(P1_N114), .IN1(P1_sub_111_n102), 
        .IN2(P1_sub_111_n103) );
  OR2X1 P1_sub_111_U123 ( .IN2(n6635), .IN1(n6636), .Q(P1_sub_111_n100) );
  NOR2X0 P1_sub_111_U122 ( .QN(P1_sub_111_n93), .IN1(P1_sub_111_n100), 
        .IN2(P1_sub_111_n101) );
  INVX0 P1_sub_111_U121 ( .ZN(P1_sub_111_n97), .INP(P1_sub_111_n93) );
  AND2X1 P1_sub_111_U120 ( .IN1(P1_sub_111_n97), .IN2(n6647), 
        .Q(P1_sub_111_n98) );
  NOR2X0 P1_sub_111_U119 ( .QN(P1_sub_111_n99), .IN1(n6647), 
        .IN2(P1_sub_111_n97) );
  NOR2X0 P1_sub_111_U118 ( .QN(P1_N115), .IN1(P1_sub_111_n98), 
        .IN2(P1_sub_111_n99) );
  OR2X1 P1_sub_111_U117 ( .IN2(n6647), .IN1(P1_sub_111_n97), 
        .Q(P1_sub_111_n96) );
  AND2X1 P1_sub_111_U116 ( .IN1(P1_sub_111_n96), .IN2(n6646), 
        .Q(P1_sub_111_n94) );
  NOR2X0 P1_sub_111_U115 ( .QN(P1_sub_111_n95), .IN1(n6646), 
        .IN2(P1_sub_111_n96) );
  NOR2X0 P1_sub_111_U114 ( .QN(P1_N116), .IN1(P1_sub_111_n94), 
        .IN2(P1_sub_111_n95) );
  NOR2X0 P1_sub_111_U113 ( .QN(P1_sub_111_n92), .IN1(n6646), .IN2(n6647) );
  NAND2X0 P1_sub_111_U112 ( .IN1(P1_sub_111_n92), .IN2(P1_sub_111_n93), 
        .QN(P1_sub_111_n86) );
  AND2X1 P1_sub_111_U111 ( .IN1(P1_sub_111_n86), .IN2(n6645), 
        .Q(P1_sub_111_n90) );
  NOR2X0 P1_sub_111_U110 ( .QN(P1_sub_111_n91), .IN1(n6645), 
        .IN2(P1_sub_111_n86) );
  NOR2X0 P1_sub_111_U109 ( .QN(P1_N117), .IN1(P1_sub_111_n90), 
        .IN2(P1_sub_111_n91) );
  OR2X1 P1_sub_111_U108 ( .IN2(n6645), .IN1(P1_sub_111_n86), 
        .Q(P1_sub_111_n89) );
  AND2X1 P1_sub_111_U107 ( .IN1(P1_sub_111_n89), .IN2(n6644), 
        .Q(P1_sub_111_n87) );
  NOR2X0 P1_sub_111_U106 ( .QN(P1_sub_111_n88), .IN1(n6644), 
        .IN2(P1_sub_111_n89) );
  NOR2X0 P1_sub_111_U105 ( .QN(P1_N118), .IN1(P1_sub_111_n87), 
        .IN2(P1_sub_111_n88) );
  OR2X1 P1_sub_111_U104 ( .IN2(n6645), .IN1(n6644), .Q(P1_sub_111_n85) );
  NOR2X0 P1_sub_111_U103 ( .QN(P1_sub_111_n78), .IN1(P1_sub_111_n85), 
        .IN2(P1_sub_111_n86) );
  INVX0 P1_sub_111_U102 ( .ZN(P1_sub_111_n82), .INP(P1_sub_111_n78) );
  AND2X1 P1_sub_111_U101 ( .IN1(P1_sub_111_n82), .IN2(n6643), 
        .Q(P1_sub_111_n83) );
  NOR2X0 P1_sub_111_U100 ( .QN(P1_sub_111_n84), .IN1(n6643), 
        .IN2(P1_sub_111_n82) );
  NOR2X0 P1_sub_111_U99 ( .QN(P1_N119), .IN1(P1_sub_111_n83), 
        .IN2(P1_sub_111_n84) );
  OR2X1 P1_sub_111_U98 ( .IN2(n6643), .IN1(P1_sub_111_n82), .Q(P1_sub_111_n81)
         );
  AND2X1 P1_sub_111_U97 ( .IN1(P1_sub_111_n81), .IN2(n6642), 
        .Q(P1_sub_111_n79) );
  NOR2X0 P1_sub_111_U96 ( .QN(P1_sub_111_n80), .IN1(n6642), 
        .IN2(P1_sub_111_n81) );
  NOR2X0 P1_sub_111_U95 ( .QN(P1_N120), .IN1(P1_sub_111_n79), 
        .IN2(P1_sub_111_n80) );
  NOR2X0 P1_sub_111_U94 ( .QN(P1_sub_111_n77), .IN1(n6642), .IN2(n6643) );
  NAND2X0 P1_sub_111_U93 ( .IN1(P1_sub_111_n77), .IN2(P1_sub_111_n78), 
        .QN(P1_sub_111_n68) );
  AND2X1 P1_sub_111_U92 ( .IN1(P1_sub_111_n68), .IN2(n6641), 
        .Q(P1_sub_111_n75) );
  NOR2X0 P1_sub_111_U91 ( .QN(P1_sub_111_n76), .IN1(n6641), 
        .IN2(P1_sub_111_n68) );
  NOR2X0 P1_sub_111_U90 ( .QN(P1_N121), .IN1(P1_sub_111_n75), 
        .IN2(P1_sub_111_n76) );
  OR2X1 P1_sub_111_U89 ( .IN2(n6625), .IN1(n18695), .Q(P1_sub_111_n72) );
  NAND2X0 P1_sub_111_U88 ( .IN1(n6625), .IN2(n18695), .QN(P1_sub_111_n73) );
  NAND2X0 P1_sub_111_U87 ( .IN1(P1_sub_111_n72), .IN2(P1_sub_111_n73), 
        .QN(P1_N103) );
  OR2X1 P1_sub_111_U86 ( .IN2(n6641), .IN1(P1_sub_111_n68), .Q(P1_sub_111_n71)
         );
  AND2X1 P1_sub_111_U85 ( .IN1(P1_sub_111_n71), .IN2(n6640), 
        .Q(P1_sub_111_n69) );
  NOR2X0 P1_sub_111_U84 ( .QN(P1_sub_111_n70), .IN1(n6640), 
        .IN2(P1_sub_111_n71) );
  NOR2X0 P1_sub_111_U83 ( .QN(P1_N122), .IN1(P1_sub_111_n69), 
        .IN2(P1_sub_111_n70) );
  OR2X1 P1_sub_111_U82 ( .IN2(n6641), .IN1(n6640), .Q(P1_sub_111_n67) );
  NOR2X0 P1_sub_111_U81 ( .QN(P1_sub_111_n60), .IN1(P1_sub_111_n67), 
        .IN2(P1_sub_111_n68) );
  INVX0 P1_sub_111_U80 ( .ZN(P1_sub_111_n64), .INP(P1_sub_111_n60) );
  AND2X1 P1_sub_111_U79 ( .IN1(P1_sub_111_n64), .IN2(n6639), 
        .Q(P1_sub_111_n65) );
  NOR2X0 P1_sub_111_U78 ( .QN(P1_sub_111_n66), .IN1(n6639), 
        .IN2(P1_sub_111_n64) );
  NOR2X0 P1_sub_111_U77 ( .QN(P1_N123), .IN1(P1_sub_111_n65), 
        .IN2(P1_sub_111_n66) );
  OR2X1 P1_sub_111_U76 ( .IN2(n6639), .IN1(P1_sub_111_n64), .Q(P1_sub_111_n63)
         );
  AND2X1 P1_sub_111_U75 ( .IN1(P1_sub_111_n63), .IN2(n6638), 
        .Q(P1_sub_111_n61) );
  NOR2X0 P1_sub_111_U74 ( .QN(P1_sub_111_n62), .IN1(n6638), 
        .IN2(P1_sub_111_n63) );
  NOR2X0 P1_sub_111_U73 ( .QN(P1_N124), .IN1(P1_sub_111_n61), 
        .IN2(P1_sub_111_n62) );
  NOR2X0 P1_sub_111_U72 ( .QN(P1_sub_111_n59), .IN1(n6638), .IN2(n6639) );
  NAND2X0 P1_sub_111_U71 ( .IN1(P1_sub_111_n59), .IN2(P1_sub_111_n60), 
        .QN(P1_sub_111_n53) );
  AND2X1 P1_sub_111_U70 ( .IN1(P1_sub_111_n53), .IN2(n6637), 
        .Q(P1_sub_111_n57) );
  NOR2X0 P1_sub_111_U69 ( .QN(P1_sub_111_n58), .IN1(n6637), 
        .IN2(P1_sub_111_n53) );
  NOR2X0 P1_sub_111_U68 ( .QN(P1_N125), .IN1(P1_sub_111_n57), 
        .IN2(P1_sub_111_n58) );
  OR2X1 P1_sub_111_U67 ( .IN2(n6637), .IN1(P1_sub_111_n53), .Q(P1_sub_111_n56)
         );
  AND2X1 P1_sub_111_U66 ( .IN1(P1_sub_111_n56), .IN2(n10195), 
        .Q(P1_sub_111_n54) );
  NOR2X0 P1_sub_111_U65 ( .QN(P1_sub_111_n55), .IN1(n10195), 
        .IN2(P1_sub_111_n56) );
  NOR2X0 P1_sub_111_U64 ( .QN(P1_N126), .IN1(P1_sub_111_n54), 
        .IN2(P1_sub_111_n55) );
  OR2X1 P1_sub_111_U63 ( .IN2(n6637), .IN1(n10195), .Q(P1_sub_111_n52) );
  NOR2X0 P1_sub_111_U62 ( .QN(P1_sub_111_n45), .IN1(P1_sub_111_n52), 
        .IN2(P1_sub_111_n53) );
  INVX0 P1_sub_111_U61 ( .ZN(P1_sub_111_n49), .INP(P1_sub_111_n45) );
  AND2X1 P1_sub_111_U60 ( .IN1(P1_sub_111_n49), .IN2(n10381), 
        .Q(P1_sub_111_n50) );
  NOR2X0 P1_sub_111_U59 ( .QN(P1_sub_111_n51), .IN1(n10381), 
        .IN2(P1_sub_111_n49) );
  NOR2X0 P1_sub_111_U58 ( .QN(P1_N127), .IN1(P1_sub_111_n50), 
        .IN2(P1_sub_111_n51) );
  OR2X1 P1_sub_111_U57 ( .IN2(n10381), .IN1(P1_sub_111_n49), 
        .Q(P1_sub_111_n48) );
  AND2X1 P1_sub_111_U56 ( .IN1(P1_sub_111_n48), .IN2(n10187), 
        .Q(P1_sub_111_n46) );
  NOR2X0 P1_sub_111_U55 ( .QN(P1_sub_111_n47), .IN1(n10187), 
        .IN2(P1_sub_111_n48) );
  NOR2X0 P1_sub_111_U54 ( .QN(P1_N128), .IN1(P1_sub_111_n46), 
        .IN2(P1_sub_111_n47) );
  NAND2X0 r792_U77 ( .IN1(r792_n78), .IN2(r792_n79), .QN(r792_n77) );
  NOR2X0 r792_U76 ( .QN(r792_n75), .IN1(r792_n71), .IN2(r792_n77) );
  AND2X1 r792_U75 ( .IN1(r792_n71), .IN2(r792_n77), .Q(r792_n76) );
  NOR2X0 r792_U74 ( .QN(n193), .IN1(r792_n75), .IN2(r792_n76) );
  INVX0 r792_U73 ( .ZN(r792_n74), .INP(P1_N344) );
  OR2X1 r792_U72 ( .IN2(n9493), .IN1(r792_n74), .Q(r792_n72) );
  NAND2X0 r792_U71 ( .IN1(n9493), .IN2(r792_n74), .QN(r792_n73) );
  NAND2X0 r792_U70 ( .IN1(r792_n72), .IN2(r792_n73), .QN(r792_n67) );
  NAND2X0 r792_U69 ( .IN1(P1_N345), .IN2(r792_n71), .QN(r792_n68) );
  OR2X1 r792_U68 ( .IN2(P1_N345), .IN1(r792_n71), .Q(r792_n70) );
  NAND2X0 r792_U67 ( .IN1(n9693), .IN2(r792_n70), .QN(r792_n69) );
  NAND2X0 r792_U66 ( .IN1(r792_n68), .IN2(r792_n69), .QN(r792_n66) );
  NOR2X0 r792_U65 ( .QN(r792_n64), .IN1(r792_n67), .IN2(r792_n66) );
  AND2X1 r792_U64 ( .IN1(r792_n66), .IN2(r792_n67), .Q(r792_n65) );
  NOR2X0 r792_U63 ( .QN(n192), .IN1(r792_n64), .IN2(r792_n65) );
  OR2X1 r792_U62 ( .IN2(n9761), .IN1(n6732), .Q(r792_n61) );
  NAND2X0 r792_U61 ( .IN1(n9761), .IN2(n6732), .QN(r792_n62) );
  NAND2X0 r792_U60 ( .IN1(r792_n61), .IN2(r792_n62), .QN(r792_n59) );
  NAND2X0 r792_U59 ( .IN1(r792_n59), .IN2(r792_n60), .QN(r792_n57) );
  OR2X1 r792_U58 ( .IN2(r792_n60), .IN1(r792_n59), .Q(r792_n58) );
  NAND2X0 r792_U57 ( .IN1(r792_n57), .IN2(r792_n58), .QN(n210) );
  OR2X1 r792_U55 ( .IN2(n9757), .IN1(n6734), .Q(r792_n54) );
  NAND2X0 r792_U54 ( .IN1(n9757), .IN2(n6734), .QN(r792_n55) );
  NAND2X0 r792_U53 ( .IN1(r792_n54), .IN2(r792_n55), .QN(r792_n53) );
  NOR2X0 r792_U52 ( .QN(r792_n50), .IN1(r792_n52), .IN2(r792_n53) );
  AND2X1 r792_U51 ( .IN1(r792_n52), .IN2(r792_n53), .Q(r792_n51) );
  NOR2X0 r792_U50 ( .QN(n209), .IN1(r792_n50), .IN2(r792_n51) );
  OR2X1 r792_U48 ( .IN2(n9753), .IN1(n6742), .Q(r792_n47) );
  NAND2X0 r792_U47 ( .IN1(n9753), .IN2(n6742), .QN(r792_n48) );
  NAND2X0 r792_U46 ( .IN1(r792_n47), .IN2(r792_n48), .QN(r792_n46) );
  NOR2X0 r792_U45 ( .QN(r792_n43), .IN1(r792_n45), .IN2(r792_n46) );
  AND2X1 r792_U44 ( .IN1(r792_n45), .IN2(r792_n46), .Q(r792_n44) );
  NOR2X0 r792_U43 ( .QN(n208), .IN1(r792_n43), .IN2(r792_n44) );
  OR2X1 r792_U41 ( .IN2(n9749), .IN1(n6744), .Q(r792_n40) );
  NAND2X0 r792_U40 ( .IN1(n9749), .IN2(n6744), .QN(r792_n41) );
  NAND2X0 r792_U39 ( .IN1(r792_n40), .IN2(r792_n41), .QN(r792_n39) );
  NOR2X0 r792_U38 ( .QN(r792_n36), .IN1(r792_n38), .IN2(r792_n39) );
  AND2X1 r792_U37 ( .IN1(r792_n38), .IN2(r792_n39), .Q(r792_n37) );
  NOR2X0 r792_U36 ( .QN(n207), .IN1(r792_n36), .IN2(r792_n37) );
  OR2X1 r792_U34 ( .IN2(n9745), .IN1(n6747), .Q(r792_n33) );
  NAND2X0 r792_U33 ( .IN1(n9745), .IN2(n6747), .QN(r792_n34) );
  NAND2X0 r792_U32 ( .IN1(r792_n33), .IN2(r792_n34), .QN(r792_n32) );
  NOR2X0 r792_U31 ( .QN(r792_n29), .IN1(r792_n31), .IN2(r792_n32) );
  AND2X1 r792_U30 ( .IN1(r792_n31), .IN2(r792_n32), .Q(r792_n30) );
  NOR2X0 r792_U29 ( .QN(n206), .IN1(r792_n29), .IN2(r792_n30) );
  OR2X1 r792_U27 ( .IN2(n9741), .IN1(n6751), .Q(r792_n26) );
  NAND2X0 r792_U26 ( .IN1(n9741), .IN2(n6751), .QN(r792_n27) );
  NAND2X0 r792_U25 ( .IN1(r792_n26), .IN2(r792_n27), .QN(r792_n25) );
  NOR2X0 r792_U24 ( .QN(r792_n22), .IN1(r792_n24), .IN2(r792_n25) );
  AND2X1 r792_U23 ( .IN1(r792_n24), .IN2(r792_n25), .Q(r792_n23) );
  NOR2X0 r792_U22 ( .QN(n205), .IN1(r792_n22), .IN2(r792_n23) );
  OR2X1 r792_U20 ( .IN2(n9737), .IN1(n6746), .Q(r792_n19) );
  NAND2X0 r792_U19 ( .IN1(n9737), .IN2(n6746), .QN(r792_n20) );
  NAND2X0 r792_U18 ( .IN1(r792_n19), .IN2(r792_n20), .QN(r792_n18) );
  NOR2X0 r792_U17 ( .QN(r792_n15), .IN1(r792_n17), .IN2(r792_n18) );
  AND2X1 r792_U16 ( .IN1(r792_n17), .IN2(r792_n18), .Q(r792_n16) );
  NOR2X0 r792_U15 ( .QN(n204), .IN1(r792_n15), .IN2(r792_n16) );
  OR2X1 r792_U13 ( .IN2(n9733), .IN1(n6750), .Q(r792_n12) );
  NAND2X0 r792_U12 ( .IN1(n9733), .IN2(n6750), .QN(r792_n13) );
  NAND2X0 r792_U11 ( .IN1(r792_n12), .IN2(r792_n13), .QN(r792_n11) );
  NOR2X0 r792_U10 ( .QN(r792_n8), .IN1(r792_n10), .IN2(r792_n11) );
  AND2X1 r792_U9 ( .IN1(r792_n10), .IN2(r792_n11), .Q(r792_n9) );
  NOR2X0 r792_U8 ( .QN(n203), .IN1(r792_n8), .IN2(r792_n9) );
  OR2X1 r792_U6 ( .IN2(n9729), .IN1(n6755), .Q(r792_n5) );
  NAND2X0 r792_U5 ( .IN1(n9729), .IN2(n6755), .QN(r792_n6) );
  NAND2X0 r792_U4 ( .IN1(r792_n5), .IN2(r792_n6), .QN(r792_n4) );
  NOR2X0 r792_U3 ( .QN(r792_n1), .IN1(r792_n3), .IN2(r792_n4) );
  AND2X1 r792_U2 ( .IN1(r792_n3), .IN2(r792_n4), .Q(r792_n2) );
  NOR2X0 r792_U1 ( .QN(n202), .IN1(r792_n1), .IN2(r792_n2) );
  NAND2X0 r792_U170 ( .IN1(n9729), .IN2(r792_n163), .QN(r792_n162) );
  NAND2X0 r792_U169 ( .IN1(r792_n161), .IN2(r792_n162), .QN(r792_n154) );
  OR2X1 r792_U167 ( .IN2(n9725), .IN1(n6759), .Q(r792_n158) );
  NAND2X0 r792_U166 ( .IN1(n9725), .IN2(n6759), .QN(r792_n159) );
  NAND2X0 r792_U165 ( .IN1(r792_n158), .IN2(r792_n159), .QN(r792_n157) );
  NOR2X0 r792_U164 ( .QN(r792_n155), .IN1(r792_n154), .IN2(r792_n157) );
  AND2X1 r792_U163 ( .IN1(r792_n154), .IN2(r792_n157), .Q(r792_n156) );
  NOR2X0 r792_U162 ( .QN(n201), .IN1(r792_n155), .IN2(r792_n156) );
  NAND2X0 r792_U161 ( .IN1(P1_N353), .IN2(r792_n154), .QN(r792_n151) );
  OR2X1 r792_U160 ( .IN2(P1_N353), .IN1(r792_n154), .Q(r792_n153) );
  NAND2X0 r792_U159 ( .IN1(n9725), .IN2(r792_n153), .QN(r792_n152) );
  NAND2X0 r792_U158 ( .IN1(r792_n151), .IN2(r792_n152), .QN(r792_n144) );
  OR2X1 r792_U156 ( .IN2(n9721), .IN1(n6754), .Q(r792_n148) );
  NAND2X0 r792_U155 ( .IN1(n9721), .IN2(n6754), .QN(r792_n149) );
  NAND2X0 r792_U154 ( .IN1(r792_n148), .IN2(r792_n149), .QN(r792_n147) );
  NOR2X0 r792_U153 ( .QN(r792_n145), .IN1(r792_n144), .IN2(r792_n147) );
  AND2X1 r792_U152 ( .IN1(r792_n144), .IN2(r792_n147), .Q(r792_n146) );
  NOR2X0 r792_U151 ( .QN(n200), .IN1(r792_n145), .IN2(r792_n146) );
  NAND2X0 r792_U150 ( .IN1(P1_N352), .IN2(r792_n144), .QN(r792_n141) );
  OR2X1 r792_U149 ( .IN2(P1_N352), .IN1(r792_n144), .Q(r792_n143) );
  NAND2X0 r792_U148 ( .IN1(n9721), .IN2(r792_n143), .QN(r792_n142) );
  NAND2X0 r792_U147 ( .IN1(r792_n141), .IN2(r792_n142), .QN(r792_n134) );
  OR2X1 r792_U145 ( .IN2(n9717), .IN1(n6758), .Q(r792_n138) );
  NAND2X0 r792_U144 ( .IN1(n9717), .IN2(n6758), .QN(r792_n139) );
  NAND2X0 r792_U143 ( .IN1(r792_n138), .IN2(r792_n139), .QN(r792_n137) );
  NOR2X0 r792_U142 ( .QN(r792_n135), .IN1(r792_n134), .IN2(r792_n137) );
  AND2X1 r792_U141 ( .IN1(r792_n134), .IN2(r792_n137), .Q(r792_n136) );
  NOR2X0 r792_U140 ( .QN(n199), .IN1(r792_n135), .IN2(r792_n136) );
  NAND2X0 r792_U139 ( .IN1(P1_N351), .IN2(r792_n134), .QN(r792_n131) );
  OR2X1 r792_U138 ( .IN2(P1_N351), .IN1(r792_n134), .Q(r792_n133) );
  NAND2X0 r792_U137 ( .IN1(n9717), .IN2(r792_n133), .QN(r792_n132) );
  NAND2X0 r792_U136 ( .IN1(r792_n131), .IN2(r792_n132), .QN(r792_n124) );
  OR2X1 r792_U134 ( .IN2(n9713), .IN1(n6763), .Q(r792_n128) );
  NAND2X0 r792_U133 ( .IN1(n9713), .IN2(n6763), .QN(r792_n129) );
  NAND2X0 r792_U132 ( .IN1(r792_n128), .IN2(r792_n129), .QN(r792_n127) );
  NOR2X0 r792_U131 ( .QN(r792_n125), .IN1(r792_n124), .IN2(r792_n127) );
  AND2X1 r792_U130 ( .IN1(r792_n124), .IN2(r792_n127), .Q(r792_n126) );
  NOR2X0 r792_U129 ( .QN(n198), .IN1(r792_n125), .IN2(r792_n126) );
  NAND2X0 r792_U128 ( .IN1(P1_N350), .IN2(r792_n124), .QN(r792_n121) );
  OR2X1 r792_U127 ( .IN2(P1_N350), .IN1(r792_n124), .Q(r792_n123) );
  NAND2X0 r792_U126 ( .IN1(n9713), .IN2(r792_n123), .QN(r792_n122) );
  NAND2X0 r792_U125 ( .IN1(r792_n121), .IN2(r792_n122), .QN(r792_n114) );
  OR2X1 r792_U123 ( .IN2(n9709), .IN1(n6767), .Q(r792_n118) );
  NAND2X0 r792_U122 ( .IN1(n9709), .IN2(n6767), .QN(r792_n119) );
  NAND2X0 r792_U121 ( .IN1(r792_n118), .IN2(r792_n119), .QN(r792_n117) );
  NOR2X0 r792_U120 ( .QN(r792_n115), .IN1(r792_n114), .IN2(r792_n117) );
  AND2X1 r792_U119 ( .IN1(r792_n114), .IN2(r792_n117), .Q(r792_n116) );
  NOR2X0 r792_U118 ( .QN(n197), .IN1(r792_n115), .IN2(r792_n116) );
  NAND2X0 r792_U117 ( .IN1(P1_N349), .IN2(r792_n114), .QN(r792_n111) );
  OR2X1 r792_U116 ( .IN2(P1_N349), .IN1(r792_n114), .Q(r792_n113) );
  NAND2X0 r792_U115 ( .IN1(n9709), .IN2(r792_n113), .QN(r792_n112) );
  NAND2X0 r792_U114 ( .IN1(r792_n111), .IN2(r792_n112), .QN(r792_n104) );
  OR2X1 r792_U112 ( .IN2(n9705), .IN1(n6762), .Q(r792_n108) );
  NAND2X0 r792_U111 ( .IN1(n9705), .IN2(n6762), .QN(r792_n109) );
  NAND2X0 r792_U110 ( .IN1(r792_n108), .IN2(r792_n109), .QN(r792_n107) );
  NOR2X0 r792_U109 ( .QN(r792_n105), .IN1(r792_n104), .IN2(r792_n107) );
  AND2X1 r792_U108 ( .IN1(r792_n104), .IN2(r792_n107), .Q(r792_n106) );
  NOR2X0 r792_U107 ( .QN(n196), .IN1(r792_n105), .IN2(r792_n106) );
  NAND2X0 r792_U106 ( .IN1(P1_N348), .IN2(r792_n104), .QN(r792_n101) );
  OR2X1 r792_U105 ( .IN2(P1_N348), .IN1(r792_n104), .Q(r792_n103) );
  NAND2X0 r792_U104 ( .IN1(n9705), .IN2(r792_n103), .QN(r792_n102) );
  NAND2X0 r792_U103 ( .IN1(r792_n101), .IN2(r792_n102), .QN(r792_n94) );
  OR2X1 r792_U101 ( .IN2(n9701), .IN1(n6766), .Q(r792_n98) );
  NAND2X0 r792_U100 ( .IN1(n9701), .IN2(n6766), .QN(r792_n99) );
  NAND2X0 r792_U99 ( .IN1(r792_n98), .IN2(r792_n99), .QN(r792_n97) );
  NOR2X0 r792_U98 ( .QN(r792_n95), .IN1(r792_n94), .IN2(r792_n97) );
  AND2X1 r792_U97 ( .IN1(r792_n94), .IN2(r792_n97), .Q(r792_n96) );
  NOR2X0 r792_U96 ( .QN(n195), .IN1(r792_n95), .IN2(r792_n96) );
  NAND2X0 r792_U95 ( .IN1(P1_N347), .IN2(r792_n94), .QN(r792_n91) );
  OR2X1 r792_U94 ( .IN2(P1_N347), .IN1(r792_n94), .Q(r792_n93) );
  NAND2X0 r792_U93 ( .IN1(n9701), .IN2(r792_n93), .QN(r792_n92) );
  NAND2X0 r792_U92 ( .IN1(r792_n91), .IN2(r792_n92), .QN(r792_n84) );
  OR2X1 r792_U90 ( .IN2(n9697), .IN1(n6770), .Q(r792_n88) );
  NAND2X0 r792_U89 ( .IN1(n9697), .IN2(n6770), .QN(r792_n89) );
  NAND2X0 r792_U88 ( .IN1(r792_n88), .IN2(r792_n89), .QN(r792_n87) );
  NOR2X0 r792_U87 ( .QN(r792_n85), .IN1(r792_n84), .IN2(r792_n87) );
  AND2X1 r792_U86 ( .IN1(r792_n84), .IN2(r792_n87), .Q(r792_n86) );
  NOR2X0 r792_U85 ( .QN(n194), .IN1(r792_n85), .IN2(r792_n86) );
  NAND2X0 r792_U84 ( .IN1(P1_N346), .IN2(r792_n84), .QN(r792_n81) );
  OR2X1 r792_U83 ( .IN2(P1_N346), .IN1(r792_n84), .Q(r792_n83) );
  NAND2X0 r792_U82 ( .IN1(n9697), .IN2(r792_n83), .QN(r792_n82) );
  NAND2X0 r792_U81 ( .IN1(r792_n81), .IN2(r792_n82), .QN(r792_n71) );
  OR2X1 r792_U79 ( .IN2(n9693), .IN1(n6773), .Q(r792_n78) );
  NAND2X0 r792_U78 ( .IN1(n9693), .IN2(n6773), .QN(r792_n79) );
  OR2X1 r792_U209 ( .IN2(n981), .IN1(n6730), .Q(r792_n188) );
  NAND2X0 r792_U208 ( .IN1(n981), .IN2(n6730), .QN(r792_n189) );
  NAND2X0 r792_U207 ( .IN1(r792_n188), .IN2(r792_n189), .QN(n211) );
  NAND2X0 r792_U205 ( .IN1(n981), .IN2(P1_N363), .QN(r792_n60) );
  OR2X1 r792_U204 ( .IN2(r792_n60), .IN1(n6732), .Q(r792_n185) );
  NAND2X0 r792_U203 ( .IN1(n6732), .IN2(r792_n60), .QN(r792_n187) );
  NAND2X0 r792_U202 ( .IN1(n9761), .IN2(r792_n187), .QN(r792_n186) );
  NAND2X0 r792_U201 ( .IN1(r792_n185), .IN2(r792_n186), .QN(r792_n52) );
  NAND2X0 r792_U200 ( .IN1(P1_N361), .IN2(r792_n52), .QN(r792_n182) );
  OR2X1 r792_U199 ( .IN2(P1_N361), .IN1(r792_n52), .Q(r792_n184) );
  NAND2X0 r792_U198 ( .IN1(n9757), .IN2(r792_n184), .QN(r792_n183) );
  NAND2X0 r792_U197 ( .IN1(r792_n182), .IN2(r792_n183), .QN(r792_n45) );
  NAND2X0 r792_U196 ( .IN1(P1_N360), .IN2(r792_n45), .QN(r792_n179) );
  OR2X1 r792_U195 ( .IN2(P1_N360), .IN1(r792_n45), .Q(r792_n181) );
  NAND2X0 r792_U194 ( .IN1(n9753), .IN2(r792_n181), .QN(r792_n180) );
  NAND2X0 r792_U193 ( .IN1(r792_n179), .IN2(r792_n180), .QN(r792_n38) );
  NAND2X0 r792_U192 ( .IN1(P1_N359), .IN2(r792_n38), .QN(r792_n176) );
  OR2X1 r792_U191 ( .IN2(P1_N359), .IN1(r792_n38), .Q(r792_n178) );
  NAND2X0 r792_U190 ( .IN1(n9749), .IN2(r792_n178), .QN(r792_n177) );
  NAND2X0 r792_U189 ( .IN1(r792_n176), .IN2(r792_n177), .QN(r792_n31) );
  NAND2X0 r792_U188 ( .IN1(P1_N358), .IN2(r792_n31), .QN(r792_n173) );
  OR2X1 r792_U187 ( .IN2(P1_N358), .IN1(r792_n31), .Q(r792_n175) );
  NAND2X0 r792_U186 ( .IN1(n9745), .IN2(r792_n175), .QN(r792_n174) );
  NAND2X0 r792_U185 ( .IN1(r792_n173), .IN2(r792_n174), .QN(r792_n24) );
  NAND2X0 r792_U184 ( .IN1(P1_N357), .IN2(r792_n24), .QN(r792_n170) );
  OR2X1 r792_U183 ( .IN2(P1_N357), .IN1(r792_n24), .Q(r792_n172) );
  NAND2X0 r792_U182 ( .IN1(n9741), .IN2(r792_n172), .QN(r792_n171) );
  NAND2X0 r792_U181 ( .IN1(r792_n170), .IN2(r792_n171), .QN(r792_n17) );
  NAND2X0 r792_U180 ( .IN1(P1_N356), .IN2(r792_n17), .QN(r792_n167) );
  OR2X1 r792_U179 ( .IN2(P1_N356), .IN1(r792_n17), .Q(r792_n169) );
  NAND2X0 r792_U178 ( .IN1(n9737), .IN2(r792_n169), .QN(r792_n168) );
  NAND2X0 r792_U177 ( .IN1(r792_n167), .IN2(r792_n168), .QN(r792_n10) );
  NAND2X0 r792_U176 ( .IN1(P1_N355), .IN2(r792_n10), .QN(r792_n164) );
  OR2X1 r792_U175 ( .IN2(P1_N355), .IN1(r792_n10), .Q(r792_n166) );
  NAND2X0 r792_U174 ( .IN1(n9733), .IN2(r792_n166), .QN(r792_n165) );
  NAND2X0 r792_U173 ( .IN1(r792_n164), .IN2(r792_n165), .QN(r792_n3) );
  NAND2X0 r792_U172 ( .IN1(P1_N354), .IN2(r792_n3), .QN(r792_n161) );
  OR2X1 r792_U171 ( .IN2(P1_N354), .IN1(r792_n3), .Q(r792_n163) );
  NOR2X0 r793_U8 ( .QN(n182), .IN1(r793_n8), .IN2(r793_n9) );
  OR2X1 r793_U6 ( .IN2(n9801), .IN1(n6755), .Q(r793_n5) );
  NAND2X0 r793_U5 ( .IN1(n9801), .IN2(n6755), .QN(r793_n6) );
  NAND2X0 r793_U4 ( .IN1(r793_n5), .IN2(r793_n6), .QN(r793_n4) );
  NOR2X0 r793_U3 ( .QN(r793_n1), .IN1(r793_n3), .IN2(r793_n4) );
  AND2X1 r793_U2 ( .IN1(r793_n3), .IN2(r793_n4), .Q(r793_n2) );
  NOR2X0 r793_U1 ( .QN(n181), .IN1(r793_n1), .IN2(r793_n2) );
  OR2X1 r793_U101 ( .IN2(n9773), .IN1(n6766), .Q(r793_n98) );
  NAND2X0 r793_U100 ( .IN1(n9773), .IN2(n6766), .QN(r793_n99) );
  NAND2X0 r793_U99 ( .IN1(r793_n98), .IN2(r793_n99), .QN(r793_n97) );
  NOR2X0 r793_U98 ( .QN(r793_n95), .IN1(r793_n94), .IN2(r793_n97) );
  AND2X1 r793_U97 ( .IN1(r793_n94), .IN2(r793_n97), .Q(r793_n96) );
  NOR2X0 r793_U96 ( .QN(n174), .IN1(r793_n95), .IN2(r793_n96) );
  NAND2X0 r793_U95 ( .IN1(P1_N347), .IN2(r793_n94), .QN(r793_n91) );
  OR2X1 r793_U94 ( .IN2(P1_N347), .IN1(r793_n94), .Q(r793_n93) );
  NAND2X0 r793_U93 ( .IN1(n9773), .IN2(r793_n93), .QN(r793_n92) );
  NAND2X0 r793_U92 ( .IN1(r793_n91), .IN2(r793_n92), .QN(r793_n84) );
  OR2X1 r793_U90 ( .IN2(n9769), .IN1(n6770), .Q(r793_n88) );
  NAND2X0 r793_U89 ( .IN1(n9769), .IN2(n6770), .QN(r793_n89) );
  NAND2X0 r793_U88 ( .IN1(r793_n88), .IN2(r793_n89), .QN(r793_n87) );
  NOR2X0 r793_U87 ( .QN(r793_n85), .IN1(r793_n84), .IN2(r793_n87) );
  AND2X1 r793_U86 ( .IN1(r793_n84), .IN2(r793_n87), .Q(r793_n86) );
  NOR2X0 r793_U85 ( .QN(n173), .IN1(r793_n85), .IN2(r793_n86) );
  NAND2X0 r793_U84 ( .IN1(P1_N346), .IN2(r793_n84), .QN(r793_n81) );
  OR2X1 r793_U83 ( .IN2(P1_N346), .IN1(r793_n84), .Q(r793_n83) );
  NAND2X0 r793_U82 ( .IN1(n9769), .IN2(r793_n83), .QN(r793_n82) );
  NAND2X0 r793_U81 ( .IN1(r793_n81), .IN2(r793_n82), .QN(r793_n71) );
  OR2X1 r793_U79 ( .IN2(n9765), .IN1(n6773), .Q(r793_n78) );
  NAND2X0 r793_U78 ( .IN1(n9765), .IN2(n6773), .QN(r793_n79) );
  NAND2X0 r793_U77 ( .IN1(r793_n78), .IN2(r793_n79), .QN(r793_n77) );
  NOR2X0 r793_U76 ( .QN(r793_n75), .IN1(r793_n71), .IN2(r793_n77) );
  AND2X1 r793_U75 ( .IN1(r793_n71), .IN2(r793_n77), .Q(r793_n76) );
  NOR2X0 r793_U74 ( .QN(n172), .IN1(r793_n75), .IN2(r793_n76) );
  INVX0 r793_U73 ( .ZN(r793_n74), .INP(P1_N344) );
  OR2X1 r793_U72 ( .IN2(n9497), .IN1(r793_n74), .Q(r793_n72) );
  NAND2X0 r793_U71 ( .IN1(n9497), .IN2(r793_n74), .QN(r793_n73) );
  NAND2X0 r793_U70 ( .IN1(r793_n72), .IN2(r793_n73), .QN(r793_n67) );
  NAND2X0 r793_U69 ( .IN1(P1_N345), .IN2(r793_n71), .QN(r793_n68) );
  OR2X1 r793_U68 ( .IN2(P1_N345), .IN1(r793_n71), .Q(r793_n70) );
  NAND2X0 r793_U67 ( .IN1(n9765), .IN2(r793_n70), .QN(r793_n69) );
  NAND2X0 r793_U66 ( .IN1(r793_n68), .IN2(r793_n69), .QN(r793_n66) );
  NOR2X0 r793_U65 ( .QN(r793_n64), .IN1(r793_n67), .IN2(r793_n66) );
  AND2X1 r793_U64 ( .IN1(r793_n66), .IN2(r793_n67), .Q(r793_n65) );
  NOR2X0 r793_U63 ( .QN(n171), .IN1(r793_n64), .IN2(r793_n65) );
  OR2X1 r793_U62 ( .IN2(n9833), .IN1(n6732), .Q(r793_n61) );
  NAND2X0 r793_U61 ( .IN1(n9833), .IN2(n6732), .QN(r793_n62) );
  NAND2X0 r793_U60 ( .IN1(r793_n61), .IN2(r793_n62), .QN(r793_n59) );
  NAND2X0 r793_U59 ( .IN1(r793_n59), .IN2(r793_n60), .QN(r793_n57) );
  OR2X1 r793_U58 ( .IN2(r793_n60), .IN1(r793_n59), .Q(r793_n58) );
  NAND2X0 r793_U57 ( .IN1(r793_n57), .IN2(r793_n58), .QN(n189) );
  OR2X1 r793_U55 ( .IN2(n9829), .IN1(n6734), .Q(r793_n54) );
  NAND2X0 r793_U54 ( .IN1(n9829), .IN2(n6734), .QN(r793_n55) );
  NAND2X0 r793_U53 ( .IN1(r793_n54), .IN2(r793_n55), .QN(r793_n53) );
  NOR2X0 r793_U52 ( .QN(r793_n50), .IN1(r793_n52), .IN2(r793_n53) );
  AND2X1 r793_U51 ( .IN1(r793_n52), .IN2(r793_n53), .Q(r793_n51) );
  NOR2X0 r793_U50 ( .QN(n188), .IN1(r793_n50), .IN2(r793_n51) );
  OR2X1 r793_U48 ( .IN2(n9825), .IN1(n6742), .Q(r793_n47) );
  NAND2X0 r793_U47 ( .IN1(n9825), .IN2(n6742), .QN(r793_n48) );
  NAND2X0 r793_U46 ( .IN1(r793_n47), .IN2(r793_n48), .QN(r793_n46) );
  NOR2X0 r793_U45 ( .QN(r793_n43), .IN1(r793_n45), .IN2(r793_n46) );
  AND2X1 r793_U44 ( .IN1(r793_n45), .IN2(r793_n46), .Q(r793_n44) );
  NOR2X0 r793_U43 ( .QN(n187), .IN1(r793_n43), .IN2(r793_n44) );
  OR2X1 r793_U41 ( .IN2(n9821), .IN1(n6744), .Q(r793_n40) );
  NAND2X0 r793_U40 ( .IN1(n9821), .IN2(n6744), .QN(r793_n41) );
  NAND2X0 r793_U39 ( .IN1(r793_n40), .IN2(r793_n41), .QN(r793_n39) );
  NOR2X0 r793_U38 ( .QN(r793_n36), .IN1(r793_n38), .IN2(r793_n39) );
  AND2X1 r793_U37 ( .IN1(r793_n38), .IN2(r793_n39), .Q(r793_n37) );
  NOR2X0 r793_U36 ( .QN(n186), .IN1(r793_n36), .IN2(r793_n37) );
  OR2X1 r793_U34 ( .IN2(n9817), .IN1(n6747), .Q(r793_n33) );
  NAND2X0 r793_U33 ( .IN1(n9817), .IN2(n6747), .QN(r793_n34) );
  NAND2X0 r793_U32 ( .IN1(r793_n33), .IN2(r793_n34), .QN(r793_n32) );
  NOR2X0 r793_U31 ( .QN(r793_n29), .IN1(r793_n31), .IN2(r793_n32) );
  AND2X1 r793_U30 ( .IN1(r793_n31), .IN2(r793_n32), .Q(r793_n30) );
  NOR2X0 r793_U29 ( .QN(n185), .IN1(r793_n29), .IN2(r793_n30) );
  OR2X1 r793_U27 ( .IN2(n9813), .IN1(n6751), .Q(r793_n26) );
  NAND2X0 r793_U26 ( .IN1(n9813), .IN2(n6751), .QN(r793_n27) );
  NAND2X0 r793_U25 ( .IN1(r793_n26), .IN2(r793_n27), .QN(r793_n25) );
  NOR2X0 r793_U24 ( .QN(r793_n22), .IN1(r793_n24), .IN2(r793_n25) );
  AND2X1 r793_U23 ( .IN1(r793_n24), .IN2(r793_n25), .Q(r793_n23) );
  NOR2X0 r793_U22 ( .QN(n184), .IN1(r793_n22), .IN2(r793_n23) );
  OR2X1 r793_U20 ( .IN2(n9809), .IN1(n6746), .Q(r793_n19) );
  NAND2X0 r793_U19 ( .IN1(n9809), .IN2(n6746), .QN(r793_n20) );
  NAND2X0 r793_U18 ( .IN1(r793_n19), .IN2(r793_n20), .QN(r793_n18) );
  NOR2X0 r793_U17 ( .QN(r793_n15), .IN1(r793_n17), .IN2(r793_n18) );
  AND2X1 r793_U16 ( .IN1(r793_n17), .IN2(r793_n18), .Q(r793_n16) );
  NOR2X0 r793_U15 ( .QN(n183), .IN1(r793_n15), .IN2(r793_n16) );
  OR2X1 r793_U13 ( .IN2(n9805), .IN1(n6750), .Q(r793_n12) );
  NAND2X0 r793_U12 ( .IN1(n9805), .IN2(n6750), .QN(r793_n13) );
  NAND2X0 r793_U11 ( .IN1(r793_n12), .IN2(r793_n13), .QN(r793_n11) );
  NOR2X0 r793_U10 ( .QN(r793_n8), .IN1(r793_n10), .IN2(r793_n11) );
  AND2X1 r793_U9 ( .IN1(r793_n10), .IN2(r793_n11), .Q(r793_n9) );
  NAND2X0 r793_U194 ( .IN1(n9825), .IN2(r793_n181), .QN(r793_n180) );
  NAND2X0 r793_U193 ( .IN1(r793_n179), .IN2(r793_n180), .QN(r793_n38) );
  NAND2X0 r793_U192 ( .IN1(P1_N359), .IN2(r793_n38), .QN(r793_n176) );
  OR2X1 r793_U191 ( .IN2(P1_N359), .IN1(r793_n38), .Q(r793_n178) );
  NAND2X0 r793_U190 ( .IN1(n9821), .IN2(r793_n178), .QN(r793_n177) );
  NAND2X0 r793_U189 ( .IN1(r793_n176), .IN2(r793_n177), .QN(r793_n31) );
  NAND2X0 r793_U188 ( .IN1(P1_N358), .IN2(r793_n31), .QN(r793_n173) );
  OR2X1 r793_U187 ( .IN2(P1_N358), .IN1(r793_n31), .Q(r793_n175) );
  NAND2X0 r793_U186 ( .IN1(n9817), .IN2(r793_n175), .QN(r793_n174) );
  NAND2X0 r793_U185 ( .IN1(r793_n173), .IN2(r793_n174), .QN(r793_n24) );
  NAND2X0 r793_U184 ( .IN1(P1_N357), .IN2(r793_n24), .QN(r793_n170) );
  OR2X1 r793_U183 ( .IN2(P1_N357), .IN1(r793_n24), .Q(r793_n172) );
  NAND2X0 r793_U182 ( .IN1(n9813), .IN2(r793_n172), .QN(r793_n171) );
  NAND2X0 r793_U181 ( .IN1(r793_n170), .IN2(r793_n171), .QN(r793_n17) );
  NAND2X0 r793_U180 ( .IN1(P1_N356), .IN2(r793_n17), .QN(r793_n167) );
  OR2X1 r793_U179 ( .IN2(P1_N356), .IN1(r793_n17), .Q(r793_n169) );
  NAND2X0 r793_U178 ( .IN1(n9809), .IN2(r793_n169), .QN(r793_n168) );
  NAND2X0 r793_U177 ( .IN1(r793_n167), .IN2(r793_n168), .QN(r793_n10) );
  NAND2X0 r793_U176 ( .IN1(P1_N355), .IN2(r793_n10), .QN(r793_n164) );
  OR2X1 r793_U175 ( .IN2(P1_N355), .IN1(r793_n10), .Q(r793_n166) );
  NAND2X0 r793_U174 ( .IN1(n9805), .IN2(r793_n166), .QN(r793_n165) );
  NAND2X0 r793_U173 ( .IN1(r793_n164), .IN2(r793_n165), .QN(r793_n3) );
  NAND2X0 r793_U172 ( .IN1(P1_N354), .IN2(r793_n3), .QN(r793_n161) );
  OR2X1 r793_U171 ( .IN2(P1_N354), .IN1(r793_n3), .Q(r793_n163) );
  NAND2X0 r793_U170 ( .IN1(n9801), .IN2(r793_n163), .QN(r793_n162) );
  NAND2X0 r793_U169 ( .IN1(r793_n161), .IN2(r793_n162), .QN(r793_n154) );
  OR2X1 r793_U167 ( .IN2(n9797), .IN1(n6759), .Q(r793_n158) );
  NAND2X0 r793_U166 ( .IN1(n9797), .IN2(n6759), .QN(r793_n159) );
  NAND2X0 r793_U165 ( .IN1(r793_n158), .IN2(r793_n159), .QN(r793_n157) );
  NOR2X0 r793_U164 ( .QN(r793_n155), .IN1(r793_n154), .IN2(r793_n157) );
  AND2X1 r793_U163 ( .IN1(r793_n154), .IN2(r793_n157), .Q(r793_n156) );
  NOR2X0 r793_U162 ( .QN(n180), .IN1(r793_n155), .IN2(r793_n156) );
  NAND2X0 r793_U161 ( .IN1(P1_N353), .IN2(r793_n154), .QN(r793_n151) );
  OR2X1 r793_U160 ( .IN2(P1_N353), .IN1(r793_n154), .Q(r793_n153) );
  NAND2X0 r793_U159 ( .IN1(n9797), .IN2(r793_n153), .QN(r793_n152) );
  NAND2X0 r793_U158 ( .IN1(r793_n151), .IN2(r793_n152), .QN(r793_n144) );
  OR2X1 r793_U156 ( .IN2(n9793), .IN1(n6754), .Q(r793_n148) );
  NAND2X0 r793_U155 ( .IN1(n9793), .IN2(n6754), .QN(r793_n149) );
  NAND2X0 r793_U154 ( .IN1(r793_n148), .IN2(r793_n149), .QN(r793_n147) );
  NOR2X0 r793_U153 ( .QN(r793_n145), .IN1(r793_n144), .IN2(r793_n147) );
  AND2X1 r793_U152 ( .IN1(r793_n144), .IN2(r793_n147), .Q(r793_n146) );
  NOR2X0 r793_U151 ( .QN(n179), .IN1(r793_n145), .IN2(r793_n146) );
  NAND2X0 r793_U150 ( .IN1(P1_N352), .IN2(r793_n144), .QN(r793_n141) );
  OR2X1 r793_U149 ( .IN2(P1_N352), .IN1(r793_n144), .Q(r793_n143) );
  NAND2X0 r793_U148 ( .IN1(n9793), .IN2(r793_n143), .QN(r793_n142) );
  NAND2X0 r793_U147 ( .IN1(r793_n141), .IN2(r793_n142), .QN(r793_n134) );
  OR2X1 r793_U145 ( .IN2(n9789), .IN1(n6758), .Q(r793_n138) );
  NAND2X0 r793_U144 ( .IN1(n9789), .IN2(n6758), .QN(r793_n139) );
  NAND2X0 r793_U143 ( .IN1(r793_n138), .IN2(r793_n139), .QN(r793_n137) );
  NOR2X0 r793_U142 ( .QN(r793_n135), .IN1(r793_n134), .IN2(r793_n137) );
  AND2X1 r793_U141 ( .IN1(r793_n134), .IN2(r793_n137), .Q(r793_n136) );
  NOR2X0 r793_U140 ( .QN(n178), .IN1(r793_n135), .IN2(r793_n136) );
  NAND2X0 r793_U139 ( .IN1(P1_N351), .IN2(r793_n134), .QN(r793_n131) );
  OR2X1 r793_U138 ( .IN2(P1_N351), .IN1(r793_n134), .Q(r793_n133) );
  NAND2X0 r793_U137 ( .IN1(n9789), .IN2(r793_n133), .QN(r793_n132) );
  NAND2X0 r793_U136 ( .IN1(r793_n131), .IN2(r793_n132), .QN(r793_n124) );
  OR2X1 r793_U134 ( .IN2(n9785), .IN1(n6763), .Q(r793_n128) );
  NAND2X0 r793_U133 ( .IN1(n9785), .IN2(n6763), .QN(r793_n129) );
  NAND2X0 r793_U132 ( .IN1(r793_n128), .IN2(r793_n129), .QN(r793_n127) );
  NOR2X0 r793_U131 ( .QN(r793_n125), .IN1(r793_n124), .IN2(r793_n127) );
  AND2X1 r793_U130 ( .IN1(r793_n124), .IN2(r793_n127), .Q(r793_n126) );
  NOR2X0 r793_U129 ( .QN(n177), .IN1(r793_n125), .IN2(r793_n126) );
  NAND2X0 r793_U128 ( .IN1(P1_N350), .IN2(r793_n124), .QN(r793_n121) );
  OR2X1 r793_U127 ( .IN2(P1_N350), .IN1(r793_n124), .Q(r793_n123) );
  NAND2X0 r793_U126 ( .IN1(n9785), .IN2(r793_n123), .QN(r793_n122) );
  NAND2X0 r793_U125 ( .IN1(r793_n121), .IN2(r793_n122), .QN(r793_n114) );
  OR2X1 r793_U123 ( .IN2(n9781), .IN1(n6767), .Q(r793_n118) );
  NAND2X0 r793_U122 ( .IN1(n9781), .IN2(n6767), .QN(r793_n119) );
  NAND2X0 r793_U121 ( .IN1(r793_n118), .IN2(r793_n119), .QN(r793_n117) );
  NOR2X0 r793_U120 ( .QN(r793_n115), .IN1(r793_n114), .IN2(r793_n117) );
  AND2X1 r793_U119 ( .IN1(r793_n114), .IN2(r793_n117), .Q(r793_n116) );
  NOR2X0 r793_U118 ( .QN(n176), .IN1(r793_n115), .IN2(r793_n116) );
  NAND2X0 r793_U117 ( .IN1(P1_N349), .IN2(r793_n114), .QN(r793_n111) );
  OR2X1 r793_U116 ( .IN2(P1_N349), .IN1(r793_n114), .Q(r793_n113) );
  NAND2X0 r793_U115 ( .IN1(n9781), .IN2(r793_n113), .QN(r793_n112) );
  NAND2X0 r793_U114 ( .IN1(r793_n111), .IN2(r793_n112), .QN(r793_n104) );
  OR2X1 r793_U112 ( .IN2(n9777), .IN1(n6762), .Q(r793_n108) );
  NAND2X0 r793_U111 ( .IN1(n9777), .IN2(n6762), .QN(r793_n109) );
  NAND2X0 r793_U110 ( .IN1(r793_n108), .IN2(r793_n109), .QN(r793_n107) );
  NOR2X0 r793_U109 ( .QN(r793_n105), .IN1(r793_n104), .IN2(r793_n107) );
  AND2X1 r793_U108 ( .IN1(r793_n104), .IN2(r793_n107), .Q(r793_n106) );
  NOR2X0 r793_U107 ( .QN(n175), .IN1(r793_n105), .IN2(r793_n106) );
  NAND2X0 r793_U106 ( .IN1(P1_N348), .IN2(r793_n104), .QN(r793_n101) );
  OR2X1 r793_U105 ( .IN2(P1_N348), .IN1(r793_n104), .Q(r793_n103) );
  NAND2X0 r793_U104 ( .IN1(n9777), .IN2(r793_n103), .QN(r793_n102) );
  NAND2X0 r793_U103 ( .IN1(r793_n101), .IN2(r793_n102), .QN(r793_n94) );
  OR2X1 r793_U209 ( .IN2(n920), .IN1(n6730), .Q(r793_n188) );
  NAND2X0 r793_U208 ( .IN1(n920), .IN2(n6730), .QN(r793_n189) );
  NAND2X0 r793_U207 ( .IN1(r793_n188), .IN2(r793_n189), .QN(n190) );
  NAND2X0 r793_U205 ( .IN1(n920), .IN2(P1_N363), .QN(r793_n60) );
  OR2X1 r793_U204 ( .IN2(r793_n60), .IN1(n6732), .Q(r793_n185) );
  NAND2X0 r793_U203 ( .IN1(n6732), .IN2(r793_n60), .QN(r793_n187) );
  NAND2X0 r793_U202 ( .IN1(n9833), .IN2(r793_n187), .QN(r793_n186) );
  NAND2X0 r793_U201 ( .IN1(r793_n185), .IN2(r793_n186), .QN(r793_n52) );
  NAND2X0 r793_U200 ( .IN1(P1_N361), .IN2(r793_n52), .QN(r793_n182) );
  OR2X1 r793_U199 ( .IN2(P1_N361), .IN1(r793_n52), .Q(r793_n184) );
  NAND2X0 r793_U198 ( .IN1(n9829), .IN2(r793_n184), .QN(r793_n183) );
  NAND2X0 r793_U197 ( .IN1(r793_n182), .IN2(r793_n183), .QN(r793_n45) );
  NAND2X0 r793_U196 ( .IN1(P1_N360), .IN2(r793_n45), .QN(r793_n179) );
  OR2X1 r793_U195 ( .IN2(P1_N360), .IN1(r793_n45), .Q(r793_n181) );
  NAND2X0 add_1104_U335 ( .IN1(add_1104_n184), .IN2(add_1104_n181), 
        .QN(add_1104_n307) );
  OR2X1 add_1104_U336 ( .IN2(add_1104_n181), .IN1(add_1104_n184), 
        .Q(add_1104_n305) );
  NAND2X0 add_1104_U337 ( .IN1(si_0_), .IN2(n9389), .QN(add_1104_n181) );
  INVX0 add_1104_U338 ( .ZN(add_1104_n184), .INP(n9337) );
  NAND2X0 add_1104_U339 ( .IN1(add_1104_n308), .IN2(add_1104_n309), .QN(N7) );
  NAND2X0 add_1104_U340 ( .IN1(si_0_), .IN2(add_1104_n310), .QN(add_1104_n309)
         );
  OR2X1 add_1104_U341 ( .IN2(si_0_), .IN1(add_1104_n310), .Q(add_1104_n308) );
  INVX0 add_1104_U342 ( .ZN(add_1104_n310), .INP(n9389) );
  OR2X1 add_1104_U327 ( .IN2(n9927), .IN1(add_1104_n45), .Q(add_1104_n301) );
  NAND2X0 add_1104_U328 ( .IN1(n9927), .IN2(add_1104_n45), .QN(add_1104_n299)
         );
  NAND2X0 add_1104_U329 ( .IN1(add_1104_n302), .IN2(add_1104_n303), 
        .QN(add_1104_n45) );
  NAND2X0 add_1104_U330 ( .IN1(si_2_), .IN2(add_1104_n304), .QN(add_1104_n303)
         );
  OR2X1 add_1104_U331 ( .IN2(n9931), .IN1(add_1104_n73), .Q(add_1104_n304) );
  NAND2X0 add_1104_U332 ( .IN1(n9931), .IN2(add_1104_n73), .QN(add_1104_n302)
         );
  NAND2X0 add_1104_U333 ( .IN1(add_1104_n305), .IN2(add_1104_n306), 
        .QN(add_1104_n73) );
  NAND2X0 add_1104_U334 ( .IN1(si_1_), .IN2(add_1104_n307), .QN(add_1104_n306)
         );
  OR2X1 add_1104_U319 ( .IN2(n9919), .IN1(add_1104_n31), .Q(add_1104_n295) );
  NAND2X0 add_1104_U320 ( .IN1(n9919), .IN2(add_1104_n31), .QN(add_1104_n293)
         );
  NAND2X0 add_1104_U321 ( .IN1(add_1104_n296), .IN2(add_1104_n297), 
        .QN(add_1104_n31) );
  NAND2X0 add_1104_U322 ( .IN1(si_4_), .IN2(add_1104_n298), .QN(add_1104_n297)
         );
  OR2X1 add_1104_U323 ( .IN2(n9923), .IN1(add_1104_n38), .Q(add_1104_n298) );
  NAND2X0 add_1104_U324 ( .IN1(n9923), .IN2(add_1104_n38), .QN(add_1104_n296)
         );
  NAND2X0 add_1104_U325 ( .IN1(add_1104_n299), .IN2(add_1104_n300), 
        .QN(add_1104_n38) );
  NAND2X0 add_1104_U326 ( .IN1(si_3_), .IN2(add_1104_n301), .QN(add_1104_n300)
         );
  OR2X1 add_1104_U311 ( .IN2(n9911), .IN1(add_1104_n17), .Q(add_1104_n289) );
  NAND2X0 add_1104_U312 ( .IN1(n9911), .IN2(add_1104_n17), .QN(add_1104_n287)
         );
  NAND2X0 add_1104_U313 ( .IN1(add_1104_n290), .IN2(add_1104_n291), 
        .QN(add_1104_n17) );
  NAND2X0 add_1104_U314 ( .IN1(si_6_), .IN2(add_1104_n292), .QN(add_1104_n291)
         );
  OR2X1 add_1104_U315 ( .IN2(n9915), .IN1(add_1104_n24), .Q(add_1104_n292) );
  NAND2X0 add_1104_U316 ( .IN1(n9915), .IN2(add_1104_n24), .QN(add_1104_n290)
         );
  NAND2X0 add_1104_U317 ( .IN1(add_1104_n293), .IN2(add_1104_n294), 
        .QN(add_1104_n24) );
  NAND2X0 add_1104_U318 ( .IN1(si_5_), .IN2(add_1104_n295), .QN(add_1104_n294)
         );
  OR2X1 add_1104_U303 ( .IN2(n9903), .IN1(add_1104_n3), .Q(add_1104_n283) );
  NAND2X0 add_1104_U304 ( .IN1(n9903), .IN2(add_1104_n3), .QN(add_1104_n281)
         );
  NAND2X0 add_1104_U305 ( .IN1(add_1104_n284), .IN2(add_1104_n285), 
        .QN(add_1104_n3) );
  NAND2X0 add_1104_U306 ( .IN1(si_8_), .IN2(add_1104_n286), .QN(add_1104_n285)
         );
  OR2X1 add_1104_U307 ( .IN2(n9907), .IN1(add_1104_n10), .Q(add_1104_n286) );
  NAND2X0 add_1104_U308 ( .IN1(n9907), .IN2(add_1104_n10), .QN(add_1104_n284)
         );
  NAND2X0 add_1104_U309 ( .IN1(add_1104_n287), .IN2(add_1104_n288), 
        .QN(add_1104_n10) );
  NAND2X0 add_1104_U310 ( .IN1(si_7_), .IN2(add_1104_n289), .QN(add_1104_n288)
         );
  AND2X1 add_1104_U295 ( .IN1(add_1104_n274), .IN2(add_1104_n277), 
        .Q(add_1104_n276) );
  NOR2X0 add_1104_U296 ( .QN(add_1104_n275), .IN1(add_1104_n274), 
        .IN2(add_1104_n277) );
  NAND2X0 add_1104_U297 ( .IN1(add_1104_n278), .IN2(add_1104_n279), 
        .QN(add_1104_n277) );
  NAND2X0 add_1104_U298 ( .IN1(si_10_), .IN2(add_1104_n280), 
        .QN(add_1104_n279) );
  OR2X1 add_1104_U299 ( .IN2(si_10_), .IN1(add_1104_n280), .Q(add_1104_n278)
         );
  INVX0 add_1104_U300 ( .ZN(add_1104_n280), .INP(n10091) );
  NAND2X0 add_1104_U301 ( .IN1(add_1104_n281), .IN2(add_1104_n282), 
        .QN(add_1104_n274) );
  NAND2X0 add_1104_U302 ( .IN1(si_9_), .IN2(add_1104_n283), .QN(add_1104_n282)
         );
  NAND2X0 add_1104_U287 ( .IN1(si_11_), .IN2(add_1104_n270), 
        .QN(add_1104_n269) );
  OR2X1 add_1104_U288 ( .IN2(si_11_), .IN1(add_1104_n270), .Q(add_1104_n268)
         );
  INVX0 add_1104_U289 ( .ZN(add_1104_n270), .INP(n10087) );
  NAND2X0 add_1104_U290 ( .IN1(add_1104_n271), .IN2(add_1104_n272), 
        .QN(add_1104_n264) );
  NAND2X0 add_1104_U291 ( .IN1(si_10_), .IN2(add_1104_n273), 
        .QN(add_1104_n272) );
  OR2X1 add_1104_U292 ( .IN2(n10091), .IN1(add_1104_n274), .Q(add_1104_n273)
         );
  NAND2X0 add_1104_U293 ( .IN1(n10091), .IN2(add_1104_n274), 
        .QN(add_1104_n271) );
  NOR2X0 add_1104_U294 ( .QN(N17), .IN1(add_1104_n275), .IN2(add_1104_n276) );
  NAND2X0 add_1104_U279 ( .IN1(add_1104_n261), .IN2(add_1104_n262), 
        .QN(add_1104_n254) );
  NAND2X0 add_1104_U280 ( .IN1(si_11_), .IN2(add_1104_n263), 
        .QN(add_1104_n262) );
  OR2X1 add_1104_U281 ( .IN2(n10087), .IN1(add_1104_n264), .Q(add_1104_n263)
         );
  NAND2X0 add_1104_U282 ( .IN1(n10087), .IN2(add_1104_n264), 
        .QN(add_1104_n261) );
  NOR2X0 add_1104_U283 ( .QN(N18), .IN1(add_1104_n265), .IN2(add_1104_n266) );
  AND2X1 add_1104_U284 ( .IN1(add_1104_n264), .IN2(add_1104_n267), 
        .Q(add_1104_n266) );
  NOR2X0 add_1104_U285 ( .QN(add_1104_n265), .IN1(add_1104_n264), 
        .IN2(add_1104_n267) );
  NAND2X0 add_1104_U286 ( .IN1(add_1104_n268), .IN2(add_1104_n269), 
        .QN(add_1104_n267) );
  NAND2X0 add_1104_U271 ( .IN1(n10083), .IN2(add_1104_n254), 
        .QN(add_1104_n251) );
  NOR2X0 add_1104_U272 ( .QN(N19), .IN1(add_1104_n255), .IN2(add_1104_n256) );
  AND2X1 add_1104_U273 ( .IN1(add_1104_n254), .IN2(add_1104_n257), 
        .Q(add_1104_n256) );
  NOR2X0 add_1104_U274 ( .QN(add_1104_n255), .IN1(add_1104_n254), 
        .IN2(add_1104_n257) );
  NAND2X0 add_1104_U275 ( .IN1(add_1104_n258), .IN2(add_1104_n259), 
        .QN(add_1104_n257) );
  NAND2X0 add_1104_U276 ( .IN1(si_12_), .IN2(add_1104_n260), 
        .QN(add_1104_n259) );
  OR2X1 add_1104_U277 ( .IN2(si_12_), .IN1(add_1104_n260), .Q(add_1104_n258)
         );
  INVX0 add_1104_U278 ( .ZN(add_1104_n260), .INP(n10083) );
  NOR2X0 add_1104_U263 ( .QN(add_1104_n245), .IN1(add_1104_n244), 
        .IN2(add_1104_n247) );
  NAND2X0 add_1104_U264 ( .IN1(add_1104_n248), .IN2(add_1104_n249), 
        .QN(add_1104_n247) );
  NAND2X0 add_1104_U265 ( .IN1(si_13_), .IN2(add_1104_n250), 
        .QN(add_1104_n249) );
  OR2X1 add_1104_U266 ( .IN2(si_13_), .IN1(add_1104_n250), .Q(add_1104_n248)
         );
  INVX0 add_1104_U267 ( .ZN(add_1104_n250), .INP(n10079) );
  NAND2X0 add_1104_U268 ( .IN1(add_1104_n251), .IN2(add_1104_n252), 
        .QN(add_1104_n244) );
  NAND2X0 add_1104_U269 ( .IN1(si_12_), .IN2(add_1104_n253), 
        .QN(add_1104_n252) );
  OR2X1 add_1104_U270 ( .IN2(n10083), .IN1(add_1104_n254), .Q(add_1104_n253)
         );
  OR2X1 add_1104_U255 ( .IN2(si_14_), .IN1(add_1104_n240), .Q(add_1104_n238)
         );
  INVX0 add_1104_U256 ( .ZN(add_1104_n240), .INP(n10075) );
  NAND2X0 add_1104_U257 ( .IN1(add_1104_n241), .IN2(add_1104_n242), 
        .QN(add_1104_n234) );
  NAND2X0 add_1104_U258 ( .IN1(si_13_), .IN2(add_1104_n243), 
        .QN(add_1104_n242) );
  OR2X1 add_1104_U259 ( .IN2(n10079), .IN1(add_1104_n244), .Q(add_1104_n243)
         );
  NAND2X0 add_1104_U260 ( .IN1(n10079), .IN2(add_1104_n244), 
        .QN(add_1104_n241) );
  NOR2X0 add_1104_U261 ( .QN(N20), .IN1(add_1104_n245), .IN2(add_1104_n246) );
  AND2X1 add_1104_U262 ( .IN1(add_1104_n244), .IN2(add_1104_n247), 
        .Q(add_1104_n246) );
  NAND2X0 add_1104_U247 ( .IN1(si_14_), .IN2(add_1104_n233), 
        .QN(add_1104_n232) );
  OR2X1 add_1104_U248 ( .IN2(n10075), .IN1(add_1104_n234), .Q(add_1104_n233)
         );
  NAND2X0 add_1104_U249 ( .IN1(n10075), .IN2(add_1104_n234), 
        .QN(add_1104_n231) );
  NOR2X0 add_1104_U250 ( .QN(N21), .IN1(add_1104_n235), .IN2(add_1104_n236) );
  AND2X1 add_1104_U251 ( .IN1(add_1104_n234), .IN2(add_1104_n237), 
        .Q(add_1104_n236) );
  NOR2X0 add_1104_U252 ( .QN(add_1104_n235), .IN1(add_1104_n234), 
        .IN2(add_1104_n237) );
  NAND2X0 add_1104_U253 ( .IN1(add_1104_n238), .IN2(add_1104_n239), 
        .QN(add_1104_n237) );
  NAND2X0 add_1104_U254 ( .IN1(si_14_), .IN2(add_1104_n240), 
        .QN(add_1104_n239) );
  NOR2X0 add_1104_U239 ( .QN(N22), .IN1(add_1104_n225), .IN2(add_1104_n226) );
  AND2X1 add_1104_U240 ( .IN1(add_1104_n224), .IN2(add_1104_n227), 
        .Q(add_1104_n226) );
  NOR2X0 add_1104_U241 ( .QN(add_1104_n225), .IN1(add_1104_n224), 
        .IN2(add_1104_n227) );
  NAND2X0 add_1104_U242 ( .IN1(add_1104_n228), .IN2(add_1104_n229), 
        .QN(add_1104_n227) );
  NAND2X0 add_1104_U243 ( .IN1(si_15_), .IN2(add_1104_n230), 
        .QN(add_1104_n229) );
  OR2X1 add_1104_U244 ( .IN2(si_15_), .IN1(add_1104_n230), .Q(add_1104_n228)
         );
  INVX0 add_1104_U245 ( .ZN(add_1104_n230), .INP(n10071) );
  NAND2X0 add_1104_U246 ( .IN1(add_1104_n231), .IN2(add_1104_n232), 
        .QN(add_1104_n224) );
  NAND2X0 add_1104_U231 ( .IN1(add_1104_n218), .IN2(add_1104_n219), 
        .QN(add_1104_n217) );
  NAND2X0 add_1104_U232 ( .IN1(si_16_), .IN2(add_1104_n220), 
        .QN(add_1104_n219) );
  OR2X1 add_1104_U233 ( .IN2(si_16_), .IN1(add_1104_n220), .Q(add_1104_n218)
         );
  INVX0 add_1104_U234 ( .ZN(add_1104_n220), .INP(n10067) );
  NAND2X0 add_1104_U235 ( .IN1(add_1104_n221), .IN2(add_1104_n222), 
        .QN(add_1104_n214) );
  NAND2X0 add_1104_U236 ( .IN1(si_15_), .IN2(add_1104_n223), 
        .QN(add_1104_n222) );
  OR2X1 add_1104_U237 ( .IN2(n10071), .IN1(add_1104_n224), .Q(add_1104_n223)
         );
  NAND2X0 add_1104_U238 ( .IN1(n10071), .IN2(add_1104_n224), 
        .QN(add_1104_n221) );
  INVX0 add_1104_U223 ( .ZN(add_1104_n210), .INP(n10063) );
  NAND2X0 add_1104_U224 ( .IN1(add_1104_n211), .IN2(add_1104_n212), 
        .QN(add_1104_n204) );
  NAND2X0 add_1104_U225 ( .IN1(si_16_), .IN2(add_1104_n213), 
        .QN(add_1104_n212) );
  OR2X1 add_1104_U226 ( .IN2(n10067), .IN1(add_1104_n214), .Q(add_1104_n213)
         );
  NAND2X0 add_1104_U227 ( .IN1(n10067), .IN2(add_1104_n214), 
        .QN(add_1104_n211) );
  NOR2X0 add_1104_U228 ( .QN(N23), .IN1(add_1104_n215), .IN2(add_1104_n216) );
  AND2X1 add_1104_U229 ( .IN1(add_1104_n214), .IN2(add_1104_n217), 
        .Q(add_1104_n216) );
  NOR2X0 add_1104_U230 ( .QN(add_1104_n215), .IN1(add_1104_n214), 
        .IN2(add_1104_n217) );
  OR2X1 add_1104_U215 ( .IN2(n10063), .IN1(add_1104_n204), .Q(add_1104_n203)
         );
  NAND2X0 add_1104_U216 ( .IN1(n10063), .IN2(add_1104_n204), 
        .QN(add_1104_n201) );
  NOR2X0 add_1104_U217 ( .QN(N24), .IN1(add_1104_n205), .IN2(add_1104_n206) );
  AND2X1 add_1104_U218 ( .IN1(add_1104_n204), .IN2(add_1104_n207), 
        .Q(add_1104_n206) );
  NOR2X0 add_1104_U219 ( .QN(add_1104_n205), .IN1(add_1104_n204), 
        .IN2(add_1104_n207) );
  NAND2X0 add_1104_U220 ( .IN1(add_1104_n208), .IN2(add_1104_n209), 
        .QN(add_1104_n207) );
  NAND2X0 add_1104_U221 ( .IN1(si_17_), .IN2(add_1104_n210), 
        .QN(add_1104_n209) );
  OR2X1 add_1104_U222 ( .IN2(si_17_), .IN1(add_1104_n210), .Q(add_1104_n208)
         );
  AND2X1 add_1104_U207 ( .IN1(add_1104_n194), .IN2(add_1104_n197), 
        .Q(add_1104_n196) );
  NOR2X0 add_1104_U208 ( .QN(add_1104_n195), .IN1(add_1104_n194), 
        .IN2(add_1104_n197) );
  NAND2X0 add_1104_U209 ( .IN1(add_1104_n198), .IN2(add_1104_n199), 
        .QN(add_1104_n197) );
  NAND2X0 add_1104_U210 ( .IN1(si_18_), .IN2(add_1104_n200), 
        .QN(add_1104_n199) );
  OR2X1 add_1104_U211 ( .IN2(si_18_), .IN1(add_1104_n200), .Q(add_1104_n198)
         );
  INVX0 add_1104_U212 ( .ZN(add_1104_n200), .INP(n10059) );
  NAND2X0 add_1104_U213 ( .IN1(add_1104_n201), .IN2(add_1104_n202), 
        .QN(add_1104_n194) );
  NAND2X0 add_1104_U214 ( .IN1(si_17_), .IN2(add_1104_n203), 
        .QN(add_1104_n202) );
  NAND2X0 add_1104_U199 ( .IN1(si_19_), .IN2(add_1104_n190), 
        .QN(add_1104_n189) );
  OR2X1 add_1104_U200 ( .IN2(si_19_), .IN1(add_1104_n190), .Q(add_1104_n188)
         );
  INVX0 add_1104_U201 ( .ZN(add_1104_n190), .INP(n10055) );
  NAND2X0 add_1104_U202 ( .IN1(add_1104_n191), .IN2(add_1104_n192), 
        .QN(add_1104_n177) );
  NAND2X0 add_1104_U203 ( .IN1(si_18_), .IN2(add_1104_n193), 
        .QN(add_1104_n192) );
  OR2X1 add_1104_U204 ( .IN2(n10059), .IN1(add_1104_n194), .Q(add_1104_n193)
         );
  NAND2X0 add_1104_U205 ( .IN1(n10059), .IN2(add_1104_n194), 
        .QN(add_1104_n191) );
  NOR2X0 add_1104_U206 ( .QN(N25), .IN1(add_1104_n195), .IN2(add_1104_n196) );
  NAND2X0 add_1104_U191 ( .IN1(add_1104_n180), .IN2(add_1104_n181), 
        .QN(add_1104_n178) );
  NAND2X0 add_1104_U192 ( .IN1(add_1104_n182), .IN2(add_1104_n183), 
        .QN(add_1104_n180) );
  NAND2X0 add_1104_U193 ( .IN1(si_1_), .IN2(add_1104_n184), .QN(add_1104_n183)
         );
  OR2X1 add_1104_U194 ( .IN2(si_1_), .IN1(add_1104_n184), .Q(add_1104_n182) );
  NOR2X0 add_1104_U195 ( .QN(N26), .IN1(add_1104_n185), .IN2(add_1104_n186) );
  AND2X1 add_1104_U196 ( .IN1(add_1104_n177), .IN2(add_1104_n187), 
        .Q(add_1104_n186) );
  NOR2X0 add_1104_U197 ( .QN(add_1104_n185), .IN1(add_1104_n177), 
        .IN2(add_1104_n187) );
  NAND2X0 add_1104_U198 ( .IN1(add_1104_n188), .IN2(add_1104_n189), 
        .QN(add_1104_n187) );
  OR2X1 add_1104_U183 ( .IN2(si_20_), .IN1(add_1104_n173), .Q(add_1104_n171)
         );
  INVX0 add_1104_U184 ( .ZN(add_1104_n173), .INP(n10051) );
  NAND2X0 add_1104_U185 ( .IN1(add_1104_n174), .IN2(add_1104_n175), 
        .QN(add_1104_n167) );
  NAND2X0 add_1104_U186 ( .IN1(si_19_), .IN2(add_1104_n176), 
        .QN(add_1104_n175) );
  OR2X1 add_1104_U187 ( .IN2(n10055), .IN1(add_1104_n177), .Q(add_1104_n176)
         );
  NAND2X0 add_1104_U188 ( .IN1(n10055), .IN2(add_1104_n177), 
        .QN(add_1104_n174) );
  NAND2X0 add_1104_U189 ( .IN1(add_1104_n178), .IN2(add_1104_n179), .QN(N8) );
  OR2X1 add_1104_U190 ( .IN2(add_1104_n181), .IN1(add_1104_n180), 
        .Q(add_1104_n179) );
  NAND2X0 add_1104_U175 ( .IN1(si_20_), .IN2(add_1104_n166), 
        .QN(add_1104_n165) );
  OR2X1 add_1104_U176 ( .IN2(n10051), .IN1(add_1104_n167), .Q(add_1104_n166)
         );
  NAND2X0 add_1104_U177 ( .IN1(n10051), .IN2(add_1104_n167), 
        .QN(add_1104_n164) );
  NOR2X0 add_1104_U178 ( .QN(N27), .IN1(add_1104_n168), .IN2(add_1104_n169) );
  AND2X1 add_1104_U179 ( .IN1(add_1104_n167), .IN2(add_1104_n170), 
        .Q(add_1104_n169) );
  NOR2X0 add_1104_U180 ( .QN(add_1104_n168), .IN1(add_1104_n167), 
        .IN2(add_1104_n170) );
  NAND2X0 add_1104_U181 ( .IN1(add_1104_n171), .IN2(add_1104_n172), 
        .QN(add_1104_n170) );
  NAND2X0 add_1104_U182 ( .IN1(si_20_), .IN2(add_1104_n173), 
        .QN(add_1104_n172) );
  NOR2X0 add_1104_U167 ( .QN(N28), .IN1(add_1104_n158), .IN2(add_1104_n159) );
  AND2X1 add_1104_U168 ( .IN1(add_1104_n157), .IN2(add_1104_n160), 
        .Q(add_1104_n159) );
  NOR2X0 add_1104_U169 ( .QN(add_1104_n158), .IN1(add_1104_n157), 
        .IN2(add_1104_n160) );
  NAND2X0 add_1104_U170 ( .IN1(add_1104_n161), .IN2(add_1104_n162), 
        .QN(add_1104_n160) );
  NAND2X0 add_1104_U171 ( .IN1(si_21_), .IN2(add_1104_n163), 
        .QN(add_1104_n162) );
  OR2X1 add_1104_U172 ( .IN2(si_21_), .IN1(add_1104_n163), .Q(add_1104_n161)
         );
  INVX0 add_1104_U173 ( .ZN(add_1104_n163), .INP(n10047) );
  NAND2X0 add_1104_U174 ( .IN1(add_1104_n164), .IN2(add_1104_n165), 
        .QN(add_1104_n157) );
  NAND2X0 add_1104_U159 ( .IN1(add_1104_n151), .IN2(add_1104_n152), 
        .QN(add_1104_n150) );
  NAND2X0 add_1104_U160 ( .IN1(si_22_), .IN2(add_1104_n153), 
        .QN(add_1104_n152) );
  OR2X1 add_1104_U161 ( .IN2(si_22_), .IN1(add_1104_n153), .Q(add_1104_n151)
         );
  INVX0 add_1104_U162 ( .ZN(add_1104_n153), .INP(n10043) );
  NAND2X0 add_1104_U163 ( .IN1(add_1104_n154), .IN2(add_1104_n155), 
        .QN(add_1104_n147) );
  NAND2X0 add_1104_U164 ( .IN1(si_21_), .IN2(add_1104_n156), 
        .QN(add_1104_n155) );
  OR2X1 add_1104_U165 ( .IN2(n10047), .IN1(add_1104_n157), .Q(add_1104_n156)
         );
  NAND2X0 add_1104_U166 ( .IN1(n10047), .IN2(add_1104_n157), 
        .QN(add_1104_n154) );
  INVX0 add_1104_U151 ( .ZN(add_1104_n143), .INP(n10039) );
  NAND2X0 add_1104_U152 ( .IN1(add_1104_n144), .IN2(add_1104_n145), 
        .QN(add_1104_n137) );
  NAND2X0 add_1104_U153 ( .IN1(si_22_), .IN2(add_1104_n146), 
        .QN(add_1104_n145) );
  OR2X1 add_1104_U154 ( .IN2(n10043), .IN1(add_1104_n147), .Q(add_1104_n146)
         );
  NAND2X0 add_1104_U155 ( .IN1(n10043), .IN2(add_1104_n147), 
        .QN(add_1104_n144) );
  NOR2X0 add_1104_U156 ( .QN(N29), .IN1(add_1104_n148), .IN2(add_1104_n149) );
  AND2X1 add_1104_U157 ( .IN1(add_1104_n147), .IN2(add_1104_n150), 
        .Q(add_1104_n149) );
  NOR2X0 add_1104_U158 ( .QN(add_1104_n148), .IN1(add_1104_n147), 
        .IN2(add_1104_n150) );
  OR2X1 add_1104_U143 ( .IN2(n10039), .IN1(add_1104_n137), .Q(add_1104_n136)
         );
  NAND2X0 add_1104_U144 ( .IN1(n10039), .IN2(add_1104_n137), 
        .QN(add_1104_n134) );
  NOR2X0 add_1104_U145 ( .QN(N30), .IN1(add_1104_n138), .IN2(add_1104_n139) );
  AND2X1 add_1104_U146 ( .IN1(add_1104_n137), .IN2(add_1104_n140), 
        .Q(add_1104_n139) );
  NOR2X0 add_1104_U147 ( .QN(add_1104_n138), .IN1(add_1104_n137), 
        .IN2(add_1104_n140) );
  NAND2X0 add_1104_U148 ( .IN1(add_1104_n141), .IN2(add_1104_n142), 
        .QN(add_1104_n140) );
  NAND2X0 add_1104_U149 ( .IN1(si_23_), .IN2(add_1104_n143), 
        .QN(add_1104_n142) );
  OR2X1 add_1104_U150 ( .IN2(si_23_), .IN1(add_1104_n143), .Q(add_1104_n141)
         );
  AND2X1 add_1104_U135 ( .IN1(add_1104_n127), .IN2(add_1104_n130), 
        .Q(add_1104_n129) );
  NOR2X0 add_1104_U136 ( .QN(add_1104_n128), .IN1(add_1104_n127), 
        .IN2(add_1104_n130) );
  NAND2X0 add_1104_U137 ( .IN1(add_1104_n131), .IN2(add_1104_n132), 
        .QN(add_1104_n130) );
  NAND2X0 add_1104_U138 ( .IN1(si_24_), .IN2(add_1104_n133), 
        .QN(add_1104_n132) );
  OR2X1 add_1104_U139 ( .IN2(si_24_), .IN1(add_1104_n133), .Q(add_1104_n131)
         );
  INVX0 add_1104_U140 ( .ZN(add_1104_n133), .INP(n10035) );
  NAND2X0 add_1104_U141 ( .IN1(add_1104_n134), .IN2(add_1104_n135), 
        .QN(add_1104_n127) );
  NAND2X0 add_1104_U142 ( .IN1(si_23_), .IN2(add_1104_n136), 
        .QN(add_1104_n135) );
  NAND2X0 add_1104_U127 ( .IN1(si_25_), .IN2(add_1104_n123), 
        .QN(add_1104_n122) );
  OR2X1 add_1104_U128 ( .IN2(si_25_), .IN1(add_1104_n123), .Q(add_1104_n121)
         );
  INVX0 add_1104_U129 ( .ZN(add_1104_n123), .INP(n10031) );
  NAND2X0 add_1104_U130 ( .IN1(add_1104_n124), .IN2(add_1104_n125), 
        .QN(add_1104_n117) );
  NAND2X0 add_1104_U131 ( .IN1(si_24_), .IN2(add_1104_n126), 
        .QN(add_1104_n125) );
  OR2X1 add_1104_U132 ( .IN2(n10035), .IN1(add_1104_n127), .Q(add_1104_n126)
         );
  NAND2X0 add_1104_U133 ( .IN1(n10035), .IN2(add_1104_n127), 
        .QN(add_1104_n124) );
  NOR2X0 add_1104_U134 ( .QN(N31), .IN1(add_1104_n128), .IN2(add_1104_n129) );
  NAND2X0 add_1104_U119 ( .IN1(add_1104_n114), .IN2(add_1104_n115), 
        .QN(add_1104_n107) );
  NAND2X0 add_1104_U120 ( .IN1(si_25_), .IN2(add_1104_n116), 
        .QN(add_1104_n115) );
  OR2X1 add_1104_U121 ( .IN2(n10031), .IN1(add_1104_n117), .Q(add_1104_n116)
         );
  NAND2X0 add_1104_U122 ( .IN1(n10031), .IN2(add_1104_n117), 
        .QN(add_1104_n114) );
  NOR2X0 add_1104_U123 ( .QN(N32), .IN1(add_1104_n118), .IN2(add_1104_n119) );
  AND2X1 add_1104_U124 ( .IN1(add_1104_n117), .IN2(add_1104_n120), 
        .Q(add_1104_n119) );
  NOR2X0 add_1104_U125 ( .QN(add_1104_n118), .IN1(add_1104_n117), 
        .IN2(add_1104_n120) );
  NAND2X0 add_1104_U126 ( .IN1(add_1104_n121), .IN2(add_1104_n122), 
        .QN(add_1104_n120) );
  NAND2X0 add_1104_U111 ( .IN1(n10027), .IN2(add_1104_n107), 
        .QN(add_1104_n104) );
  NOR2X0 add_1104_U112 ( .QN(N33), .IN1(add_1104_n108), .IN2(add_1104_n109) );
  AND2X1 add_1104_U113 ( .IN1(add_1104_n107), .IN2(add_1104_n110), 
        .Q(add_1104_n109) );
  NOR2X0 add_1104_U114 ( .QN(add_1104_n108), .IN1(add_1104_n107), 
        .IN2(add_1104_n110) );
  NAND2X0 add_1104_U115 ( .IN1(add_1104_n111), .IN2(add_1104_n112), 
        .QN(add_1104_n110) );
  NAND2X0 add_1104_U116 ( .IN1(si_26_), .IN2(add_1104_n113), 
        .QN(add_1104_n112) );
  OR2X1 add_1104_U117 ( .IN2(si_26_), .IN1(add_1104_n113), .Q(add_1104_n111)
         );
  INVX0 add_1104_U118 ( .ZN(add_1104_n113), .INP(n10027) );
  NOR2X0 add_1104_U103 ( .QN(add_1104_n98), .IN1(add_1104_n97), 
        .IN2(add_1104_n100) );
  NAND2X0 add_1104_U104 ( .IN1(add_1104_n101), .IN2(add_1104_n102), 
        .QN(add_1104_n100) );
  NAND2X0 add_1104_U105 ( .IN1(si_27_), .IN2(add_1104_n103), 
        .QN(add_1104_n102) );
  OR2X1 add_1104_U106 ( .IN2(si_27_), .IN1(add_1104_n103), .Q(add_1104_n101)
         );
  INVX0 add_1104_U107 ( .ZN(add_1104_n103), .INP(n10023) );
  NAND2X0 add_1104_U108 ( .IN1(add_1104_n104), .IN2(add_1104_n105), 
        .QN(add_1104_n97) );
  NAND2X0 add_1104_U109 ( .IN1(si_26_), .IN2(add_1104_n106), 
        .QN(add_1104_n105) );
  OR2X1 add_1104_U110 ( .IN2(n10027), .IN1(add_1104_n107), .Q(add_1104_n106)
         );
  OR2X1 add_1104_U95 ( .IN2(si_28_), .IN1(add_1104_n93), .Q(add_1104_n91) );
  INVX0 add_1104_U96 ( .ZN(add_1104_n93), .INP(n10019) );
  NAND2X0 add_1104_U97 ( .IN1(add_1104_n94), .IN2(add_1104_n95), 
        .QN(add_1104_n87) );
  NAND2X0 add_1104_U98 ( .IN1(si_27_), .IN2(add_1104_n96), .QN(add_1104_n95)
         );
  OR2X1 add_1104_U99 ( .IN2(n10023), .IN1(add_1104_n97), .Q(add_1104_n96) );
  NAND2X0 add_1104_U100 ( .IN1(n10023), .IN2(add_1104_n97), .QN(add_1104_n94)
         );
  NOR2X0 add_1104_U101 ( .QN(N34), .IN1(add_1104_n98), .IN2(add_1104_n99) );
  AND2X1 add_1104_U102 ( .IN1(add_1104_n97), .IN2(add_1104_n100), 
        .Q(add_1104_n99) );
  NAND2X0 add_1104_U87 ( .IN1(si_28_), .IN2(add_1104_n86), .QN(add_1104_n85)
         );
  OR2X1 add_1104_U88 ( .IN2(n10019), .IN1(add_1104_n87), .Q(add_1104_n86) );
  NAND2X0 add_1104_U89 ( .IN1(n10019), .IN2(add_1104_n87), .QN(add_1104_n84)
         );
  NOR2X0 add_1104_U90 ( .QN(N35), .IN1(add_1104_n88), .IN2(add_1104_n89) );
  AND2X1 add_1104_U91 ( .IN1(add_1104_n87), .IN2(add_1104_n90), 
        .Q(add_1104_n89) );
  NOR2X0 add_1104_U92 ( .QN(add_1104_n88), .IN1(add_1104_n87), 
        .IN2(add_1104_n90) );
  NAND2X0 add_1104_U93 ( .IN1(add_1104_n91), .IN2(add_1104_n92), 
        .QN(add_1104_n90) );
  NAND2X0 add_1104_U94 ( .IN1(si_28_), .IN2(add_1104_n93), .QN(add_1104_n92)
         );
  NOR2X0 add_1104_U79 ( .QN(N36), .IN1(add_1104_n78), .IN2(add_1104_n79) );
  AND2X1 add_1104_U80 ( .IN1(add_1104_n70), .IN2(add_1104_n80), 
        .Q(add_1104_n79) );
  NOR2X0 add_1104_U81 ( .QN(add_1104_n78), .IN1(add_1104_n70), 
        .IN2(add_1104_n80) );
  NAND2X0 add_1104_U82 ( .IN1(add_1104_n81), .IN2(add_1104_n82), 
        .QN(add_1104_n80) );
  NAND2X0 add_1104_U83 ( .IN1(si_29_), .IN2(add_1104_n83), .QN(add_1104_n82)
         );
  OR2X1 add_1104_U84 ( .IN2(si_29_), .IN1(add_1104_n83), .Q(add_1104_n81) );
  INVX0 add_1104_U85 ( .ZN(add_1104_n83), .INP(n10099) );
  NAND2X0 add_1104_U86 ( .IN1(add_1104_n84), .IN2(add_1104_n85), 
        .QN(add_1104_n70) );
  NAND2X0 add_1104_U71 ( .IN1(n10099), .IN2(add_1104_n70), .QN(add_1104_n67)
         );
  NOR2X0 add_1104_U72 ( .QN(N9), .IN1(add_1104_n71), .IN2(add_1104_n72) );
  AND2X1 add_1104_U73 ( .IN1(add_1104_n73), .IN2(add_1104_n74), 
        .Q(add_1104_n72) );
  NOR2X0 add_1104_U74 ( .QN(add_1104_n71), .IN1(add_1104_n73), 
        .IN2(add_1104_n74) );
  NAND2X0 add_1104_U75 ( .IN1(add_1104_n75), .IN2(add_1104_n76), 
        .QN(add_1104_n74) );
  NAND2X0 add_1104_U76 ( .IN1(si_2_), .IN2(add_1104_n77), .QN(add_1104_n76) );
  OR2X1 add_1104_U77 ( .IN2(si_2_), .IN1(add_1104_n77), .Q(add_1104_n75) );
  INVX0 add_1104_U78 ( .ZN(add_1104_n77), .INP(n9931) );
  NOR2X0 add_1104_U63 ( .QN(add_1104_n61), .IN1(add_1104_n57), 
        .IN2(add_1104_n63) );
  NAND2X0 add_1104_U64 ( .IN1(add_1104_n64), .IN2(add_1104_n65), 
        .QN(add_1104_n63) );
  NAND2X0 add_1104_U65 ( .IN1(si_30_), .IN2(add_1104_n66), .QN(add_1104_n65)
         );
  OR2X1 add_1104_U66 ( .IN2(si_30_), .IN1(add_1104_n66), .Q(add_1104_n64) );
  INVX0 add_1104_U67 ( .ZN(add_1104_n66), .INP(n10107) );
  NAND2X0 add_1104_U68 ( .IN1(add_1104_n67), .IN2(add_1104_n68), 
        .QN(add_1104_n57) );
  NAND2X0 add_1104_U69 ( .IN1(si_29_), .IN2(add_1104_n69), .QN(add_1104_n68)
         );
  OR2X1 add_1104_U70 ( .IN2(n10099), .IN1(add_1104_n70), .Q(add_1104_n69) );
  OR2X1 add_1104_U55 ( .IN2(n10107), .IN1(add_1104_n57), .Q(add_1104_n56) );
  NAND2X0 add_1104_U56 ( .IN1(n10107), .IN2(add_1104_n57), .QN(add_1104_n54)
         );
  NAND2X0 add_1104_U57 ( .IN1(add_1104_n58), .IN2(add_1104_n59), 
        .QN(add_1104_n53) );
  NAND2X0 add_1104_U58 ( .IN1(si_31_), .IN2(add_1104_n60), .QN(add_1104_n59)
         );
  OR2X1 add_1104_U59 ( .IN2(si_31_), .IN1(add_1104_n60), .Q(add_1104_n58) );
  INVX0 add_1104_U60 ( .ZN(add_1104_n60), .INP(n9341) );
  NOR2X0 add_1104_U61 ( .QN(N37), .IN1(add_1104_n61), .IN2(add_1104_n62) );
  AND2X1 add_1104_U62 ( .IN1(add_1104_n57), .IN2(add_1104_n63), 
        .Q(add_1104_n62) );
  NAND2X0 add_1104_U47 ( .IN1(si_3_), .IN2(add_1104_n49), .QN(add_1104_n48) );
  OR2X1 add_1104_U48 ( .IN2(si_3_), .IN1(add_1104_n49), .Q(add_1104_n47) );
  INVX0 add_1104_U49 ( .ZN(add_1104_n49), .INP(n9927) );
  NOR2X0 add_1104_U50 ( .QN(N38), .IN1(add_1104_n50), .IN2(add_1104_n51) );
  AND2X1 add_1104_U51 ( .IN1(add_1104_n52), .IN2(add_1104_n53), 
        .Q(add_1104_n51) );
  NOR2X0 add_1104_U52 ( .QN(add_1104_n50), .IN1(add_1104_n53), 
        .IN2(add_1104_n52) );
  NAND2X0 add_1104_U53 ( .IN1(add_1104_n54), .IN2(add_1104_n55), 
        .QN(add_1104_n52) );
  NAND2X0 add_1104_U54 ( .IN1(si_30_), .IN2(add_1104_n56), .QN(add_1104_n55)
         );
  NAND2X0 add_1104_U39 ( .IN1(add_1104_n40), .IN2(add_1104_n41), 
        .QN(add_1104_n39) );
  NAND2X0 add_1104_U40 ( .IN1(si_4_), .IN2(add_1104_n42), .QN(add_1104_n41) );
  OR2X1 add_1104_U41 ( .IN2(si_4_), .IN1(add_1104_n42), .Q(add_1104_n40) );
  INVX0 add_1104_U42 ( .ZN(add_1104_n42), .INP(n9923) );
  NOR2X0 add_1104_U43 ( .QN(N10), .IN1(add_1104_n43), .IN2(add_1104_n44) );
  AND2X1 add_1104_U44 ( .IN1(add_1104_n45), .IN2(add_1104_n46), 
        .Q(add_1104_n44) );
  NOR2X0 add_1104_U45 ( .QN(add_1104_n43), .IN1(add_1104_n45), 
        .IN2(add_1104_n46) );
  NAND2X0 add_1104_U46 ( .IN1(add_1104_n47), .IN2(add_1104_n48), 
        .QN(add_1104_n46) );
  NOR2X0 add_1104_U31 ( .QN(add_1104_n29), .IN1(add_1104_n31), 
        .IN2(add_1104_n32) );
  NAND2X0 add_1104_U32 ( .IN1(add_1104_n33), .IN2(add_1104_n34), 
        .QN(add_1104_n32) );
  NAND2X0 add_1104_U33 ( .IN1(si_5_), .IN2(add_1104_n35), .QN(add_1104_n34) );
  OR2X1 add_1104_U34 ( .IN2(si_5_), .IN1(add_1104_n35), .Q(add_1104_n33) );
  INVX0 add_1104_U35 ( .ZN(add_1104_n35), .INP(n9919) );
  NOR2X0 add_1104_U36 ( .QN(N11), .IN1(add_1104_n36), .IN2(add_1104_n37) );
  AND2X1 add_1104_U37 ( .IN1(add_1104_n38), .IN2(add_1104_n39), 
        .Q(add_1104_n37) );
  NOR2X0 add_1104_U38 ( .QN(add_1104_n36), .IN1(add_1104_n38), 
        .IN2(add_1104_n39) );
  AND2X1 add_1104_U23 ( .IN1(add_1104_n24), .IN2(add_1104_n25), 
        .Q(add_1104_n23) );
  NOR2X0 add_1104_U24 ( .QN(add_1104_n22), .IN1(add_1104_n24), 
        .IN2(add_1104_n25) );
  NAND2X0 add_1104_U25 ( .IN1(add_1104_n26), .IN2(add_1104_n27), 
        .QN(add_1104_n25) );
  NAND2X0 add_1104_U26 ( .IN1(si_6_), .IN2(add_1104_n28), .QN(add_1104_n27) );
  OR2X1 add_1104_U27 ( .IN2(si_6_), .IN1(add_1104_n28), .Q(add_1104_n26) );
  INVX0 add_1104_U28 ( .ZN(add_1104_n28), .INP(n9915) );
  NOR2X0 add_1104_U29 ( .QN(N12), .IN1(add_1104_n29), .IN2(add_1104_n30) );
  AND2X1 add_1104_U30 ( .IN1(add_1104_n31), .IN2(add_1104_n32), 
        .Q(add_1104_n30) );
  NOR2X0 add_1104_U15 ( .QN(N14), .IN1(add_1104_n15), .IN2(add_1104_n16) );
  AND2X1 add_1104_U16 ( .IN1(add_1104_n17), .IN2(add_1104_n18), 
        .Q(add_1104_n16) );
  NOR2X0 add_1104_U17 ( .QN(add_1104_n15), .IN1(add_1104_n17), 
        .IN2(add_1104_n18) );
  NAND2X0 add_1104_U18 ( .IN1(add_1104_n19), .IN2(add_1104_n20), 
        .QN(add_1104_n18) );
  NAND2X0 add_1104_U19 ( .IN1(si_7_), .IN2(add_1104_n21), .QN(add_1104_n20) );
  OR2X1 add_1104_U20 ( .IN2(si_7_), .IN1(add_1104_n21), .Q(add_1104_n19) );
  INVX0 add_1104_U21 ( .ZN(add_1104_n21), .INP(n9911) );
  NOR2X0 add_1104_U22 ( .QN(N13), .IN1(add_1104_n22), .IN2(add_1104_n23) );
  INVX0 add_1104_U7 ( .ZN(add_1104_n7), .INP(n9903) );
  NOR2X0 add_1104_U8 ( .QN(N15), .IN1(add_1104_n8), .IN2(add_1104_n9) );
  AND2X1 add_1104_U9 ( .IN1(add_1104_n10), .IN2(add_1104_n11), .Q(add_1104_n9)
         );
  NOR2X0 add_1104_U10 ( .QN(add_1104_n8), .IN1(add_1104_n10), 
        .IN2(add_1104_n11) );
  NAND2X0 add_1104_U11 ( .IN1(add_1104_n12), .IN2(add_1104_n13), 
        .QN(add_1104_n11) );
  NAND2X0 add_1104_U12 ( .IN1(si_8_), .IN2(add_1104_n14), .QN(add_1104_n13) );
  OR2X1 add_1104_U13 ( .IN2(si_8_), .IN1(add_1104_n14), .Q(add_1104_n12) );
  INVX0 add_1104_U14 ( .ZN(add_1104_n14), .INP(n9907) );
  NOR2X0 add_1104_U1 ( .QN(N16), .IN1(add_1104_n1), .IN2(add_1104_n2) );
  AND2X1 add_1104_U2 ( .IN1(add_1104_n3), .IN2(add_1104_n4), .Q(add_1104_n2)
         );
  NOR2X0 add_1104_U3 ( .QN(add_1104_n1), .IN1(add_1104_n3), .IN2(add_1104_n4)
         );
  NAND2X0 add_1104_U4 ( .IN1(add_1104_n5), .IN2(add_1104_n6), .QN(add_1104_n4)
         );
  NAND2X0 add_1104_U5 ( .IN1(si_9_), .IN2(add_1104_n7), .QN(add_1104_n6) );
  OR2X1 add_1104_U6 ( .IN2(si_9_), .IN1(add_1104_n7), .Q(add_1104_n5) );
  NOR2X0 r794_U31 ( .QN(P1_N814), .IN1(r794_n28), .IN2(r794_n29) );
  OR2X1 r794_U30 ( .IN2(P1_N660), .IN1(r794_n27), .Q(r794_n26) );
  AND2X1 r794_U29 ( .IN1(r794_n26), .IN2(P1_N661), .Q(r794_n24) );
  NOR2X0 r794_U28 ( .QN(r794_n25), .IN1(P1_N661), .IN2(r794_n26) );
  NOR2X0 r794_U27 ( .QN(P1_N815), .IN1(r794_n24), .IN2(r794_n25) );
  AND2X1 r794_U26 ( .IN1(r794_n21), .IN2(P1_N633), .Q(r794_n22) );
  NOR2X0 r794_U25 ( .QN(r794_n23), .IN1(P1_N633), .IN2(r794_n21) );
  NOR2X0 r794_U24 ( .QN(P1_N787), .IN1(r794_n22), .IN2(r794_n23) );
  OR2X1 r794_U23 ( .IN2(P1_N633), .IN1(r794_n21), .Q(r794_n20) );
  AND2X1 r794_U22 ( .IN1(r794_n20), .IN2(P1_N634), .Q(r794_n18) );
  NOR2X0 r794_U21 ( .QN(r794_n19), .IN1(P1_N634), .IN2(r794_n20) );
  NOR2X0 r794_U20 ( .QN(P1_N788), .IN1(r794_n18), .IN2(r794_n19) );
  INVX0 r794_U19 ( .ZN(r794_n14), .INP(r794_n17) );
  AND2X1 r794_U18 ( .IN1(r794_n14), .IN2(P1_N635), .Q(r794_n15) );
  NOR2X0 r794_U17 ( .QN(r794_n16), .IN1(P1_N635), .IN2(r794_n14) );
  NOR2X0 r794_U16 ( .QN(P1_N789), .IN1(r794_n15), .IN2(r794_n16) );
  OR2X1 r794_U15 ( .IN2(P1_N635), .IN1(r794_n14), .Q(r794_n13) );
  AND2X1 r794_U14 ( .IN1(r794_n13), .IN2(P1_N636), .Q(r794_n11) );
  NOR2X0 r794_U13 ( .QN(r794_n12), .IN1(P1_N636), .IN2(r794_n13) );
  NOR2X0 r794_U12 ( .QN(P1_N790), .IN1(r794_n11), .IN2(r794_n12) );
  AND2X1 r794_U11 ( .IN1(r794_n8), .IN2(P1_N637), .Q(r794_n9) );
  NOR2X0 r794_U10 ( .QN(r794_n10), .IN1(P1_N637), .IN2(r794_n8) );
  NOR2X0 r794_U9 ( .QN(P1_N791), .IN1(r794_n9), .IN2(r794_n10) );
  OR2X1 r794_U8 ( .IN2(P1_N637), .IN1(r794_n8), .Q(r794_n7) );
  AND2X1 r794_U7 ( .IN1(r794_n7), .IN2(P1_N638), .Q(r794_n5) );
  NOR2X0 r794_U6 ( .QN(r794_n6), .IN1(P1_N638), .IN2(r794_n7) );
  NOR2X0 r794_U5 ( .QN(P1_N792), .IN1(r794_n5), .IN2(r794_n6) );
  AND2X1 r794_U4 ( .IN1(r794_n4), .IN2(P1_N639), .Q(r794_n2) );
  NOR2X0 r794_U3 ( .QN(r794_n3), .IN1(P1_N639), .IN2(r794_n4) );
  NOR2X0 r794_U2 ( .QN(P1_N793), .IN1(r794_n2), .IN2(r794_n3) );
  NOR2X0 r794_U124 ( .QN(P1_N796), .IN1(r794_n102), .IN2(r794_n103) );
  OR2X1 r794_U123 ( .IN2(P1_N641), .IN1(P1_N642), .Q(r794_n100) );
  NOR2X0 r794_U122 ( .QN(r794_n93), .IN1(r794_n100), .IN2(r794_n101) );
  INVX0 r794_U121 ( .ZN(r794_n97), .INP(r794_n93) );
  AND2X1 r794_U120 ( .IN1(r794_n97), .IN2(P1_N643), .Q(r794_n98) );
  NOR2X0 r794_U119 ( .QN(r794_n99), .IN1(P1_N643), .IN2(r794_n97) );
  NOR2X0 r794_U118 ( .QN(P1_N797), .IN1(r794_n98), .IN2(r794_n99) );
  OR2X1 r794_U117 ( .IN2(P1_N643), .IN1(r794_n97), .Q(r794_n96) );
  AND2X1 r794_U116 ( .IN1(r794_n96), .IN2(P1_N644), .Q(r794_n94) );
  NOR2X0 r794_U115 ( .QN(r794_n95), .IN1(P1_N644), .IN2(r794_n96) );
  NOR2X0 r794_U114 ( .QN(P1_N798), .IN1(r794_n94), .IN2(r794_n95) );
  NOR2X0 r794_U113 ( .QN(r794_n92), .IN1(P1_N644), .IN2(P1_N643) );
  NAND2X0 r794_U112 ( .IN1(r794_n92), .IN2(r794_n93), .QN(r794_n86) );
  AND2X1 r794_U111 ( .IN1(r794_n86), .IN2(P1_N645), .Q(r794_n90) );
  NOR2X0 r794_U110 ( .QN(r794_n91), .IN1(P1_N645), .IN2(r794_n86) );
  NOR2X0 r794_U109 ( .QN(P1_N799), .IN1(r794_n90), .IN2(r794_n91) );
  OR2X1 r794_U108 ( .IN2(P1_N645), .IN1(r794_n86), .Q(r794_n89) );
  AND2X1 r794_U107 ( .IN1(r794_n89), .IN2(P1_N646), .Q(r794_n87) );
  NOR2X0 r794_U106 ( .QN(r794_n88), .IN1(P1_N646), .IN2(r794_n89) );
  NOR2X0 r794_U105 ( .QN(P1_N800), .IN1(r794_n87), .IN2(r794_n88) );
  OR2X1 r794_U104 ( .IN2(P1_N645), .IN1(P1_N646), .Q(r794_n85) );
  NOR2X0 r794_U103 ( .QN(r794_n78), .IN1(r794_n85), .IN2(r794_n86) );
  INVX0 r794_U102 ( .ZN(r794_n82), .INP(r794_n78) );
  AND2X1 r794_U101 ( .IN1(r794_n82), .IN2(P1_N647), .Q(r794_n83) );
  NOR2X0 r794_U100 ( .QN(r794_n84), .IN1(P1_N647), .IN2(r794_n82) );
  NOR2X0 r794_U99 ( .QN(P1_N801), .IN1(r794_n83), .IN2(r794_n84) );
  OR2X1 r794_U98 ( .IN2(P1_N647), .IN1(r794_n82), .Q(r794_n81) );
  AND2X1 r794_U97 ( .IN1(r794_n81), .IN2(P1_N648), .Q(r794_n79) );
  NOR2X0 r794_U96 ( .QN(r794_n80), .IN1(P1_N648), .IN2(r794_n81) );
  NOR2X0 r794_U95 ( .QN(P1_N802), .IN1(r794_n79), .IN2(r794_n80) );
  NOR2X0 r794_U94 ( .QN(r794_n77), .IN1(P1_N648), .IN2(P1_N647) );
  NAND2X0 r794_U93 ( .IN1(r794_n77), .IN2(r794_n78), .QN(r794_n68) );
  AND2X1 r794_U92 ( .IN1(r794_n68), .IN2(P1_N649), .Q(r794_n75) );
  NOR2X0 r794_U91 ( .QN(r794_n76), .IN1(P1_N649), .IN2(r794_n68) );
  NOR2X0 r794_U90 ( .QN(P1_N803), .IN1(r794_n75), .IN2(r794_n76) );
  OR2X1 r794_U89 ( .IN2(P1_N631), .IN1(n7274), .Q(r794_n72) );
  NAND2X0 r794_U88 ( .IN1(P1_N631), .IN2(n7274), .QN(r794_n73) );
  NAND2X0 r794_U87 ( .IN1(r794_n72), .IN2(r794_n73), .QN(P1_N785) );
  OR2X1 r794_U86 ( .IN2(P1_N649), .IN1(r794_n68), .Q(r794_n71) );
  AND2X1 r794_U85 ( .IN1(r794_n71), .IN2(P1_N650), .Q(r794_n69) );
  NOR2X0 r794_U84 ( .QN(r794_n70), .IN1(P1_N650), .IN2(r794_n71) );
  NOR2X0 r794_U83 ( .QN(P1_N804), .IN1(r794_n69), .IN2(r794_n70) );
  OR2X1 r794_U82 ( .IN2(P1_N649), .IN1(P1_N650), .Q(r794_n67) );
  NOR2X0 r794_U81 ( .QN(r794_n60), .IN1(r794_n67), .IN2(r794_n68) );
  INVX0 r794_U80 ( .ZN(r794_n64), .INP(r794_n60) );
  AND2X1 r794_U79 ( .IN1(r794_n64), .IN2(P1_N651), .Q(r794_n65) );
  NOR2X0 r794_U78 ( .QN(r794_n66), .IN1(P1_N651), .IN2(r794_n64) );
  NOR2X0 r794_U77 ( .QN(P1_N805), .IN1(r794_n65), .IN2(r794_n66) );
  OR2X1 r794_U76 ( .IN2(P1_N651), .IN1(r794_n64), .Q(r794_n63) );
  AND2X1 r794_U75 ( .IN1(r794_n63), .IN2(P1_N652), .Q(r794_n61) );
  NOR2X0 r794_U74 ( .QN(r794_n62), .IN1(P1_N652), .IN2(r794_n63) );
  NOR2X0 r794_U73 ( .QN(P1_N806), .IN1(r794_n61), .IN2(r794_n62) );
  NOR2X0 r794_U72 ( .QN(r794_n59), .IN1(P1_N652), .IN2(P1_N651) );
  NAND2X0 r794_U71 ( .IN1(r794_n59), .IN2(r794_n60), .QN(r794_n53) );
  AND2X1 r794_U70 ( .IN1(r794_n53), .IN2(P1_N653), .Q(r794_n57) );
  NOR2X0 r794_U69 ( .QN(r794_n58), .IN1(P1_N653), .IN2(r794_n53) );
  NOR2X0 r794_U68 ( .QN(P1_N807), .IN1(r794_n57), .IN2(r794_n58) );
  OR2X1 r794_U67 ( .IN2(P1_N653), .IN1(r794_n53), .Q(r794_n56) );
  AND2X1 r794_U66 ( .IN1(r794_n56), .IN2(P1_N654), .Q(r794_n54) );
  NOR2X0 r794_U65 ( .QN(r794_n55), .IN1(P1_N654), .IN2(r794_n56) );
  NOR2X0 r794_U64 ( .QN(P1_N808), .IN1(r794_n54), .IN2(r794_n55) );
  OR2X1 r794_U63 ( .IN2(P1_N653), .IN1(P1_N654), .Q(r794_n52) );
  NOR2X0 r794_U62 ( .QN(r794_n45), .IN1(r794_n52), .IN2(r794_n53) );
  INVX0 r794_U61 ( .ZN(r794_n49), .INP(r794_n45) );
  AND2X1 r794_U60 ( .IN1(r794_n49), .IN2(P1_N655), .Q(r794_n50) );
  NOR2X0 r794_U59 ( .QN(r794_n51), .IN1(P1_N655), .IN2(r794_n49) );
  NOR2X0 r794_U58 ( .QN(P1_N809), .IN1(r794_n50), .IN2(r794_n51) );
  OR2X1 r794_U57 ( .IN2(P1_N655), .IN1(r794_n49), .Q(r794_n48) );
  AND2X1 r794_U56 ( .IN1(r794_n48), .IN2(P1_N656), .Q(r794_n46) );
  NOR2X0 r794_U55 ( .QN(r794_n47), .IN1(P1_N656), .IN2(r794_n48) );
  NOR2X0 r794_U54 ( .QN(P1_N810), .IN1(r794_n46), .IN2(r794_n47) );
  NOR2X0 r794_U53 ( .QN(r794_n44), .IN1(P1_N656), .IN2(P1_N655) );
  NAND2X0 r794_U52 ( .IN1(r794_n44), .IN2(r794_n45), .QN(r794_n38) );
  AND2X1 r794_U51 ( .IN1(r794_n38), .IN2(P1_N657), .Q(r794_n42) );
  NOR2X0 r794_U50 ( .QN(r794_n43), .IN1(P1_N657), .IN2(r794_n38) );
  NOR2X0 r794_U49 ( .QN(P1_N811), .IN1(r794_n42), .IN2(r794_n43) );
  OR2X1 r794_U48 ( .IN2(P1_N657), .IN1(r794_n38), .Q(r794_n41) );
  AND2X1 r794_U47 ( .IN1(r794_n41), .IN2(P1_N658), .Q(r794_n39) );
  NOR2X0 r794_U46 ( .QN(r794_n40), .IN1(P1_N658), .IN2(r794_n41) );
  NOR2X0 r794_U45 ( .QN(P1_N812), .IN1(r794_n39), .IN2(r794_n40) );
  NOR2X0 r794_U44 ( .QN(r794_n36), .IN1(P1_N658), .IN2(P1_N657) );
  INVX0 r794_U43 ( .ZN(r794_n37), .INP(r794_n38) );
  NAND2X0 r794_U42 ( .IN1(r794_n36), .IN2(r794_n37), .QN(r794_n30) );
  AND2X1 r794_U41 ( .IN1(r794_n30), .IN2(P1_N659), .Q(r794_n34) );
  NOR2X0 r794_U40 ( .QN(r794_n35), .IN1(P1_N659), .IN2(r794_n30) );
  NOR2X0 r794_U39 ( .QN(P1_N813), .IN1(r794_n34), .IN2(r794_n35) );
  OR2X1 r794_U38 ( .IN2(P1_N630), .IN1(P1_N631), .Q(r794_n33) );
  AND2X1 r794_U37 ( .IN1(r794_n33), .IN2(P1_N632), .Q(r794_n31) );
  NOR2X0 r794_U36 ( .QN(r794_n32), .IN1(P1_N632), .IN2(r794_n33) );
  NOR2X0 r794_U35 ( .QN(P1_N786), .IN1(r794_n31), .IN2(r794_n32) );
  OR2X1 r794_U34 ( .IN2(P1_N659), .IN1(r794_n30), .Q(r794_n27) );
  AND2X1 r794_U33 ( .IN1(r794_n27), .IN2(P1_N660), .Q(r794_n28) );
  NOR2X0 r794_U32 ( .QN(r794_n29), .IN1(P1_N660), .IN2(r794_n27) );
  OR2X1 r794_U146 ( .IN2(P1_N637), .IN1(P1_N638), .Q(r794_n112) );
  NOR2X0 r794_U145 ( .QN(r794_n113), .IN1(P1_N636), .IN2(P1_N635) );
  OR2X1 r794_U144 ( .IN2(P1_N633), .IN1(P1_N634), .Q(r794_n114) );
  NOR2X0 r794_U143 ( .QN(r794_n115), .IN1(P1_N632), .IN2(P1_N631) );
  NAND2X0 r794_U141 ( .IN1(r794_n115), .IN2(n7274), .QN(r794_n21) );
  NOR2X0 r794_U140 ( .QN(r794_n17), .IN1(r794_n114), .IN2(r794_n21) );
  NAND2X0 r794_U139 ( .IN1(r794_n113), .IN2(r794_n17), .QN(r794_n8) );
  NOR2X0 r794_U138 ( .QN(r794_n108), .IN1(r794_n112), .IN2(r794_n8) );
  INVX0 r794_U137 ( .ZN(r794_n4), .INP(r794_n108) );
  OR2X1 r794_U136 ( .IN2(P1_N639), .IN1(r794_n4), .Q(r794_n111) );
  AND2X1 r794_U135 ( .IN1(r794_n111), .IN2(P1_N640), .Q(r794_n109) );
  NOR2X0 r794_U134 ( .QN(r794_n110), .IN1(P1_N640), .IN2(r794_n111) );
  NOR2X0 r794_U133 ( .QN(P1_N794), .IN1(r794_n109), .IN2(r794_n110) );
  NOR2X0 r794_U132 ( .QN(r794_n107), .IN1(P1_N639), .IN2(P1_N640) );
  NAND2X0 r794_U131 ( .IN1(r794_n107), .IN2(r794_n108), .QN(r794_n101) );
  AND2X1 r794_U130 ( .IN1(r794_n101), .IN2(P1_N641), .Q(r794_n105) );
  NOR2X0 r794_U129 ( .QN(r794_n106), .IN1(P1_N641), .IN2(r794_n101) );
  NOR2X0 r794_U128 ( .QN(P1_N795), .IN1(r794_n105), .IN2(r794_n106) );
  OR2X1 r794_U127 ( .IN2(P1_N641), .IN1(r794_n101), .Q(r794_n104) );
  AND2X1 r794_U126 ( .IN1(r794_n104), .IN2(P1_N642), .Q(r794_n102) );
  NOR2X0 r794_U125 ( .QN(r794_n103), .IN1(P1_N642), .IN2(r794_n104) );
  NAND2X0 P1_add_122_U67 ( .IN1(P1_add_122_n58), .IN2(P1_add_122_n59), 
        .QN(P1_N384) );
  INVX0 P1_add_122_U66 ( .ZN(P1_add_122_n54), .INP(n9649) );
  OR2X1 P1_add_122_U65 ( .IN2(P1_add_122_n53), .IN1(P1_add_122_n54), 
        .Q(P1_add_122_n57) );
  OR2X1 P1_add_122_U64 ( .IN2(n9413), .IN1(P1_add_122_n57), .Q(P1_add_122_n55)
         );
  NAND2X0 P1_add_122_U63 ( .IN1(n9413), .IN2(P1_add_122_n57), 
        .QN(P1_add_122_n56) );
  NAND2X0 P1_add_122_U62 ( .IN1(P1_add_122_n55), .IN2(P1_add_122_n56), 
        .QN(P1_N385) );
  NOR2X0 P1_add_122_U61 ( .QN(P1_add_122_n52), .IN1(P1_add_122_n53), 
        .IN2(P1_add_122_n54) );
  NAND2X0 P1_add_122_U60 ( .IN1(P1_add_122_n52), .IN2(n9413), 
        .QN(P1_add_122_n45) );
  OR2X1 P1_add_122_U59 ( .IN2(n9645), .IN1(P1_add_122_n45), .Q(P1_add_122_n50)
         );
  NAND2X0 P1_add_122_U58 ( .IN1(n9645), .IN2(P1_add_122_n45), 
        .QN(P1_add_122_n51) );
  NAND2X0 P1_add_122_U57 ( .IN1(P1_add_122_n50), .IN2(P1_add_122_n51), 
        .QN(P1_N386) );
  INVX0 P1_add_122_U56 ( .ZN(P1_add_122_n46), .INP(n9645) );
  OR2X1 P1_add_122_U55 ( .IN2(P1_add_122_n45), .IN1(P1_add_122_n46), 
        .Q(P1_add_122_n49) );
  OR2X1 P1_add_122_U54 ( .IN2(n9409), .IN1(P1_add_122_n49), .Q(P1_add_122_n47)
         );
  NAND2X0 P1_add_122_U53 ( .IN1(n9409), .IN2(P1_add_122_n49), 
        .QN(P1_add_122_n48) );
  NAND2X0 P1_add_122_U52 ( .IN1(P1_add_122_n47), .IN2(P1_add_122_n48), 
        .QN(P1_N387) );
  NOR2X0 P1_add_122_U51 ( .QN(P1_add_122_n44), .IN1(P1_add_122_n45), 
        .IN2(P1_add_122_n46) );
  NAND2X0 P1_add_122_U50 ( .IN1(P1_add_122_n44), .IN2(n9409), 
        .QN(P1_add_122_n37) );
  OR2X1 P1_add_122_U49 ( .IN2(n9641), .IN1(P1_add_122_n37), .Q(P1_add_122_n42)
         );
  NAND2X0 P1_add_122_U48 ( .IN1(n9641), .IN2(P1_add_122_n37), 
        .QN(P1_add_122_n43) );
  NAND2X0 P1_add_122_U47 ( .IN1(P1_add_122_n42), .IN2(P1_add_122_n43), 
        .QN(P1_N388) );
  INVX0 P1_add_122_U46 ( .ZN(P1_add_122_n38), .INP(n9641) );
  OR2X1 P1_add_122_U45 ( .IN2(P1_add_122_n37), .IN1(P1_add_122_n38), 
        .Q(P1_add_122_n41) );
  OR2X1 P1_add_122_U44 ( .IN2(n9405), .IN1(P1_add_122_n41), .Q(P1_add_122_n39)
         );
  NAND2X0 P1_add_122_U43 ( .IN1(n9405), .IN2(P1_add_122_n41), 
        .QN(P1_add_122_n40) );
  NAND2X0 P1_add_122_U42 ( .IN1(P1_add_122_n39), .IN2(P1_add_122_n40), 
        .QN(P1_N389) );
  NOR2X0 P1_add_122_U41 ( .QN(P1_add_122_n36), .IN1(P1_add_122_n37), 
        .IN2(P1_add_122_n38) );
  NAND2X0 P1_add_122_U40 ( .IN1(P1_add_122_n36), .IN2(n9405), 
        .QN(P1_add_122_n29) );
  OR2X1 P1_add_122_U39 ( .IN2(n9637), .IN1(P1_add_122_n29), .Q(P1_add_122_n34)
         );
  NAND2X0 P1_add_122_U38 ( .IN1(n9637), .IN2(P1_add_122_n29), 
        .QN(P1_add_122_n35) );
  NAND2X0 P1_add_122_U37 ( .IN1(P1_add_122_n34), .IN2(P1_add_122_n35), 
        .QN(P1_N390) );
  INVX0 P1_add_122_U36 ( .ZN(P1_add_122_n30), .INP(n9637) );
  OR2X1 P1_add_122_U35 ( .IN2(P1_add_122_n29), .IN1(P1_add_122_n30), 
        .Q(P1_add_122_n33) );
  OR2X1 P1_add_122_U34 ( .IN2(n9401), .IN1(P1_add_122_n33), .Q(P1_add_122_n31)
         );
  NAND2X0 P1_add_122_U33 ( .IN1(n9401), .IN2(P1_add_122_n33), 
        .QN(P1_add_122_n32) );
  NAND2X0 P1_add_122_U32 ( .IN1(P1_add_122_n31), .IN2(P1_add_122_n32), 
        .QN(P1_N391) );
  NOR2X0 P1_add_122_U31 ( .QN(P1_add_122_n28), .IN1(P1_add_122_n29), 
        .IN2(P1_add_122_n30) );
  NAND2X0 P1_add_122_U30 ( .IN1(P1_add_122_n28), .IN2(n9401), 
        .QN(P1_add_122_n24) );
  OR2X1 P1_add_122_U29 ( .IN2(n9633), .IN1(P1_add_122_n24), .Q(P1_add_122_n26)
         );
  NAND2X0 P1_add_122_U28 ( .IN1(n9633), .IN2(P1_add_122_n24), 
        .QN(P1_add_122_n27) );
  NAND2X0 P1_add_122_U27 ( .IN1(P1_add_122_n26), .IN2(P1_add_122_n27), 
        .QN(P1_N392) );
  INVX0 P1_add_122_U26 ( .ZN(P1_add_122_n25), .INP(n9633) );
  NOR2X0 P1_add_122_U25 ( .QN(P1_N393), .IN1(P1_add_122_n24), 
        .IN2(P1_add_122_n25) );
  NAND2X0 P1_add_122_U24 ( .IN1(n6594), .IN2(P1_add_122_n23), 
        .QN(P1_add_122_n21) );
  NAND2X0 P1_add_122_U23 ( .IN1(n9657), .IN2(n18451), .QN(P1_add_122_n22) );
  NAND2X0 P1_add_122_U22 ( .IN1(P1_add_122_n21), .IN2(P1_add_122_n22), 
        .QN(P1_N368) );
  NAND2X0 P1_add_122_U21 ( .IN1(n9657), .IN2(n6594), .QN(P1_add_122_n20) );
  OR2X1 P1_add_122_U20 ( .IN2(n9689), .IN1(P1_add_122_n20), .Q(P1_add_122_n18)
         );
  NAND2X0 P1_add_122_U19 ( .IN1(n9689), .IN2(P1_add_122_n20), 
        .QN(P1_add_122_n19) );
  NAND2X0 P1_add_122_U18 ( .IN1(P1_add_122_n18), .IN2(P1_add_122_n19), 
        .QN(P1_N369) );
  OR2X1 P1_add_122_U17 ( .IN2(n10015), .IN1(P1_add_122_n15), 
        .Q(P1_add_122_n16) );
  NAND2X0 P1_add_122_U16 ( .IN1(n10015), .IN2(P1_add_122_n15), 
        .QN(P1_add_122_n17) );
  NAND2X0 P1_add_122_U15 ( .IN1(P1_add_122_n16), .IN2(P1_add_122_n17), 
        .QN(P1_N370) );
  OR2X1 P1_add_122_U14 ( .IN2(P1_add_122_n15), .IN1(P1_add_122_n14), 
        .Q(P1_add_122_n13) );
  OR2X1 P1_add_122_U13 ( .IN2(n9685), .IN1(P1_add_122_n13), .Q(P1_add_122_n11)
         );
  NAND2X0 P1_add_122_U12 ( .IN1(n9685), .IN2(P1_add_122_n13), 
        .QN(P1_add_122_n12) );
  NAND2X0 P1_add_122_U11 ( .IN1(P1_add_122_n11), .IN2(P1_add_122_n12), 
        .QN(P1_N371) );
  OR2X1 P1_add_122_U10 ( .IN2(n10011), .IN1(P1_add_122_n8), .Q(P1_add_122_n9)
         );
  NAND2X0 P1_add_122_U9 ( .IN1(n10011), .IN2(P1_add_122_n8), 
        .QN(P1_add_122_n10) );
  NAND2X0 P1_add_122_U8 ( .IN1(P1_add_122_n9), .IN2(P1_add_122_n10), 
        .QN(P1_N372) );
  OR2X1 P1_add_122_U7 ( .IN2(P1_add_122_n8), .IN1(P1_add_122_n7), 
        .Q(P1_add_122_n6) );
  OR2X1 P1_add_122_U6 ( .IN2(n9681), .IN1(P1_add_122_n6), .Q(P1_add_122_n4) );
  NAND2X0 P1_add_122_U5 ( .IN1(n9681), .IN2(P1_add_122_n6), .QN(P1_add_122_n5)
         );
  INVX0 P1_add_122_U128 ( .ZN(P1_add_122_n23), .INP(n9657) );
  NOR2X0 P1_add_122_U127 ( .QN(P1_add_122_n102), .IN1(n18451), 
        .IN2(P1_add_122_n23) );
  NAND2X0 P1_add_122_U126 ( .IN1(P1_add_122_n102), .IN2(n9689), 
        .QN(P1_add_122_n15) );
  INVX0 P1_add_122_U125 ( .ZN(P1_add_122_n14), .INP(n10015) );
  NOR2X0 P1_add_122_U124 ( .QN(P1_add_122_n101), .IN1(P1_add_122_n15), 
        .IN2(P1_add_122_n14) );
  NAND2X0 P1_add_122_U123 ( .IN1(P1_add_122_n101), .IN2(n9685), 
        .QN(P1_add_122_n8) );
  INVX0 P1_add_122_U122 ( .ZN(P1_add_122_n7), .INP(n10011) );
  NOR2X0 P1_add_122_U121 ( .QN(P1_add_122_n100), .IN1(P1_add_122_n8), 
        .IN2(P1_add_122_n7) );
  NAND2X0 P1_add_122_U120 ( .IN1(P1_add_122_n100), .IN2(n9681), 
        .QN(P1_add_122_n93) );
  OR2X1 P1_add_122_U119 ( .IN2(n9867), .IN1(P1_add_122_n93), 
        .Q(P1_add_122_n98) );
  NAND2X0 P1_add_122_U118 ( .IN1(n9867), .IN2(P1_add_122_n93), 
        .QN(P1_add_122_n99) );
  NAND2X0 P1_add_122_U117 ( .IN1(P1_add_122_n98), .IN2(P1_add_122_n99), 
        .QN(P1_N374) );
  INVX0 P1_add_122_U116 ( .ZN(P1_add_122_n94), .INP(n9867) );
  OR2X1 P1_add_122_U115 ( .IN2(P1_add_122_n93), .IN1(P1_add_122_n94), 
        .Q(P1_add_122_n97) );
  OR2X1 P1_add_122_U114 ( .IN2(n9677), .IN1(P1_add_122_n97), 
        .Q(P1_add_122_n95) );
  NAND2X0 P1_add_122_U113 ( .IN1(n9677), .IN2(P1_add_122_n97), 
        .QN(P1_add_122_n96) );
  NAND2X0 P1_add_122_U112 ( .IN1(P1_add_122_n95), .IN2(P1_add_122_n96), 
        .QN(P1_N375) );
  NOR2X0 P1_add_122_U111 ( .QN(P1_add_122_n92), .IN1(P1_add_122_n93), 
        .IN2(P1_add_122_n94) );
  NAND2X0 P1_add_122_U110 ( .IN1(P1_add_122_n92), .IN2(n9677), 
        .QN(P1_add_122_n85) );
  OR2X1 P1_add_122_U109 ( .IN2(n9863), .IN1(P1_add_122_n85), 
        .Q(P1_add_122_n90) );
  NAND2X0 P1_add_122_U108 ( .IN1(n9863), .IN2(P1_add_122_n85), 
        .QN(P1_add_122_n91) );
  NAND2X0 P1_add_122_U107 ( .IN1(P1_add_122_n90), .IN2(P1_add_122_n91), 
        .QN(P1_N376) );
  INVX0 P1_add_122_U106 ( .ZN(P1_add_122_n86), .INP(n9863) );
  OR2X1 P1_add_122_U105 ( .IN2(P1_add_122_n85), .IN1(P1_add_122_n86), 
        .Q(P1_add_122_n89) );
  OR2X1 P1_add_122_U104 ( .IN2(n9673), .IN1(P1_add_122_n89), 
        .Q(P1_add_122_n87) );
  NAND2X0 P1_add_122_U103 ( .IN1(n9673), .IN2(P1_add_122_n89), 
        .QN(P1_add_122_n88) );
  NAND2X0 P1_add_122_U102 ( .IN1(P1_add_122_n87), .IN2(P1_add_122_n88), 
        .QN(P1_N377) );
  NOR2X0 P1_add_122_U101 ( .QN(P1_add_122_n84), .IN1(P1_add_122_n85), 
        .IN2(P1_add_122_n86) );
  NAND2X0 P1_add_122_U100 ( .IN1(P1_add_122_n84), .IN2(n9673), 
        .QN(P1_add_122_n77) );
  OR2X1 P1_add_122_U99 ( .IN2(n9859), .IN1(P1_add_122_n77), .Q(P1_add_122_n82)
         );
  NAND2X0 P1_add_122_U98 ( .IN1(n9859), .IN2(P1_add_122_n77), 
        .QN(P1_add_122_n83) );
  NAND2X0 P1_add_122_U97 ( .IN1(P1_add_122_n82), .IN2(P1_add_122_n83), 
        .QN(P1_N378) );
  INVX0 P1_add_122_U96 ( .ZN(P1_add_122_n78), .INP(n9859) );
  OR2X1 P1_add_122_U95 ( .IN2(P1_add_122_n77), .IN1(P1_add_122_n78), 
        .Q(P1_add_122_n81) );
  OR2X1 P1_add_122_U94 ( .IN2(n9669), .IN1(P1_add_122_n81), .Q(P1_add_122_n79)
         );
  NAND2X0 P1_add_122_U93 ( .IN1(n9669), .IN2(P1_add_122_n81), 
        .QN(P1_add_122_n80) );
  NAND2X0 P1_add_122_U92 ( .IN1(P1_add_122_n79), .IN2(P1_add_122_n80), 
        .QN(P1_N379) );
  NOR2X0 P1_add_122_U91 ( .QN(P1_add_122_n76), .IN1(P1_add_122_n77), 
        .IN2(P1_add_122_n78) );
  NAND2X0 P1_add_122_U90 ( .IN1(P1_add_122_n76), .IN2(n9669), 
        .QN(P1_add_122_n69) );
  OR2X1 P1_add_122_U89 ( .IN2(n9855), .IN1(P1_add_122_n69), .Q(P1_add_122_n74)
         );
  NAND2X0 P1_add_122_U88 ( .IN1(n9855), .IN2(P1_add_122_n69), 
        .QN(P1_add_122_n75) );
  NAND2X0 P1_add_122_U87 ( .IN1(P1_add_122_n74), .IN2(P1_add_122_n75), 
        .QN(P1_N380) );
  INVX0 P1_add_122_U86 ( .ZN(P1_add_122_n70), .INP(n9855) );
  OR2X1 P1_add_122_U85 ( .IN2(P1_add_122_n69), .IN1(P1_add_122_n70), 
        .Q(P1_add_122_n73) );
  OR2X1 P1_add_122_U84 ( .IN2(n9665), .IN1(P1_add_122_n73), .Q(P1_add_122_n71)
         );
  NAND2X0 P1_add_122_U83 ( .IN1(n9665), .IN2(P1_add_122_n73), 
        .QN(P1_add_122_n72) );
  NAND2X0 P1_add_122_U82 ( .IN1(P1_add_122_n71), .IN2(P1_add_122_n72), 
        .QN(P1_N381) );
  NOR2X0 P1_add_122_U81 ( .QN(P1_add_122_n68), .IN1(P1_add_122_n69), 
        .IN2(P1_add_122_n70) );
  NAND2X0 P1_add_122_U80 ( .IN1(P1_add_122_n68), .IN2(n9665), 
        .QN(P1_add_122_n61) );
  OR2X1 P1_add_122_U79 ( .IN2(n9851), .IN1(P1_add_122_n61), .Q(P1_add_122_n66)
         );
  NAND2X0 P1_add_122_U78 ( .IN1(n9851), .IN2(P1_add_122_n61), 
        .QN(P1_add_122_n67) );
  NAND2X0 P1_add_122_U77 ( .IN1(P1_add_122_n66), .IN2(P1_add_122_n67), 
        .QN(P1_N382) );
  INVX0 P1_add_122_U76 ( .ZN(P1_add_122_n62), .INP(n9851) );
  OR2X1 P1_add_122_U75 ( .IN2(P1_add_122_n61), .IN1(P1_add_122_n62), 
        .Q(P1_add_122_n65) );
  OR2X1 P1_add_122_U74 ( .IN2(n9661), .IN1(P1_add_122_n65), .Q(P1_add_122_n63)
         );
  NAND2X0 P1_add_122_U73 ( .IN1(n9661), .IN2(P1_add_122_n65), 
        .QN(P1_add_122_n64) );
  NAND2X0 P1_add_122_U72 ( .IN1(P1_add_122_n63), .IN2(P1_add_122_n64), 
        .QN(P1_N383) );
  NOR2X0 P1_add_122_U71 ( .QN(P1_add_122_n60), .IN1(P1_add_122_n61), 
        .IN2(P1_add_122_n62) );
  NAND2X0 P1_add_122_U70 ( .IN1(P1_add_122_n60), .IN2(n9661), 
        .QN(P1_add_122_n53) );
  OR2X1 P1_add_122_U69 ( .IN2(n9649), .IN1(P1_add_122_n53), .Q(P1_add_122_n58)
         );
  NAND2X0 P1_add_122_U68 ( .IN1(n9649), .IN2(P1_add_122_n53), 
        .QN(P1_add_122_n59) );
  NAND2X1 P1_add_122_U4 ( .IN1(P1_add_122_n4), .IN2(P1_add_122_n5), 
        .QN(P1_N373) );
  NOR2X0 r796_U15 ( .QN(P1_N1771), .IN1(r796_n15), .IN2(r796_n16) );
  OR2X1 r796_U13 ( .IN2(P1_N1620), .IN1(n7073), .Q(r796_n12) );
  NAND2X0 r796_U12 ( .IN1(P1_N1620), .IN2(n7073), .QN(r796_n13) );
  NAND2X0 r796_U11 ( .IN1(r796_n12), .IN2(r796_n13), .QN(r796_n11) );
  NOR2X0 r796_U10 ( .QN(r796_n8), .IN1(r796_n10), .IN2(r796_n11) );
  AND2X1 r796_U9 ( .IN1(r796_n10), .IN2(r796_n11), .Q(r796_n9) );
  NOR2X0 r796_U8 ( .QN(P1_N1772), .IN1(r796_n8), .IN2(r796_n9) );
  OR2X1 r796_U6 ( .IN2(P1_N1621), .IN1(n7071), .Q(r796_n5) );
  NAND2X0 r796_U5 ( .IN1(P1_N1621), .IN2(n7071), .QN(r796_n6) );
  NAND2X0 r796_U4 ( .IN1(r796_n5), .IN2(r796_n6), .QN(r796_n4) );
  NOR2X0 r796_U3 ( .QN(r796_n1), .IN1(r796_n3), .IN2(r796_n4) );
  AND2X1 r796_U2 ( .IN1(r796_n3), .IN2(r796_n4), .Q(r796_n2) );
  NOR2X0 r796_U1 ( .QN(P1_N1773), .IN1(r796_n1), .IN2(r796_n2) );
  NAND2X0 r796_U108 ( .IN1(r796_n104), .IN2(r796_n105), .QN(r796_n97) );
  OR2X1 r796_U106 ( .IN2(P1_N1637), .IN1(n7130), .Q(r796_n101) );
  NAND2X0 r796_U105 ( .IN1(P1_N1637), .IN2(n7130), .QN(r796_n102) );
  NAND2X0 r796_U104 ( .IN1(r796_n101), .IN2(r796_n102), .QN(r796_n100) );
  NOR2X0 r796_U103 ( .QN(r796_n98), .IN1(r796_n97), .IN2(r796_n100) );
  AND2X1 r796_U102 ( .IN1(r796_n97), .IN2(r796_n100), .Q(r796_n99) );
  NOR2X0 r796_U101 ( .QN(P1_N1789), .IN1(r796_n98), .IN2(r796_n99) );
  NAND2X0 r796_U100 ( .IN1(n7129), .IN2(r796_n97), .QN(r796_n94) );
  OR2X1 r796_U99 ( .IN2(n7129), .IN1(r796_n97), .Q(r796_n96) );
  NAND2X0 r796_U98 ( .IN1(P1_N1637), .IN2(r796_n96), .QN(r796_n95) );
  NAND2X0 r796_U97 ( .IN1(r796_n94), .IN2(r796_n95), .QN(r796_n87) );
  OR2X1 r796_U95 ( .IN2(P1_N1638), .IN1(n7125), .Q(r796_n91) );
  NAND2X0 r796_U94 ( .IN1(P1_N1638), .IN2(n7125), .QN(r796_n92) );
  NAND2X0 r796_U93 ( .IN1(r796_n91), .IN2(r796_n92), .QN(r796_n90) );
  NOR2X0 r796_U92 ( .QN(r796_n88), .IN1(r796_n87), .IN2(r796_n90) );
  AND2X1 r796_U91 ( .IN1(r796_n87), .IN2(r796_n90), .Q(r796_n89) );
  NOR2X0 r796_U90 ( .QN(P1_N1790), .IN1(r796_n88), .IN2(r796_n89) );
  NAND2X0 r796_U89 ( .IN1(n7124), .IN2(r796_n87), .QN(r796_n84) );
  OR2X1 r796_U88 ( .IN2(n7124), .IN1(r796_n87), .Q(r796_n86) );
  NAND2X0 r796_U87 ( .IN1(P1_N1638), .IN2(r796_n86), .QN(r796_n85) );
  NAND2X0 r796_U86 ( .IN1(r796_n84), .IN2(r796_n85), .QN(r796_n77) );
  OR2X1 r796_U84 ( .IN2(P1_N1639), .IN1(n7119), .Q(r796_n81) );
  NAND2X0 r796_U83 ( .IN1(P1_N1639), .IN2(n7119), .QN(r796_n82) );
  NAND2X0 r796_U82 ( .IN1(r796_n81), .IN2(r796_n82), .QN(r796_n80) );
  NOR2X0 r796_U81 ( .QN(r796_n78), .IN1(r796_n77), .IN2(r796_n80) );
  AND2X1 r796_U80 ( .IN1(r796_n77), .IN2(r796_n80), .Q(r796_n79) );
  NOR2X0 r796_U79 ( .QN(P1_N1791), .IN1(r796_n78), .IN2(r796_n79) );
  NAND2X0 r796_U78 ( .IN1(P1_N5176), .IN2(r796_n77), .QN(r796_n74) );
  OR2X1 r796_U77 ( .IN2(P1_N5176), .IN1(r796_n77), .Q(r796_n76) );
  NAND2X0 r796_U76 ( .IN1(P1_N1639), .IN2(r796_n76), .QN(r796_n75) );
  NAND2X0 r796_U75 ( .IN1(r796_n74), .IN2(r796_n75), .QN(r796_n64) );
  OR2X1 r796_U73 ( .IN2(P1_N1640), .IN1(n7117), .Q(r796_n71) );
  NAND2X0 r796_U72 ( .IN1(P1_N1640), .IN2(n7117), .QN(r796_n72) );
  NAND2X0 r796_U71 ( .IN1(r796_n71), .IN2(r796_n72), .QN(r796_n70) );
  NOR2X0 r796_U70 ( .QN(r796_n68), .IN1(r796_n64), .IN2(r796_n70) );
  AND2X1 r796_U69 ( .IN1(r796_n64), .IN2(r796_n70), .Q(r796_n69) );
  NOR2X0 r796_U68 ( .QN(P1_N1792), .IN1(r796_n68), .IN2(r796_n69) );
  OR2X1 r796_U66 ( .IN2(P1_N1641), .IN1(n7146), .Q(r796_n65) );
  NAND2X0 r796_U65 ( .IN1(P1_N1641), .IN2(n7146), .QN(r796_n66) );
  NAND2X0 r796_U64 ( .IN1(r796_n65), .IN2(r796_n66), .QN(r796_n60) );
  NAND2X0 r796_U63 ( .IN1(P1_N5177), .IN2(r796_n64), .QN(r796_n61) );
  OR2X1 r796_U62 ( .IN2(P1_N5177), .IN1(r796_n64), .Q(r796_n63) );
  NAND2X0 r796_U61 ( .IN1(P1_N1640), .IN2(r796_n63), .QN(r796_n62) );
  NAND2X0 r796_U60 ( .IN1(r796_n61), .IN2(r796_n62), .QN(r796_n59) );
  NOR2X0 r796_U59 ( .QN(r796_n57), .IN1(r796_n60), .IN2(r796_n59) );
  AND2X1 r796_U58 ( .IN1(r796_n59), .IN2(r796_n60), .Q(r796_n58) );
  NOR2X0 r796_U57 ( .QN(P1_N1793), .IN1(r796_n57), .IN2(r796_n58) );
  OR2X1 r796_U55 ( .IN2(P1_N1614), .IN1(n7045), .Q(r796_n54) );
  NAND2X0 r796_U54 ( .IN1(P1_N1614), .IN2(n7045), .QN(r796_n55) );
  NAND2X0 r796_U53 ( .IN1(r796_n54), .IN2(r796_n55), .QN(r796_n53) );
  NOR2X0 r796_U52 ( .QN(r796_n50), .IN1(r796_n52), .IN2(r796_n53) );
  AND2X1 r796_U51 ( .IN1(r796_n52), .IN2(r796_n53), .Q(r796_n51) );
  NOR2X0 r796_U50 ( .QN(P1_N1766), .IN1(r796_n50), .IN2(r796_n51) );
  OR2X1 r796_U48 ( .IN2(P1_N1615), .IN1(n7043), .Q(r796_n47) );
  NAND2X0 r796_U47 ( .IN1(P1_N1615), .IN2(n7043), .QN(r796_n48) );
  NAND2X0 r796_U46 ( .IN1(r796_n47), .IN2(r796_n48), .QN(r796_n46) );
  NOR2X0 r796_U45 ( .QN(r796_n43), .IN1(r796_n45), .IN2(r796_n46) );
  AND2X1 r796_U44 ( .IN1(r796_n45), .IN2(r796_n46), .Q(r796_n44) );
  NOR2X0 r796_U43 ( .QN(P1_N1767), .IN1(r796_n43), .IN2(r796_n44) );
  OR2X1 r796_U41 ( .IN2(P1_N1616), .IN1(n7037), .Q(r796_n40) );
  NAND2X0 r796_U40 ( .IN1(P1_N1616), .IN2(n7037), .QN(r796_n41) );
  NAND2X0 r796_U39 ( .IN1(r796_n40), .IN2(r796_n41), .QN(r796_n39) );
  NOR2X0 r796_U38 ( .QN(r796_n36), .IN1(r796_n38), .IN2(r796_n39) );
  AND2X1 r796_U37 ( .IN1(r796_n38), .IN2(r796_n39), .Q(r796_n37) );
  NOR2X0 r796_U36 ( .QN(P1_N1768), .IN1(r796_n36), .IN2(r796_n37) );
  OR2X1 r796_U34 ( .IN2(P1_N1617), .IN1(n7082), .Q(r796_n33) );
  NAND2X0 r796_U33 ( .IN1(P1_N1617), .IN2(n7082), .QN(r796_n34) );
  NAND2X0 r796_U32 ( .IN1(r796_n33), .IN2(r796_n34), .QN(r796_n32) );
  NOR2X0 r796_U31 ( .QN(r796_n29), .IN1(r796_n31), .IN2(r796_n32) );
  AND2X1 r796_U30 ( .IN1(r796_n31), .IN2(r796_n32), .Q(r796_n30) );
  NOR2X0 r796_U29 ( .QN(P1_N1769), .IN1(r796_n29), .IN2(r796_n30) );
  OR2X1 r796_U27 ( .IN2(P1_N1618), .IN1(n7079), .Q(r796_n26) );
  NAND2X0 r796_U26 ( .IN1(P1_N1618), .IN2(n7079), .QN(r796_n27) );
  NAND2X0 r796_U25 ( .IN1(r796_n26), .IN2(r796_n27), .QN(r796_n25) );
  NOR2X0 r796_U24 ( .QN(r796_n22), .IN1(r796_n24), .IN2(r796_n25) );
  AND2X1 r796_U23 ( .IN1(r796_n24), .IN2(r796_n25), .Q(r796_n23) );
  NOR2X0 r796_U22 ( .QN(P1_N1770), .IN1(r796_n22), .IN2(r796_n23) );
  OR2X1 r796_U20 ( .IN2(P1_N1619), .IN1(n7076), .Q(r796_n19) );
  NAND2X0 r796_U19 ( .IN1(P1_N1619), .IN2(n7076), .QN(r796_n20) );
  NAND2X0 r796_U18 ( .IN1(r796_n19), .IN2(r796_n20), .QN(r796_n18) );
  NOR2X0 r796_U17 ( .QN(r796_n15), .IN1(r796_n17), .IN2(r796_n18) );
  AND2X1 r796_U16 ( .IN1(r796_n17), .IN2(r796_n18), .Q(r796_n16) );
  OR2X1 r796_U200 ( .IN2(P1_N1629), .IN1(n7105), .Q(r796_n188) );
  NAND2X0 r796_U199 ( .IN1(P1_N1629), .IN2(n7105), .QN(r796_n189) );
  NAND2X0 r796_U198 ( .IN1(r796_n188), .IN2(r796_n189), .QN(r796_n187) );
  NOR2X0 r796_U197 ( .QN(r796_n185), .IN1(r796_n184), .IN2(r796_n187) );
  AND2X1 r796_U196 ( .IN1(r796_n184), .IN2(r796_n187), .Q(r796_n186) );
  NOR2X0 r796_U195 ( .QN(P1_N1781), .IN1(r796_n185), .IN2(r796_n186) );
  NAND2X0 r796_U194 ( .IN1(n7106), .IN2(r796_n184), .QN(r796_n181) );
  OR2X1 r796_U193 ( .IN2(n7106), .IN1(r796_n184), .Q(r796_n183) );
  NAND2X0 r796_U192 ( .IN1(P1_N1629), .IN2(r796_n183), .QN(r796_n182) );
  NAND2X0 r796_U191 ( .IN1(r796_n181), .IN2(r796_n182), .QN(r796_n174) );
  OR2X1 r796_U189 ( .IN2(P1_N1630), .IN1(n7102), .Q(r796_n178) );
  NAND2X0 r796_U188 ( .IN1(P1_N1630), .IN2(n7102), .QN(r796_n179) );
  NAND2X0 r796_U187 ( .IN1(r796_n178), .IN2(r796_n179), .QN(r796_n177) );
  NOR2X0 r796_U186 ( .QN(r796_n175), .IN1(r796_n174), .IN2(r796_n177) );
  AND2X1 r796_U185 ( .IN1(r796_n174), .IN2(r796_n177), .Q(r796_n176) );
  NOR2X0 r796_U184 ( .QN(P1_N1782), .IN1(r796_n175), .IN2(r796_n176) );
  NAND2X0 r796_U183 ( .IN1(P1_N5167), .IN2(r796_n174), .QN(r796_n171) );
  OR2X1 r796_U182 ( .IN2(P1_N5167), .IN1(r796_n174), .Q(r796_n173) );
  NAND2X0 r796_U181 ( .IN1(P1_N1630), .IN2(r796_n173), .QN(r796_n172) );
  NAND2X0 r796_U180 ( .IN1(r796_n171), .IN2(r796_n172), .QN(r796_n157) );
  OR2X1 r796_U178 ( .IN2(P1_N1631), .IN1(n7098), .Q(r796_n168) );
  NAND2X0 r796_U177 ( .IN1(P1_N1631), .IN2(n7098), .QN(r796_n169) );
  NAND2X0 r796_U176 ( .IN1(r796_n168), .IN2(r796_n169), .QN(r796_n167) );
  NOR2X0 r796_U175 ( .QN(r796_n165), .IN1(r796_n157), .IN2(r796_n167) );
  AND2X1 r796_U174 ( .IN1(r796_n157), .IN2(r796_n167), .Q(r796_n166) );
  NOR2X0 r796_U173 ( .QN(P1_N1783), .IN1(r796_n165), .IN2(r796_n166) );
  OR2X1 r796_U172 ( .IN2(P1_N1613), .IN1(n7051), .Q(r796_n162) );
  NAND2X0 r796_U171 ( .IN1(P1_N1613), .IN2(n7051), .QN(r796_n163) );
  NAND2X0 r796_U170 ( .IN1(r796_n162), .IN2(r796_n163), .QN(r796_n160) );
  NAND2X0 r796_U169 ( .IN1(r796_n160), .IN2(r796_n161), .QN(r796_n158) );
  OR2X1 r796_U168 ( .IN2(r796_n161), .IN1(r796_n160), .Q(r796_n159) );
  NAND2X0 r796_U167 ( .IN1(r796_n158), .IN2(r796_n159), .QN(P1_N1765) );
  NAND2X0 r796_U166 ( .IN1(n7099), .IN2(r796_n157), .QN(r796_n154) );
  OR2X1 r796_U165 ( .IN2(n7099), .IN1(r796_n157), .Q(r796_n156) );
  NAND2X0 r796_U164 ( .IN1(P1_N1631), .IN2(r796_n156), .QN(r796_n155) );
  NAND2X0 r796_U163 ( .IN1(r796_n154), .IN2(r796_n155), .QN(r796_n147) );
  OR2X1 r796_U161 ( .IN2(P1_N1632), .IN1(n7095), .Q(r796_n151) );
  NAND2X0 r796_U160 ( .IN1(P1_N1632), .IN2(n7095), .QN(r796_n152) );
  NAND2X0 r796_U159 ( .IN1(r796_n151), .IN2(r796_n152), .QN(r796_n150) );
  NOR2X0 r796_U158 ( .QN(r796_n148), .IN1(r796_n147), .IN2(r796_n150) );
  AND2X1 r796_U157 ( .IN1(r796_n147), .IN2(r796_n150), .Q(r796_n149) );
  NOR2X0 r796_U156 ( .QN(P1_N1784), .IN1(r796_n148), .IN2(r796_n149) );
  NAND2X0 r796_U155 ( .IN1(P1_N5169), .IN2(r796_n147), .QN(r796_n144) );
  OR2X1 r796_U154 ( .IN2(P1_N5169), .IN1(r796_n147), .Q(r796_n146) );
  NAND2X0 r796_U153 ( .IN1(P1_N1632), .IN2(r796_n146), .QN(r796_n145) );
  NAND2X0 r796_U152 ( .IN1(r796_n144), .IN2(r796_n145), .QN(r796_n137) );
  OR2X1 r796_U150 ( .IN2(P1_N1633), .IN1(n7092), .Q(r796_n141) );
  NAND2X0 r796_U149 ( .IN1(P1_N1633), .IN2(n7092), .QN(r796_n142) );
  NAND2X0 r796_U148 ( .IN1(r796_n141), .IN2(r796_n142), .QN(r796_n140) );
  NOR2X0 r796_U147 ( .QN(r796_n138), .IN1(r796_n137), .IN2(r796_n140) );
  AND2X1 r796_U146 ( .IN1(r796_n137), .IN2(r796_n140), .Q(r796_n139) );
  NOR2X0 r796_U145 ( .QN(P1_N1785), .IN1(r796_n138), .IN2(r796_n139) );
  NAND2X0 r796_U144 ( .IN1(P1_N5170), .IN2(r796_n137), .QN(r796_n134) );
  OR2X1 r796_U143 ( .IN2(P1_N5170), .IN1(r796_n137), .Q(r796_n136) );
  NAND2X0 r796_U142 ( .IN1(P1_N1633), .IN2(r796_n136), .QN(r796_n135) );
  NAND2X0 r796_U141 ( .IN1(r796_n134), .IN2(r796_n135), .QN(r796_n127) );
  OR2X1 r796_U139 ( .IN2(P1_N1634), .IN1(n7090), .Q(r796_n131) );
  NAND2X0 r796_U138 ( .IN1(P1_N1634), .IN2(n7090), .QN(r796_n132) );
  NAND2X0 r796_U137 ( .IN1(r796_n131), .IN2(r796_n132), .QN(r796_n130) );
  NOR2X0 r796_U136 ( .QN(r796_n128), .IN1(r796_n127), .IN2(r796_n130) );
  AND2X1 r796_U135 ( .IN1(r796_n127), .IN2(r796_n130), .Q(r796_n129) );
  NOR2X0 r796_U134 ( .QN(P1_N1786), .IN1(r796_n128), .IN2(r796_n129) );
  NAND2X0 r796_U133 ( .IN1(n7089), .IN2(r796_n127), .QN(r796_n124) );
  OR2X1 r796_U132 ( .IN2(n7089), .IN1(r796_n127), .Q(r796_n126) );
  NAND2X0 r796_U131 ( .IN1(P1_N1634), .IN2(r796_n126), .QN(r796_n125) );
  NAND2X0 r796_U130 ( .IN1(r796_n124), .IN2(r796_n125), .QN(r796_n117) );
  OR2X1 r796_U128 ( .IN2(P1_N1635), .IN1(n7144), .Q(r796_n121) );
  NAND2X0 r796_U127 ( .IN1(P1_N1635), .IN2(n7144), .QN(r796_n122) );
  NAND2X0 r796_U126 ( .IN1(r796_n121), .IN2(r796_n122), .QN(r796_n120) );
  NOR2X0 r796_U125 ( .QN(r796_n118), .IN1(r796_n117), .IN2(r796_n120) );
  AND2X1 r796_U124 ( .IN1(r796_n117), .IN2(r796_n120), .Q(r796_n119) );
  NOR2X0 r796_U123 ( .QN(P1_N1787), .IN1(r796_n118), .IN2(r796_n119) );
  NAND2X0 r796_U122 ( .IN1(n7141), .IN2(r796_n117), .QN(r796_n114) );
  OR2X1 r796_U121 ( .IN2(n7141), .IN1(r796_n117), .Q(r796_n116) );
  NAND2X0 r796_U120 ( .IN1(P1_N1635), .IN2(r796_n116), .QN(r796_n115) );
  NAND2X0 r796_U119 ( .IN1(r796_n114), .IN2(r796_n115), .QN(r796_n107) );
  OR2X1 r796_U117 ( .IN2(P1_N1636), .IN1(n7136), .Q(r796_n111) );
  NAND2X0 r796_U116 ( .IN1(P1_N1636), .IN2(n7136), .QN(r796_n112) );
  NAND2X0 r796_U115 ( .IN1(r796_n111), .IN2(r796_n112), .QN(r796_n110) );
  NOR2X0 r796_U114 ( .QN(r796_n108), .IN1(r796_n107), .IN2(r796_n110) );
  AND2X1 r796_U113 ( .IN1(r796_n107), .IN2(r796_n110), .Q(r796_n109) );
  NOR2X0 r796_U112 ( .QN(P1_N1788), .IN1(r796_n108), .IN2(r796_n109) );
  NAND2X0 r796_U111 ( .IN1(n7138), .IN2(r796_n107), .QN(r796_n104) );
  OR2X1 r796_U110 ( .IN2(n7138), .IN1(r796_n107), .Q(r796_n106) );
  NAND2X0 r796_U109 ( .IN1(P1_N1636), .IN2(r796_n106), .QN(r796_n105) );
  NAND2X0 r796_U294 ( .IN1(P1_N5155), .IN2(r796_n24), .QN(r796_n270) );
  OR2X1 r796_U293 ( .IN2(P1_N5155), .IN1(r796_n24), .Q(r796_n272) );
  NAND2X0 r796_U292 ( .IN1(P1_N1618), .IN2(r796_n272), .QN(r796_n271) );
  NAND2X0 r796_U291 ( .IN1(r796_n270), .IN2(r796_n271), .QN(r796_n17) );
  NAND2X0 r796_U290 ( .IN1(n7075), .IN2(r796_n17), .QN(r796_n267) );
  OR2X1 r796_U289 ( .IN2(n7075), .IN1(r796_n17), .Q(r796_n269) );
  NAND2X0 r796_U288 ( .IN1(P1_N1619), .IN2(r796_n269), .QN(r796_n268) );
  NAND2X0 r796_U287 ( .IN1(r796_n267), .IN2(r796_n268), .QN(r796_n10) );
  NAND2X0 r796_U286 ( .IN1(n7072), .IN2(r796_n10), .QN(r796_n264) );
  OR2X1 r796_U285 ( .IN2(n7072), .IN1(r796_n10), .Q(r796_n266) );
  NAND2X0 r796_U284 ( .IN1(P1_N1620), .IN2(r796_n266), .QN(r796_n265) );
  NAND2X0 r796_U283 ( .IN1(r796_n264), .IN2(r796_n265), .QN(r796_n3) );
  NAND2X0 r796_U282 ( .IN1(P1_N5158), .IN2(r796_n3), .QN(r796_n261) );
  OR2X1 r796_U281 ( .IN2(P1_N5158), .IN1(r796_n3), .Q(r796_n263) );
  NAND2X0 r796_U280 ( .IN1(P1_N1621), .IN2(r796_n263), .QN(r796_n262) );
  NAND2X0 r796_U279 ( .IN1(r796_n261), .IN2(r796_n262), .QN(r796_n254) );
  OR2X1 r796_U277 ( .IN2(P1_N1622), .IN1(n7067), .Q(r796_n258) );
  NAND2X0 r796_U276 ( .IN1(P1_N1622), .IN2(n7067), .QN(r796_n259) );
  NAND2X0 r796_U275 ( .IN1(r796_n258), .IN2(r796_n259), .QN(r796_n257) );
  NOR2X0 r796_U274 ( .QN(r796_n255), .IN1(r796_n254), .IN2(r796_n257) );
  AND2X1 r796_U273 ( .IN1(r796_n254), .IN2(r796_n257), .Q(r796_n256) );
  NOR2X0 r796_U272 ( .QN(P1_N1774), .IN1(r796_n255), .IN2(r796_n256) );
  NAND2X0 r796_U271 ( .IN1(n7066), .IN2(r796_n254), .QN(r796_n251) );
  OR2X1 r796_U270 ( .IN2(n7066), .IN1(r796_n254), .Q(r796_n253) );
  NAND2X0 r796_U269 ( .IN1(P1_N1622), .IN2(r796_n253), .QN(r796_n252) );
  NAND2X0 r796_U268 ( .IN1(r796_n251), .IN2(r796_n252), .QN(r796_n244) );
  OR2X1 r796_U266 ( .IN2(P1_N1623), .IN1(n7063), .Q(r796_n248) );
  NAND2X0 r796_U265 ( .IN1(P1_N1623), .IN2(n7063), .QN(r796_n249) );
  NAND2X0 r796_U264 ( .IN1(r796_n248), .IN2(r796_n249), .QN(r796_n247) );
  NOR2X0 r796_U263 ( .QN(r796_n245), .IN1(r796_n244), .IN2(r796_n247) );
  AND2X1 r796_U262 ( .IN1(r796_n244), .IN2(r796_n247), .Q(r796_n246) );
  NOR2X0 r796_U261 ( .QN(P1_N1775), .IN1(r796_n245), .IN2(r796_n246) );
  NAND2X0 r796_U260 ( .IN1(n7062), .IN2(r796_n244), .QN(r796_n241) );
  OR2X1 r796_U259 ( .IN2(n7062), .IN1(r796_n244), .Q(r796_n243) );
  NAND2X0 r796_U258 ( .IN1(P1_N1623), .IN2(r796_n243), .QN(r796_n242) );
  NAND2X0 r796_U257 ( .IN1(r796_n241), .IN2(r796_n242), .QN(r796_n234) );
  OR2X1 r796_U255 ( .IN2(P1_N1624), .IN1(n7058), .Q(r796_n238) );
  NAND2X0 r796_U254 ( .IN1(P1_N1624), .IN2(n7058), .QN(r796_n239) );
  NAND2X0 r796_U253 ( .IN1(r796_n238), .IN2(r796_n239), .QN(r796_n237) );
  NOR2X0 r796_U252 ( .QN(r796_n235), .IN1(r796_n234), .IN2(r796_n237) );
  AND2X1 r796_U251 ( .IN1(r796_n234), .IN2(r796_n237), .Q(r796_n236) );
  NOR2X0 r796_U250 ( .QN(P1_N1776), .IN1(r796_n235), .IN2(r796_n236) );
  NAND2X0 r796_U249 ( .IN1(n7059), .IN2(r796_n234), .QN(r796_n231) );
  OR2X1 r796_U248 ( .IN2(n7059), .IN1(r796_n234), .Q(r796_n233) );
  NAND2X0 r796_U247 ( .IN1(P1_N1624), .IN2(r796_n233), .QN(r796_n232) );
  NAND2X0 r796_U246 ( .IN1(r796_n231), .IN2(r796_n232), .QN(r796_n224) );
  OR2X1 r796_U244 ( .IN2(P1_N1625), .IN1(n7056), .Q(r796_n228) );
  NAND2X0 r796_U243 ( .IN1(P1_N1625), .IN2(n7056), .QN(r796_n229) );
  NAND2X0 r796_U242 ( .IN1(r796_n228), .IN2(r796_n229), .QN(r796_n227) );
  NOR2X0 r796_U241 ( .QN(r796_n225), .IN1(r796_n224), .IN2(r796_n227) );
  AND2X1 r796_U240 ( .IN1(r796_n224), .IN2(r796_n227), .Q(r796_n226) );
  NOR2X0 r796_U239 ( .QN(P1_N1777), .IN1(r796_n225), .IN2(r796_n226) );
  NAND2X0 r796_U238 ( .IN1(P1_N5162), .IN2(r796_n224), .QN(r796_n221) );
  OR2X1 r796_U237 ( .IN2(P1_N5162), .IN1(r796_n224), .Q(r796_n223) );
  NAND2X0 r796_U236 ( .IN1(P1_N1625), .IN2(r796_n223), .QN(r796_n222) );
  NAND2X0 r796_U235 ( .IN1(r796_n221), .IN2(r796_n222), .QN(r796_n214) );
  OR2X1 r796_U233 ( .IN2(P1_N1626), .IN1(n7115), .Q(r796_n218) );
  NAND2X0 r796_U232 ( .IN1(P1_N1626), .IN2(n7115), .QN(r796_n219) );
  NAND2X0 r796_U231 ( .IN1(r796_n218), .IN2(r796_n219), .QN(r796_n217) );
  NOR2X0 r796_U230 ( .QN(r796_n215), .IN1(r796_n214), .IN2(r796_n217) );
  AND2X1 r796_U229 ( .IN1(r796_n214), .IN2(r796_n217), .Q(r796_n216) );
  NOR2X0 r796_U228 ( .QN(P1_N1778), .IN1(r796_n215), .IN2(r796_n216) );
  NAND2X0 r796_U227 ( .IN1(P1_N5163), .IN2(r796_n214), .QN(r796_n211) );
  OR2X1 r796_U226 ( .IN2(P1_N5163), .IN1(r796_n214), .Q(r796_n213) );
  NAND2X0 r796_U225 ( .IN1(P1_N1626), .IN2(r796_n213), .QN(r796_n212) );
  NAND2X0 r796_U224 ( .IN1(r796_n211), .IN2(r796_n212), .QN(r796_n204) );
  OR2X1 r796_U222 ( .IN2(P1_N1627), .IN1(n7112), .Q(r796_n208) );
  NAND2X0 r796_U221 ( .IN1(P1_N1627), .IN2(n7112), .QN(r796_n209) );
  NAND2X0 r796_U220 ( .IN1(r796_n208), .IN2(r796_n209), .QN(r796_n207) );
  NOR2X0 r796_U219 ( .QN(r796_n205), .IN1(r796_n204), .IN2(r796_n207) );
  AND2X1 r796_U218 ( .IN1(r796_n204), .IN2(r796_n207), .Q(r796_n206) );
  NOR2X0 r796_U217 ( .QN(P1_N1779), .IN1(r796_n205), .IN2(r796_n206) );
  NAND2X0 r796_U216 ( .IN1(P1_N5164), .IN2(r796_n204), .QN(r796_n201) );
  OR2X1 r796_U215 ( .IN2(P1_N5164), .IN1(r796_n204), .Q(r796_n203) );
  NAND2X0 r796_U214 ( .IN1(P1_N1627), .IN2(r796_n203), .QN(r796_n202) );
  NAND2X0 r796_U213 ( .IN1(r796_n201), .IN2(r796_n202), .QN(r796_n194) );
  OR2X1 r796_U211 ( .IN2(P1_N1628), .IN1(n7109), .Q(r796_n198) );
  NAND2X0 r796_U210 ( .IN1(P1_N1628), .IN2(n7109), .QN(r796_n199) );
  NAND2X0 r796_U209 ( .IN1(r796_n198), .IN2(r796_n199), .QN(r796_n197) );
  NOR2X0 r796_U208 ( .QN(r796_n195), .IN1(r796_n194), .IN2(r796_n197) );
  AND2X1 r796_U207 ( .IN1(r796_n194), .IN2(r796_n197), .Q(r796_n196) );
  NOR2X0 r796_U206 ( .QN(P1_N1780), .IN1(r796_n195), .IN2(r796_n196) );
  NAND2X0 r796_U205 ( .IN1(P1_N5165), .IN2(r796_n194), .QN(r796_n191) );
  OR2X1 r796_U204 ( .IN2(P1_N5165), .IN1(r796_n194), .Q(r796_n193) );
  NAND2X0 r796_U203 ( .IN1(P1_N1628), .IN2(r796_n193), .QN(r796_n192) );
  NAND2X0 r796_U202 ( .IN1(r796_n191), .IN2(r796_n192), .QN(r796_n184) );
  OR2X1 r796_U319 ( .IN2(P1_N1612), .IN1(n4803), .Q(r796_n288) );
  NAND2X0 r796_U318 ( .IN1(P1_N1612), .IN2(n4803), .QN(r796_n289) );
  NAND2X0 r796_U317 ( .IN1(r796_n288), .IN2(r796_n289), .QN(P1_N1764) );
  NAND2X0 r796_U315 ( .IN1(P1_N1612), .IN2(n7034), .QN(r796_n161) );
  OR2X1 r796_U314 ( .IN2(r796_n161), .IN1(n7051), .Q(r796_n285) );
  NAND2X0 r796_U313 ( .IN1(n7051), .IN2(r796_n161), .QN(r796_n287) );
  NAND2X0 r796_U312 ( .IN1(P1_N1613), .IN2(r796_n287), .QN(r796_n286) );
  NAND2X0 r796_U311 ( .IN1(r796_n285), .IN2(r796_n286), .QN(r796_n52) );
  NAND2X0 r796_U310 ( .IN1(P1_N5151), .IN2(r796_n52), .QN(r796_n282) );
  OR2X1 r796_U309 ( .IN2(P1_N5151), .IN1(r796_n52), .Q(r796_n284) );
  NAND2X0 r796_U308 ( .IN1(P1_N1614), .IN2(r796_n284), .QN(r796_n283) );
  NAND2X0 r796_U307 ( .IN1(r796_n282), .IN2(r796_n283), .QN(r796_n45) );
  NAND2X0 r796_U306 ( .IN1(n7041), .IN2(r796_n45), .QN(r796_n279) );
  OR2X1 r796_U305 ( .IN2(n7041), .IN1(r796_n45), .Q(r796_n281) );
  NAND2X0 r796_U304 ( .IN1(P1_N1615), .IN2(r796_n281), .QN(r796_n280) );
  NAND2X0 r796_U303 ( .IN1(r796_n279), .IN2(r796_n280), .QN(r796_n38) );
  NAND2X0 r796_U302 ( .IN1(n7036), .IN2(r796_n38), .QN(r796_n276) );
  OR2X1 r796_U301 ( .IN2(n7036), .IN1(r796_n38), .Q(r796_n278) );
  NAND2X0 r796_U300 ( .IN1(P1_N1616), .IN2(r796_n278), .QN(r796_n277) );
  NAND2X0 r796_U299 ( .IN1(r796_n276), .IN2(r796_n277), .QN(r796_n31) );
  NAND2X0 r796_U298 ( .IN1(P1_N5154), .IN2(r796_n31), .QN(r796_n273) );
  OR2X1 r796_U297 ( .IN2(P1_N5154), .IN1(r796_n31), .Q(r796_n275) );
  NAND2X0 r796_U296 ( .IN1(P1_N1617), .IN2(r796_n275), .QN(r796_n274) );
  NAND2X0 r796_U295 ( .IN1(r796_n273), .IN2(r796_n274), .QN(r796_n24) );
  OR2X1 r798_U55 ( .IN2(P1_N1987), .IN1(n7045), .Q(r798_n54) );
  NAND2X0 r798_U54 ( .IN1(P1_N1987), .IN2(n7045), .QN(r798_n55) );
  NAND2X0 r798_U53 ( .IN1(r798_n54), .IN2(r798_n55), .QN(r798_n53) );
  NOR2X0 r798_U52 ( .QN(r798_n50), .IN1(r798_n52), .IN2(r798_n53) );
  AND2X1 r798_U51 ( .IN1(r798_n52), .IN2(r798_n53), .Q(r798_n51) );
  NOR2X0 r798_U50 ( .QN(P1_N2139), .IN1(r798_n50), .IN2(r798_n51) );
  OR2X1 r798_U48 ( .IN2(P1_N1988), .IN1(n7043), .Q(r798_n47) );
  NAND2X0 r798_U47 ( .IN1(P1_N1988), .IN2(n7043), .QN(r798_n48) );
  NAND2X0 r798_U46 ( .IN1(r798_n47), .IN2(r798_n48), .QN(r798_n46) );
  NOR2X0 r798_U45 ( .QN(r798_n43), .IN1(r798_n45), .IN2(r798_n46) );
  AND2X1 r798_U44 ( .IN1(r798_n45), .IN2(r798_n46), .Q(r798_n44) );
  NOR2X0 r798_U43 ( .QN(P1_N2140), .IN1(r798_n43), .IN2(r798_n44) );
  OR2X1 r798_U41 ( .IN2(P1_N1989), .IN1(n7037), .Q(r798_n40) );
  NAND2X0 r798_U40 ( .IN1(P1_N1989), .IN2(n7037), .QN(r798_n41) );
  NAND2X0 r798_U39 ( .IN1(r798_n40), .IN2(r798_n41), .QN(r798_n39) );
  NOR2X0 r798_U38 ( .QN(r798_n36), .IN1(r798_n38), .IN2(r798_n39) );
  AND2X1 r798_U37 ( .IN1(r798_n38), .IN2(r798_n39), .Q(r798_n37) );
  NOR2X0 r798_U36 ( .QN(P1_N2141), .IN1(r798_n36), .IN2(r798_n37) );
  OR2X1 r798_U34 ( .IN2(P1_N1990), .IN1(n7082), .Q(r798_n33) );
  NAND2X0 r798_U33 ( .IN1(P1_N1990), .IN2(n7082), .QN(r798_n34) );
  NAND2X0 r798_U32 ( .IN1(r798_n33), .IN2(r798_n34), .QN(r798_n32) );
  NOR2X0 r798_U31 ( .QN(r798_n29), .IN1(r798_n31), .IN2(r798_n32) );
  AND2X1 r798_U30 ( .IN1(r798_n31), .IN2(r798_n32), .Q(r798_n30) );
  NOR2X0 r798_U29 ( .QN(P1_N2142), .IN1(r798_n29), .IN2(r798_n30) );
  OR2X1 r798_U27 ( .IN2(P1_N1991), .IN1(n7079), .Q(r798_n26) );
  NAND2X0 r798_U26 ( .IN1(P1_N1991), .IN2(n7079), .QN(r798_n27) );
  NAND2X0 r798_U25 ( .IN1(r798_n26), .IN2(r798_n27), .QN(r798_n25) );
  NOR2X0 r798_U24 ( .QN(r798_n22), .IN1(r798_n24), .IN2(r798_n25) );
  AND2X1 r798_U23 ( .IN1(r798_n24), .IN2(r798_n25), .Q(r798_n23) );
  NOR2X0 r798_U22 ( .QN(P1_N2143), .IN1(r798_n22), .IN2(r798_n23) );
  OR2X1 r798_U20 ( .IN2(P1_N1992), .IN1(n7076), .Q(r798_n19) );
  NAND2X0 r798_U19 ( .IN1(P1_N1992), .IN2(n7076), .QN(r798_n20) );
  NAND2X0 r798_U18 ( .IN1(r798_n19), .IN2(r798_n20), .QN(r798_n18) );
  NOR2X0 r798_U17 ( .QN(r798_n15), .IN1(r798_n17), .IN2(r798_n18) );
  AND2X1 r798_U16 ( .IN1(r798_n17), .IN2(r798_n18), .Q(r798_n16) );
  NOR2X0 r798_U15 ( .QN(P1_N2144), .IN1(r798_n15), .IN2(r798_n16) );
  OR2X1 r798_U13 ( .IN2(P1_N1993), .IN1(n7073), .Q(r798_n12) );
  NAND2X0 r798_U12 ( .IN1(P1_N1993), .IN2(n7073), .QN(r798_n13) );
  NAND2X0 r798_U11 ( .IN1(r798_n12), .IN2(r798_n13), .QN(r798_n11) );
  NOR2X0 r798_U10 ( .QN(r798_n8), .IN1(r798_n10), .IN2(r798_n11) );
  AND2X1 r798_U9 ( .IN1(r798_n10), .IN2(r798_n11), .Q(r798_n9) );
  NOR2X0 r798_U8 ( .QN(P1_N2145), .IN1(r798_n8), .IN2(r798_n9) );
  OR2X1 r798_U6 ( .IN2(P1_N1994), .IN1(n7071), .Q(r798_n5) );
  NAND2X0 r798_U5 ( .IN1(P1_N1994), .IN2(n7071), .QN(r798_n6) );
  NAND2X0 r798_U4 ( .IN1(r798_n5), .IN2(r798_n6), .QN(r798_n4) );
  NOR2X0 r798_U3 ( .QN(r798_n1), .IN1(r798_n3), .IN2(r798_n4) );
  AND2X1 r798_U2 ( .IN1(r798_n3), .IN2(r798_n4), .Q(r798_n2) );
  NOR2X0 r798_U1 ( .QN(P1_N2146), .IN1(r798_n1), .IN2(r798_n2) );
  NAND2X0 r798_U149 ( .IN1(P1_N2006), .IN2(n7092), .QN(r798_n142) );
  NAND2X0 r798_U148 ( .IN1(r798_n141), .IN2(r798_n142), .QN(r798_n140) );
  NOR2X0 r798_U147 ( .QN(r798_n138), .IN1(r798_n137), .IN2(r798_n140) );
  AND2X1 r798_U146 ( .IN1(r798_n137), .IN2(r798_n140), .Q(r798_n139) );
  NOR2X0 r798_U145 ( .QN(P1_N2158), .IN1(r798_n138), .IN2(r798_n139) );
  NAND2X0 r798_U144 ( .IN1(P1_N5170), .IN2(r798_n137), .QN(r798_n134) );
  OR2X1 r798_U143 ( .IN2(P1_N5170), .IN1(r798_n137), .Q(r798_n136) );
  NAND2X0 r798_U142 ( .IN1(P1_N2006), .IN2(r798_n136), .QN(r798_n135) );
  NAND2X0 r798_U141 ( .IN1(r798_n134), .IN2(r798_n135), .QN(r798_n127) );
  OR2X1 r798_U139 ( .IN2(P1_N2007), .IN1(n7090), .Q(r798_n131) );
  NAND2X0 r798_U138 ( .IN1(P1_N2007), .IN2(n7090), .QN(r798_n132) );
  NAND2X0 r798_U137 ( .IN1(r798_n131), .IN2(r798_n132), .QN(r798_n130) );
  NOR2X0 r798_U136 ( .QN(r798_n128), .IN1(r798_n127), .IN2(r798_n130) );
  AND2X1 r798_U135 ( .IN1(r798_n127), .IN2(r798_n130), .Q(r798_n129) );
  NOR2X0 r798_U134 ( .QN(P1_N2159), .IN1(r798_n128), .IN2(r798_n129) );
  NAND2X0 r798_U133 ( .IN1(n7089), .IN2(r798_n127), .QN(r798_n124) );
  OR2X1 r798_U132 ( .IN2(n7089), .IN1(r798_n127), .Q(r798_n126) );
  NAND2X0 r798_U131 ( .IN1(P1_N2007), .IN2(r798_n126), .QN(r798_n125) );
  NAND2X0 r798_U130 ( .IN1(r798_n124), .IN2(r798_n125), .QN(r798_n117) );
  OR2X1 r798_U128 ( .IN2(P1_N2008), .IN1(n7144), .Q(r798_n121) );
  NAND2X0 r798_U127 ( .IN1(P1_N2008), .IN2(n7144), .QN(r798_n122) );
  NAND2X0 r798_U126 ( .IN1(r798_n121), .IN2(r798_n122), .QN(r798_n120) );
  NOR2X0 r798_U125 ( .QN(r798_n118), .IN1(r798_n117), .IN2(r798_n120) );
  AND2X1 r798_U124 ( .IN1(r798_n117), .IN2(r798_n120), .Q(r798_n119) );
  NOR2X0 r798_U123 ( .QN(P1_N2160), .IN1(r798_n118), .IN2(r798_n119) );
  NAND2X0 r798_U122 ( .IN1(n7141), .IN2(r798_n117), .QN(r798_n114) );
  OR2X1 r798_U121 ( .IN2(n7141), .IN1(r798_n117), .Q(r798_n116) );
  NAND2X0 r798_U120 ( .IN1(P1_N2008), .IN2(r798_n116), .QN(r798_n115) );
  NAND2X0 r798_U119 ( .IN1(r798_n114), .IN2(r798_n115), .QN(r798_n107) );
  OR2X1 r798_U117 ( .IN2(P1_N2009), .IN1(r798_n314), .Q(r798_n111) );
  NAND2X0 r798_U116 ( .IN1(P1_N2009), .IN2(r798_n314), .QN(r798_n112) );
  NAND2X0 r798_U115 ( .IN1(r798_n111), .IN2(r798_n112), .QN(r798_n110) );
  NOR2X0 r798_U114 ( .QN(r798_n108), .IN1(r798_n107), .IN2(r798_n110) );
  AND2X1 r798_U113 ( .IN1(r798_n107), .IN2(r798_n110), .Q(r798_n109) );
  NOR2X0 r798_U112 ( .QN(P1_N2161), .IN1(r798_n108), .IN2(r798_n109) );
  NAND2X0 r798_U111 ( .IN1(n7138), .IN2(r798_n107), .QN(r798_n104) );
  OR2X1 r798_U110 ( .IN2(n7138), .IN1(r798_n107), .Q(r798_n106) );
  NAND2X0 r798_U109 ( .IN1(P1_N2009), .IN2(r798_n106), .QN(r798_n105) );
  NAND2X0 r798_U108 ( .IN1(r798_n104), .IN2(r798_n105), .QN(r798_n97) );
  OR2X1 r798_U106 ( .IN2(P1_N2010), .IN1(n7130), .Q(r798_n101) );
  NAND2X0 r798_U105 ( .IN1(P1_N2010), .IN2(n7130), .QN(r798_n102) );
  NAND2X0 r798_U104 ( .IN1(r798_n101), .IN2(r798_n102), .QN(r798_n100) );
  NOR2X0 r798_U103 ( .QN(r798_n98), .IN1(r798_n97), .IN2(r798_n100) );
  AND2X1 r798_U102 ( .IN1(r798_n97), .IN2(r798_n100), .Q(r798_n99) );
  NOR2X0 r798_U101 ( .QN(P1_N2162), .IN1(r798_n98), .IN2(r798_n99) );
  NAND2X0 r798_U100 ( .IN1(P1_N5174), .IN2(r798_n97), .QN(r798_n94) );
  OR2X1 r798_U99 ( .IN2(P1_N5174), .IN1(r798_n97), .Q(r798_n96) );
  NAND2X0 r798_U98 ( .IN1(P1_N2010), .IN2(r798_n96), .QN(r798_n95) );
  NAND2X0 r798_U97 ( .IN1(r798_n94), .IN2(r798_n95), .QN(r798_n87) );
  OR2X1 r798_U95 ( .IN2(P1_N2011), .IN1(n7125), .Q(r798_n91) );
  NAND2X0 r798_U94 ( .IN1(P1_N2011), .IN2(n7125), .QN(r798_n92) );
  NAND2X0 r798_U93 ( .IN1(r798_n91), .IN2(r798_n92), .QN(r798_n90) );
  NOR2X0 r798_U92 ( .QN(r798_n88), .IN1(r798_n87), .IN2(r798_n90) );
  AND2X1 r798_U91 ( .IN1(r798_n87), .IN2(r798_n90), .Q(r798_n89) );
  NOR2X0 r798_U90 ( .QN(P1_N2163), .IN1(r798_n88), .IN2(r798_n89) );
  NAND2X0 r798_U89 ( .IN1(n7124), .IN2(r798_n87), .QN(r798_n84) );
  OR2X1 r798_U88 ( .IN2(n7124), .IN1(r798_n87), .Q(r798_n86) );
  NAND2X0 r798_U87 ( .IN1(P1_N2011), .IN2(r798_n86), .QN(r798_n85) );
  NAND2X0 r798_U86 ( .IN1(r798_n84), .IN2(r798_n85), .QN(r798_n77) );
  OR2X1 r798_U84 ( .IN2(P1_N2012), .IN1(n7119), .Q(r798_n81) );
  NAND2X0 r798_U83 ( .IN1(P1_N2012), .IN2(n7119), .QN(r798_n82) );
  NAND2X0 r798_U82 ( .IN1(r798_n81), .IN2(r798_n82), .QN(r798_n80) );
  NOR2X0 r798_U81 ( .QN(r798_n78), .IN1(r798_n77), .IN2(r798_n80) );
  AND2X1 r798_U80 ( .IN1(r798_n77), .IN2(r798_n80), .Q(r798_n79) );
  NOR2X0 r798_U79 ( .QN(P1_N2164), .IN1(r798_n78), .IN2(r798_n79) );
  NAND2X0 r798_U78 ( .IN1(P1_N5176), .IN2(r798_n77), .QN(r798_n74) );
  OR2X1 r798_U77 ( .IN2(P1_N5176), .IN1(r798_n77), .Q(r798_n76) );
  NAND2X0 r798_U76 ( .IN1(P1_N2012), .IN2(r798_n76), .QN(r798_n75) );
  NAND2X0 r798_U75 ( .IN1(r798_n74), .IN2(r798_n75), .QN(r798_n64) );
  OR2X1 r798_U73 ( .IN2(P1_N2013), .IN1(n7117), .Q(r798_n71) );
  NAND2X0 r798_U72 ( .IN1(P1_N2013), .IN2(n7117), .QN(r798_n72) );
  NAND2X0 r798_U71 ( .IN1(r798_n71), .IN2(r798_n72), .QN(r798_n70) );
  NOR2X0 r798_U70 ( .QN(r798_n68), .IN1(r798_n64), .IN2(r798_n70) );
  AND2X1 r798_U69 ( .IN1(r798_n64), .IN2(r798_n70), .Q(r798_n69) );
  NOR2X0 r798_U68 ( .QN(P1_N2165), .IN1(r798_n68), .IN2(r798_n69) );
  OR2X1 r798_U66 ( .IN2(P1_N2014), .IN1(n7146), .Q(r798_n65) );
  NAND2X0 r798_U65 ( .IN1(P1_N2014), .IN2(n7146), .QN(r798_n66) );
  NAND2X0 r798_U64 ( .IN1(r798_n65), .IN2(r798_n66), .QN(r798_n60) );
  NAND2X0 r798_U63 ( .IN1(P1_N5177), .IN2(r798_n64), .QN(r798_n61) );
  OR2X1 r798_U62 ( .IN2(P1_N5177), .IN1(r798_n64), .Q(r798_n63) );
  NAND2X0 r798_U61 ( .IN1(P1_N2013), .IN2(r798_n63), .QN(r798_n62) );
  NAND2X0 r798_U60 ( .IN1(r798_n61), .IN2(r798_n62), .QN(r798_n59) );
  NOR2X0 r798_U59 ( .QN(r798_n57), .IN1(r798_n60), .IN2(r798_n59) );
  AND2X1 r798_U58 ( .IN1(r798_n59), .IN2(r798_n60), .Q(r798_n58) );
  NOR2X0 r798_U57 ( .QN(P1_N2166), .IN1(r798_n57), .IN2(r798_n58) );
  NAND2X0 r798_U242 ( .IN1(r798_n228), .IN2(r798_n229), .QN(r798_n227) );
  NOR2X0 r798_U241 ( .QN(r798_n225), .IN1(r798_n224), .IN2(r798_n227) );
  AND2X1 r798_U240 ( .IN1(r798_n224), .IN2(r798_n227), .Q(r798_n226) );
  NOR2X0 r798_U239 ( .QN(P1_N2150), .IN1(r798_n225), .IN2(r798_n226) );
  NAND2X0 r798_U238 ( .IN1(P1_N5162), .IN2(r798_n224), .QN(r798_n221) );
  OR2X1 r798_U237 ( .IN2(P1_N5162), .IN1(r798_n224), .Q(r798_n223) );
  NAND2X0 r798_U236 ( .IN1(P1_N1998), .IN2(r798_n223), .QN(r798_n222) );
  NAND2X0 r798_U235 ( .IN1(r798_n221), .IN2(r798_n222), .QN(r798_n214) );
  OR2X1 r798_U233 ( .IN2(P1_N1999), .IN1(n7115), .Q(r798_n218) );
  NAND2X0 r798_U232 ( .IN1(P1_N1999), .IN2(n7115), .QN(r798_n219) );
  NAND2X0 r798_U231 ( .IN1(r798_n218), .IN2(r798_n219), .QN(r798_n217) );
  NOR2X0 r798_U230 ( .QN(r798_n215), .IN1(r798_n214), .IN2(r798_n217) );
  AND2X1 r798_U229 ( .IN1(r798_n214), .IN2(r798_n217), .Q(r798_n216) );
  NOR2X0 r798_U228 ( .QN(P1_N2151), .IN1(r798_n215), .IN2(r798_n216) );
  NAND2X0 r798_U227 ( .IN1(P1_N5163), .IN2(r798_n214), .QN(r798_n211) );
  OR2X1 r798_U226 ( .IN2(P1_N5163), .IN1(r798_n214), .Q(r798_n213) );
  NAND2X0 r798_U225 ( .IN1(P1_N1999), .IN2(r798_n213), .QN(r798_n212) );
  NAND2X0 r798_U224 ( .IN1(r798_n211), .IN2(r798_n212), .QN(r798_n204) );
  OR2X1 r798_U222 ( .IN2(P1_N2000), .IN1(n7112), .Q(r798_n208) );
  NAND2X0 r798_U221 ( .IN1(P1_N2000), .IN2(n7112), .QN(r798_n209) );
  NAND2X0 r798_U220 ( .IN1(r798_n208), .IN2(r798_n209), .QN(r798_n207) );
  NOR2X0 r798_U219 ( .QN(r798_n205), .IN1(r798_n204), .IN2(r798_n207) );
  AND2X1 r798_U218 ( .IN1(r798_n204), .IN2(r798_n207), .Q(r798_n206) );
  NOR2X0 r798_U217 ( .QN(P1_N2152), .IN1(r798_n205), .IN2(r798_n206) );
  NAND2X0 r798_U216 ( .IN1(P1_N5164), .IN2(r798_n204), .QN(r798_n201) );
  OR2X1 r798_U215 ( .IN2(P1_N5164), .IN1(r798_n204), .Q(r798_n203) );
  NAND2X0 r798_U214 ( .IN1(P1_N2000), .IN2(r798_n203), .QN(r798_n202) );
  NAND2X0 r798_U213 ( .IN1(r798_n201), .IN2(r798_n202), .QN(r798_n194) );
  OR2X1 r798_U211 ( .IN2(P1_N2001), .IN1(n7109), .Q(r798_n198) );
  NAND2X0 r798_U210 ( .IN1(P1_N2001), .IN2(n7109), .QN(r798_n199) );
  NAND2X0 r798_U209 ( .IN1(r798_n198), .IN2(r798_n199), .QN(r798_n197) );
  NOR2X0 r798_U208 ( .QN(r798_n195), .IN1(r798_n194), .IN2(r798_n197) );
  AND2X1 r798_U207 ( .IN1(r798_n194), .IN2(r798_n197), .Q(r798_n196) );
  NOR2X0 r798_U206 ( .QN(P1_N2153), .IN1(r798_n195), .IN2(r798_n196) );
  NAND2X0 r798_U205 ( .IN1(P1_N5165), .IN2(r798_n194), .QN(r798_n191) );
  OR2X1 r798_U204 ( .IN2(P1_N5165), .IN1(r798_n194), .Q(r798_n193) );
  NAND2X0 r798_U203 ( .IN1(P1_N2001), .IN2(r798_n193), .QN(r798_n192) );
  NAND2X0 r798_U202 ( .IN1(r798_n191), .IN2(r798_n192), .QN(r798_n184) );
  OR2X1 r798_U200 ( .IN2(P1_N2002), .IN1(n7105), .Q(r798_n188) );
  NAND2X0 r798_U199 ( .IN1(P1_N2002), .IN2(n7105), .QN(r798_n189) );
  NAND2X0 r798_U198 ( .IN1(r798_n188), .IN2(r798_n189), .QN(r798_n187) );
  NOR2X0 r798_U197 ( .QN(r798_n185), .IN1(r798_n184), .IN2(r798_n187) );
  AND2X1 r798_U196 ( .IN1(r798_n184), .IN2(r798_n187), .Q(r798_n186) );
  NOR2X0 r798_U195 ( .QN(P1_N2154), .IN1(r798_n185), .IN2(r798_n186) );
  NAND2X0 r798_U194 ( .IN1(P1_N5166), .IN2(r798_n184), .QN(r798_n181) );
  OR2X1 r798_U193 ( .IN2(P1_N5166), .IN1(r798_n184), .Q(r798_n183) );
  NAND2X0 r798_U192 ( .IN1(P1_N2002), .IN2(r798_n183), .QN(r798_n182) );
  NAND2X0 r798_U191 ( .IN1(r798_n181), .IN2(r798_n182), .QN(r798_n174) );
  OR2X1 r798_U189 ( .IN2(P1_N2003), .IN1(n7102), .Q(r798_n178) );
  NAND2X0 r798_U188 ( .IN1(P1_N2003), .IN2(n7102), .QN(r798_n179) );
  NAND2X0 r798_U187 ( .IN1(r798_n178), .IN2(r798_n179), .QN(r798_n177) );
  NOR2X0 r798_U186 ( .QN(r798_n175), .IN1(r798_n174), .IN2(r798_n177) );
  AND2X1 r798_U185 ( .IN1(r798_n174), .IN2(r798_n177), .Q(r798_n176) );
  NOR2X0 r798_U184 ( .QN(P1_N2155), .IN1(r798_n175), .IN2(r798_n176) );
  NAND2X0 r798_U183 ( .IN1(P1_N5167), .IN2(r798_n174), .QN(r798_n171) );
  OR2X1 r798_U182 ( .IN2(P1_N5167), .IN1(r798_n174), .Q(r798_n173) );
  NAND2X0 r798_U181 ( .IN1(P1_N2003), .IN2(r798_n173), .QN(r798_n172) );
  NAND2X0 r798_U180 ( .IN1(r798_n171), .IN2(r798_n172), .QN(r798_n157) );
  OR2X1 r798_U178 ( .IN2(P1_N2004), .IN1(n7098), .Q(r798_n168) );
  NAND2X0 r798_U177 ( .IN1(P1_N2004), .IN2(n7098), .QN(r798_n169) );
  NAND2X0 r798_U176 ( .IN1(r798_n168), .IN2(r798_n169), .QN(r798_n167) );
  NOR2X0 r798_U175 ( .QN(r798_n165), .IN1(r798_n157), .IN2(r798_n167) );
  AND2X1 r798_U174 ( .IN1(r798_n157), .IN2(r798_n167), .Q(r798_n166) );
  NOR2X0 r798_U173 ( .QN(P1_N2156), .IN1(r798_n165), .IN2(r798_n166) );
  OR2X1 r798_U172 ( .IN2(P1_N1986), .IN1(n7048), .Q(r798_n162) );
  NAND2X0 r798_U171 ( .IN1(P1_N1986), .IN2(n7048), .QN(r798_n163) );
  NAND2X0 r798_U170 ( .IN1(r798_n162), .IN2(r798_n163), .QN(r798_n160) );
  NAND2X0 r798_U169 ( .IN1(r798_n160), .IN2(r798_n161), .QN(r798_n158) );
  OR2X1 r798_U168 ( .IN2(r798_n161), .IN1(r798_n160), .Q(r798_n159) );
  NAND2X0 r798_U167 ( .IN1(r798_n158), .IN2(r798_n159), .QN(P1_N2138) );
  NAND2X0 r798_U166 ( .IN1(n7099), .IN2(r798_n157), .QN(r798_n154) );
  OR2X1 r798_U165 ( .IN2(n7099), .IN1(r798_n157), .Q(r798_n156) );
  NAND2X0 r798_U164 ( .IN1(P1_N2004), .IN2(r798_n156), .QN(r798_n155) );
  NAND2X0 r798_U163 ( .IN1(r798_n154), .IN2(r798_n155), .QN(r798_n147) );
  OR2X1 r798_U161 ( .IN2(P1_N2005), .IN1(n7095), .Q(r798_n151) );
  NAND2X0 r798_U160 ( .IN1(P1_N2005), .IN2(n7095), .QN(r798_n152) );
  NAND2X0 r798_U159 ( .IN1(r798_n151), .IN2(r798_n152), .QN(r798_n150) );
  NOR2X0 r798_U158 ( .QN(r798_n148), .IN1(r798_n147), .IN2(r798_n150) );
  AND2X1 r798_U157 ( .IN1(r798_n147), .IN2(r798_n150), .Q(r798_n149) );
  NOR2X0 r798_U156 ( .QN(P1_N2157), .IN1(r798_n148), .IN2(r798_n149) );
  NAND2X0 r798_U155 ( .IN1(P1_N5169), .IN2(r798_n147), .QN(r798_n144) );
  OR2X1 r798_U154 ( .IN2(P1_N5169), .IN1(r798_n147), .Q(r798_n146) );
  NAND2X0 r798_U153 ( .IN1(P1_N2005), .IN2(r798_n146), .QN(r798_n145) );
  NAND2X0 r798_U152 ( .IN1(r798_n144), .IN2(r798_n145), .QN(r798_n137) );
  OR2X1 r798_U150 ( .IN2(P1_N2006), .IN1(n7092), .Q(r798_n141) );
  OR2X1 r798_U319 ( .IN2(P1_N1985), .IN1(n4803), .Q(r798_n288) );
  NAND2X0 r798_U318 ( .IN1(P1_N1985), .IN2(n4803), .QN(r798_n289) );
  NAND2X0 r798_U317 ( .IN1(r798_n288), .IN2(r798_n289), .QN(P1_N2137) );
  NAND2X0 r798_U315 ( .IN1(P1_N1985), .IN2(n7034), .QN(r798_n161) );
  OR2X1 r798_U314 ( .IN2(r798_n161), .IN1(n7048), .Q(r798_n285) );
  NAND2X0 r798_U313 ( .IN1(n7048), .IN2(r798_n161), .QN(r798_n287) );
  NAND2X0 r798_U312 ( .IN1(P1_N1986), .IN2(r798_n287), .QN(r798_n286) );
  NAND2X0 r798_U311 ( .IN1(r798_n285), .IN2(r798_n286), .QN(r798_n52) );
  NAND2X0 r798_U310 ( .IN1(P1_N5151), .IN2(r798_n52), .QN(r798_n282) );
  OR2X1 r798_U309 ( .IN2(P1_N5151), .IN1(r798_n52), .Q(r798_n284) );
  NAND2X0 r798_U308 ( .IN1(P1_N1987), .IN2(r798_n284), .QN(r798_n283) );
  NAND2X0 r798_U307 ( .IN1(r798_n282), .IN2(r798_n283), .QN(r798_n45) );
  NAND2X0 r798_U306 ( .IN1(n7041), .IN2(r798_n45), .QN(r798_n279) );
  OR2X1 r798_U305 ( .IN2(P1_N5152), .IN1(r798_n45), .Q(r798_n281) );
  NAND2X0 r798_U304 ( .IN1(P1_N1988), .IN2(r798_n281), .QN(r798_n280) );
  NAND2X0 r798_U303 ( .IN1(r798_n279), .IN2(r798_n280), .QN(r798_n38) );
  NAND2X0 r798_U302 ( .IN1(n7036), .IN2(r798_n38), .QN(r798_n276) );
  OR2X1 r798_U301 ( .IN2(n7036), .IN1(r798_n38), .Q(r798_n278) );
  NAND2X0 r798_U300 ( .IN1(P1_N1989), .IN2(r798_n278), .QN(r798_n277) );
  NAND2X0 r798_U299 ( .IN1(r798_n276), .IN2(r798_n277), .QN(r798_n31) );
  NAND2X0 r798_U298 ( .IN1(P1_N5154), .IN2(r798_n31), .QN(r798_n273) );
  OR2X1 r798_U297 ( .IN2(P1_N5154), .IN1(r798_n31), .Q(r798_n275) );
  NAND2X0 r798_U296 ( .IN1(P1_N1990), .IN2(r798_n275), .QN(r798_n274) );
  NAND2X0 r798_U295 ( .IN1(r798_n273), .IN2(r798_n274), .QN(r798_n24) );
  NAND2X0 r798_U294 ( .IN1(P1_N5155), .IN2(r798_n24), .QN(r798_n270) );
  OR2X1 r798_U293 ( .IN2(P1_N5155), .IN1(r798_n24), .Q(r798_n272) );
  NAND2X0 r798_U292 ( .IN1(P1_N1991), .IN2(r798_n272), .QN(r798_n271) );
  NAND2X0 r798_U291 ( .IN1(r798_n270), .IN2(r798_n271), .QN(r798_n17) );
  NAND2X0 r798_U290 ( .IN1(n7075), .IN2(r798_n17), .QN(r798_n267) );
  OR2X1 r798_U289 ( .IN2(n7075), .IN1(r798_n17), .Q(r798_n269) );
  NAND2X0 r798_U288 ( .IN1(P1_N1992), .IN2(r798_n269), .QN(r798_n268) );
  NAND2X0 r798_U287 ( .IN1(r798_n267), .IN2(r798_n268), .QN(r798_n10) );
  NAND2X0 r798_U286 ( .IN1(n7072), .IN2(r798_n10), .QN(r798_n264) );
  OR2X1 r798_U285 ( .IN2(n7072), .IN1(r798_n10), .Q(r798_n266) );
  NAND2X0 r798_U284 ( .IN1(P1_N1993), .IN2(r798_n266), .QN(r798_n265) );
  NAND2X0 r798_U283 ( .IN1(r798_n264), .IN2(r798_n265), .QN(r798_n3) );
  NAND2X0 r798_U282 ( .IN1(P1_N5158), .IN2(r798_n3), .QN(r798_n261) );
  OR2X1 r798_U281 ( .IN2(P1_N5158), .IN1(r798_n3), .Q(r798_n263) );
  NAND2X0 r798_U280 ( .IN1(P1_N1994), .IN2(r798_n263), .QN(r798_n262) );
  NAND2X0 r798_U279 ( .IN1(r798_n261), .IN2(r798_n262), .QN(r798_n254) );
  OR2X1 r798_U277 ( .IN2(P1_N1995), .IN1(n7067), .Q(r798_n258) );
  NAND2X0 r798_U276 ( .IN1(P1_N1995), .IN2(n7067), .QN(r798_n259) );
  NAND2X0 r798_U275 ( .IN1(r798_n258), .IN2(r798_n259), .QN(r798_n257) );
  NOR2X0 r798_U274 ( .QN(r798_n255), .IN1(r798_n254), .IN2(r798_n257) );
  AND2X1 r798_U273 ( .IN1(r798_n254), .IN2(r798_n257), .Q(r798_n256) );
  NOR2X0 r798_U272 ( .QN(P1_N2147), .IN1(r798_n255), .IN2(r798_n256) );
  NAND2X0 r798_U271 ( .IN1(P1_N5159), .IN2(r798_n254), .QN(r798_n251) );
  OR2X1 r798_U270 ( .IN2(P1_N5159), .IN1(r798_n254), .Q(r798_n253) );
  NAND2X0 r798_U269 ( .IN1(P1_N1995), .IN2(r798_n253), .QN(r798_n252) );
  NAND2X0 r798_U268 ( .IN1(r798_n251), .IN2(r798_n252), .QN(r798_n244) );
  OR2X1 r798_U266 ( .IN2(P1_N1996), .IN1(n7063), .Q(r798_n248) );
  NAND2X0 r798_U265 ( .IN1(P1_N1996), .IN2(n7063), .QN(r798_n249) );
  NAND2X0 r798_U264 ( .IN1(r798_n248), .IN2(r798_n249), .QN(r798_n247) );
  NOR2X0 r798_U263 ( .QN(r798_n245), .IN1(r798_n244), .IN2(r798_n247) );
  AND2X1 r798_U262 ( .IN1(r798_n244), .IN2(r798_n247), .Q(r798_n246) );
  NOR2X0 r798_U261 ( .QN(P1_N2148), .IN1(r798_n245), .IN2(r798_n246) );
  NAND2X0 r798_U260 ( .IN1(P1_N5160), .IN2(r798_n244), .QN(r798_n241) );
  OR2X1 r798_U259 ( .IN2(P1_N5160), .IN1(r798_n244), .Q(r798_n243) );
  NAND2X0 r798_U258 ( .IN1(P1_N1996), .IN2(r798_n243), .QN(r798_n242) );
  NAND2X0 r798_U257 ( .IN1(r798_n241), .IN2(r798_n242), .QN(r798_n234) );
  OR2X1 r798_U255 ( .IN2(P1_N1997), .IN1(n7058), .Q(r798_n238) );
  NAND2X0 r798_U254 ( .IN1(P1_N1997), .IN2(n7058), .QN(r798_n239) );
  NAND2X0 r798_U253 ( .IN1(r798_n238), .IN2(r798_n239), .QN(r798_n237) );
  NOR2X0 r798_U252 ( .QN(r798_n235), .IN1(r798_n234), .IN2(r798_n237) );
  AND2X1 r798_U251 ( .IN1(r798_n234), .IN2(r798_n237), .Q(r798_n236) );
  NOR2X0 r798_U250 ( .QN(P1_N2149), .IN1(r798_n235), .IN2(r798_n236) );
  NAND2X0 r798_U249 ( .IN1(P1_N5161), .IN2(r798_n234), .QN(r798_n231) );
  OR2X1 r798_U248 ( .IN2(P1_N5161), .IN1(r798_n234), .Q(r798_n233) );
  NAND2X0 r798_U247 ( .IN1(P1_N1997), .IN2(r798_n233), .QN(r798_n232) );
  NAND2X0 r798_U246 ( .IN1(r798_n231), .IN2(r798_n232), .QN(r798_n224) );
  OR2X1 r798_U244 ( .IN2(P1_N1998), .IN1(n7056), .Q(r798_n228) );
  NAND2X0 r798_U243 ( .IN1(P1_N1998), .IN2(n7056), .QN(r798_n229) );
  INVX0 r798_U7 ( .ZN(r798_n314), .INP(n7138) );
endmodule

